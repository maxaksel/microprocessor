magic
tech scmos
timestamp 1682952543
<< metal1 >>
rect 14 4107 4211 4127
rect 38 4083 4187 4103
rect 14 4067 4211 4073
rect 108 4013 133 4016
rect 204 4013 237 4016
rect 388 4013 397 4016
rect 660 4013 677 4016
rect 778 4013 788 4016
rect 844 4013 853 4016
rect 890 4013 916 4016
rect 954 4013 964 4016
rect 994 4013 1020 4016
rect 1330 4013 1356 4016
rect 1524 4013 1549 4016
rect 1698 4013 1724 4016
rect 1762 4013 1780 4016
rect 2234 4013 2260 4016
rect 2340 4013 2365 4016
rect 2396 4013 2405 4016
rect 2412 4013 2421 4016
rect 2468 4013 2485 4016
rect 2524 4013 2533 4016
rect 2676 4013 2701 4016
rect 2706 4013 2716 4016
rect 2834 4013 2844 4016
rect 2882 4013 2908 4016
rect 2962 4013 2972 4016
rect 2978 4013 2996 4016
rect 3026 4013 3052 4016
rect 3106 4013 3132 4016
rect 3162 4013 3188 4016
rect 3516 4013 3533 4016
rect 3612 4013 3637 4016
rect 3804 4013 3829 4016
rect 3868 4013 3885 4016
rect 4100 4013 4117 4016
rect 196 4003 221 4006
rect 370 4003 380 4006
rect 1596 4003 1605 4006
rect 1642 4003 1652 4006
rect 2402 4005 2405 4013
rect 2690 4003 2708 4006
rect 2818 4003 2836 4006
rect 2978 4005 2981 4013
rect 3106 4005 3109 4013
rect 38 3967 4187 3973
rect 978 3943 1004 3946
rect 308 3933 349 3936
rect 354 3933 364 3936
rect 380 3933 389 3936
rect 498 3926 501 3936
rect 524 3933 557 3936
rect 572 3933 597 3936
rect 666 3933 676 3936
rect 724 3933 740 3936
rect 762 3933 772 3936
rect 820 3933 829 3936
rect 858 3933 868 3936
rect 900 3933 916 3936
rect 938 3933 948 3936
rect 1058 3933 1068 3936
rect 1098 3926 1101 3936
rect 1106 3933 1116 3936
rect 1146 3933 1164 3936
rect 1202 3933 1212 3936
rect 1228 3933 1244 3936
rect 1298 3933 1316 3936
rect 1338 3933 1364 3936
rect 1386 3933 1397 3936
rect 1426 3933 1452 3936
rect 1586 3933 1596 3936
rect 1612 3933 1636 3936
rect 1772 3933 1805 3936
rect 108 3923 117 3926
rect 220 3923 229 3926
rect 316 3923 325 3926
rect 338 3923 356 3926
rect 434 3923 444 3926
rect 474 3925 501 3926
rect 474 3923 500 3925
rect 532 3923 557 3926
rect 578 3923 596 3926
rect 628 3923 636 3926
rect 674 3923 684 3926
rect 786 3923 796 3926
rect 866 3923 876 3926
rect 956 3923 965 3926
rect 980 3923 1005 3926
rect 1060 3923 1069 3926
rect 1076 3923 1101 3926
rect 1340 3923 1356 3926
rect 1386 3925 1389 3933
rect 1394 3925 1397 3933
rect 2154 3926 2157 3935
rect 2186 3933 2204 3936
rect 2388 3933 2397 3936
rect 2402 3933 2412 3936
rect 2450 3933 2468 3936
rect 2530 3933 2540 3936
rect 2554 3933 2572 3936
rect 2722 3926 2725 3935
rect 2738 3933 2748 3936
rect 2820 3933 2828 3936
rect 2866 3933 2892 3936
rect 2930 3933 2956 3936
rect 3506 3933 3516 3936
rect 3594 3933 3612 3936
rect 3834 3926 3837 3935
rect 3930 3933 3980 3936
rect 1450 3923 1460 3926
rect 1466 3923 1516 3926
rect 1546 3923 1556 3926
rect 1794 3923 1804 3926
rect 1842 3923 1860 3926
rect 1906 3923 1916 3926
rect 1996 3923 2021 3926
rect 2092 3923 2117 3926
rect 2148 3923 2157 3926
rect 2164 3923 2197 3926
rect 2228 3923 2252 3926
rect 2492 3923 2548 3926
rect 2562 3923 2580 3926
rect 2586 3923 2596 3926
rect 2660 3923 2677 3926
rect 2716 3923 2725 3926
rect 2732 3923 2756 3926
rect 2786 3923 2796 3926
rect 2882 3923 2900 3926
rect 2938 3923 2964 3926
rect 3026 3923 3052 3926
rect 3258 3923 3268 3926
rect 3298 3923 3308 3926
rect 3338 3923 3348 3926
rect 3354 3923 3380 3926
rect 3442 3923 3468 3926
rect 3540 3923 3557 3926
rect 3594 3923 3620 3926
rect 3652 3923 3676 3926
rect 3772 3923 3797 3926
rect 3828 3923 3837 3926
rect 3850 3923 3860 3926
rect 3890 3923 3900 3926
rect 3954 3923 3988 3926
rect 14 3867 4211 3873
rect 122 3813 148 3816
rect 180 3813 205 3816
rect 226 3813 260 3816
rect 124 3803 141 3806
rect 146 3803 156 3806
rect 172 3803 197 3806
rect 268 3803 285 3806
rect 314 3803 317 3814
rect 322 3813 332 3816
rect 556 3813 565 3816
rect 612 3813 621 3816
rect 748 3813 757 3816
rect 794 3813 820 3816
rect 1036 3813 1061 3816
rect 1100 3813 1109 3816
rect 1164 3813 1197 3816
rect 1442 3813 1468 3816
rect 1556 3813 1573 3816
rect 1578 3813 1588 3816
rect 1722 3813 1748 3816
rect 1834 3813 1852 3816
rect 1900 3813 1909 3816
rect 1922 3813 1956 3816
rect 2116 3813 2141 3816
rect 2172 3813 2181 3816
rect 2188 3813 2228 3816
rect 2266 3813 2284 3816
rect 2356 3813 2365 3816
rect 2484 3813 2509 3816
rect 2540 3813 2549 3816
rect 2556 3813 2580 3816
rect 2652 3813 2677 3816
rect 2714 3813 2732 3816
rect 2812 3813 2837 3816
rect 2868 3813 2877 3816
rect 2922 3813 2948 3816
rect 3076 3813 3101 3816
rect 3212 3813 3237 3816
rect 3282 3813 3292 3816
rect 3322 3813 3348 3816
rect 3484 3813 3509 3816
rect 3540 3813 3557 3816
rect 3564 3813 3573 3816
rect 3690 3813 3700 3816
rect 3812 3813 3861 3816
rect 4100 3813 4132 3816
rect 330 3803 340 3806
rect 362 3803 372 3806
rect 964 3803 973 3806
rect 1108 3803 1125 3806
rect 1130 3803 1140 3806
rect 1172 3803 1205 3806
rect 1234 3803 1252 3806
rect 1370 3803 1396 3806
rect 1538 3803 1548 3806
rect 1618 3803 1628 3806
rect 1650 3803 1676 3806
rect 1786 3803 1804 3806
rect 1842 3803 1860 3806
rect 1882 3803 1892 3806
rect 2178 3805 2181 3813
rect 2258 3803 2276 3806
rect 2314 3803 2348 3806
rect 2546 3805 2549 3813
rect 2874 3805 2877 3813
rect 3282 3805 3285 3813
rect 3554 3805 3557 3813
rect 3570 3805 3573 3813
rect 3770 3803 3788 3806
rect 3858 3805 3861 3813
rect 4140 3803 4149 3806
rect 38 3767 4187 3773
rect 922 3743 948 3746
rect 108 3723 133 3726
rect 170 3725 173 3736
rect 316 3733 325 3736
rect 556 3733 581 3736
rect 586 3733 596 3736
rect 612 3733 621 3736
rect 756 3733 789 3736
rect 812 3733 828 3736
rect 842 3733 868 3736
rect 890 3733 908 3736
rect 930 3733 956 3736
rect 1076 3733 1085 3736
rect 1108 3733 1132 3736
rect 1204 3733 1213 3736
rect 1218 3733 1228 3736
rect 1306 3733 1364 3736
rect 1386 3733 1396 3736
rect 2146 3726 2149 3735
rect 2244 3733 2277 3736
rect 2316 3733 2341 3736
rect 2346 3733 2364 3736
rect 2402 3733 2420 3736
rect 2458 3733 2468 3736
rect 2500 3733 2509 3736
rect 2602 3733 2612 3736
rect 2684 3733 2693 3736
rect 2690 3726 2693 3733
rect 2714 3733 2724 3736
rect 2820 3733 2829 3736
rect 3082 3733 3100 3736
rect 3132 3733 3141 3736
rect 3178 3733 3220 3736
rect 3348 3733 3364 3736
rect 2714 3726 2717 3733
rect 2826 3726 2829 3733
rect 3506 3726 3509 3735
rect 3562 3726 3565 3735
rect 3674 3726 3677 3735
rect 3794 3726 3797 3735
rect 244 3723 261 3726
rect 314 3723 324 3726
rect 468 3723 477 3726
rect 564 3723 573 3726
rect 762 3723 788 3726
rect 826 3723 860 3726
rect 1004 3723 1021 3726
rect 1116 3723 1125 3726
rect 1156 3723 1165 3726
rect 1236 3723 1245 3726
rect 1300 3723 1325 3726
rect 1330 3723 1356 3726
rect 1442 3723 1468 3726
rect 1530 3723 1540 3726
rect 1570 3723 1596 3726
rect 1634 3723 1644 3726
rect 1674 3723 1700 3726
rect 1834 3723 1844 3726
rect 2002 3723 2012 3726
rect 2084 3723 2109 3726
rect 2140 3723 2149 3726
rect 2156 3723 2196 3726
rect 2250 3723 2300 3726
rect 2410 3723 2428 3726
rect 2466 3723 2476 3726
rect 2506 3723 2524 3726
rect 2554 3723 2572 3726
rect 2602 3723 2620 3726
rect 2650 3723 2660 3726
rect 2690 3723 2717 3726
rect 2748 3723 2796 3726
rect 2826 3723 2836 3726
rect 2842 3723 2860 3726
rect 2890 3723 2900 3726
rect 2930 3723 2940 3726
rect 3146 3723 3164 3726
rect 3266 3723 3284 3726
rect 3314 3723 3324 3726
rect 3444 3723 3469 3726
rect 3500 3723 3509 3726
rect 3554 3723 3565 3726
rect 3612 3723 3637 3726
rect 3668 3723 3677 3726
rect 3684 3723 3700 3726
rect 3730 3723 3740 3726
rect 3794 3723 3805 3726
rect 3842 3723 3852 3726
rect 3882 3723 3892 3726
rect 3962 3723 3972 3726
rect 4002 3723 4012 3726
rect 14 3667 4211 3673
rect 2764 3623 2780 3626
rect 3028 3623 3036 3626
rect 3892 3623 3909 3626
rect 108 3613 133 3616
rect 220 3613 245 3616
rect 290 3613 308 3616
rect 340 3614 372 3616
rect 338 3613 372 3614
rect 404 3613 413 3616
rect 460 3613 485 3616
rect 602 3613 620 3616
rect 658 3613 668 3616
rect 842 3613 868 3616
rect 924 3613 949 3616
rect 1004 3613 1029 3616
rect 1090 3613 1108 3616
rect 1258 3613 1284 3616
rect 1322 3613 1332 3616
rect 1338 3613 1348 3616
rect 1434 3613 1460 3616
rect 1548 3613 1572 3616
rect 1636 3613 1645 3616
rect 1652 3613 1661 3616
rect 1668 3613 1677 3616
rect 1826 3613 1836 3616
rect 1850 3613 1876 3616
rect 1908 3613 1917 3616
rect 1932 3613 1949 3616
rect 1986 3613 2012 3616
rect 2092 3613 2117 3616
rect 2148 3613 2173 3616
rect 2180 3613 2196 3616
rect 2226 3613 2236 3616
rect 2276 3613 2285 3616
rect 2332 3613 2341 3616
rect 2394 3613 2404 3616
rect 2442 3613 2468 3616
rect 2530 3613 2564 3616
rect 2642 3613 2684 3616
rect 2738 3613 2748 3616
rect 2796 3613 2805 3616
rect 2844 3613 2861 3616
rect 2866 3613 2876 3616
rect 2898 3613 2917 3616
rect 2994 3613 3012 3616
rect 3052 3613 3061 3616
rect 3186 3613 3196 3616
rect 3210 3613 3220 3616
rect 3348 3613 3373 3616
rect 3404 3613 3413 3616
rect 3420 3613 3436 3616
rect 3562 3613 3572 3616
rect 3612 3613 3637 3616
rect 3668 3613 3677 3616
rect 3684 3613 3708 3616
rect 3754 3613 3764 3616
rect 3818 3613 3836 3616
rect 292 3603 309 3606
rect 338 3603 341 3613
rect 402 3603 436 3606
rect 468 3603 485 3606
rect 594 3603 628 3606
rect 650 3603 660 3606
rect 748 3603 764 3606
rect 786 3603 796 3606
rect 956 3603 965 3606
rect 1076 3603 1109 3606
rect 1132 3603 1172 3606
rect 1204 3603 1221 3606
rect 1346 3603 1356 3606
rect 1378 3603 1388 3606
rect 1634 3603 1644 3606
rect 1778 3603 1796 3606
rect 1858 3603 1884 3606
rect 1906 3603 1924 3606
rect 2170 3605 2173 3613
rect 2338 3605 2341 3613
rect 2420 3603 2453 3606
rect 2498 3603 2508 3606
rect 2532 3603 2549 3606
rect 2594 3603 2620 3606
rect 2644 3603 2661 3606
rect 2666 3603 2676 3606
rect 2730 3603 2740 3606
rect 2810 3603 2836 3606
rect 2892 3603 2917 3606
rect 3202 3603 3212 3606
rect 3410 3605 3413 3613
rect 3674 3605 3677 3613
rect 3922 3606 3925 3625
rect 3738 3603 3756 3606
rect 3852 3603 3869 3606
rect 3890 3603 3908 3606
rect 3922 3603 3932 3606
rect 4010 3603 4020 3606
rect 922 3593 948 3596
rect 962 3593 965 3603
rect 2666 3596 2669 3603
rect 2650 3593 2669 3596
rect 38 3567 4187 3573
rect 842 3543 860 3546
rect 874 3543 892 3546
rect 906 3543 924 3546
rect 938 3543 956 3546
rect 3706 3543 3733 3546
rect 180 3533 189 3536
rect 258 3533 268 3536
rect 378 3526 381 3535
rect 418 3533 436 3536
rect 108 3523 117 3526
rect 178 3523 188 3526
rect 372 3523 381 3526
rect 434 3523 444 3526
rect 618 3525 621 3536
rect 650 3533 668 3536
rect 722 3533 732 3536
rect 786 3533 804 3536
rect 836 3533 845 3536
rect 868 3533 885 3536
rect 900 3533 909 3536
rect 964 3533 981 3536
rect 1100 3533 1117 3536
rect 666 3523 676 3526
rect 748 3523 764 3526
rect 794 3523 812 3526
rect 876 3523 893 3526
rect 908 3523 925 3526
rect 940 3523 949 3526
rect 972 3523 989 3526
rect 1028 3523 1037 3526
rect 1098 3523 1116 3526
rect 1146 3525 1149 3536
rect 1154 3533 1164 3536
rect 1186 3533 1196 3536
rect 1346 3525 1349 3536
rect 1378 3533 1388 3536
rect 1532 3533 1549 3536
rect 1588 3533 1613 3536
rect 1380 3523 1389 3526
rect 1434 3523 1460 3526
rect 1594 3523 1612 3526
rect 1642 3525 1645 3536
rect 1746 3533 1764 3536
rect 1682 3523 1708 3526
rect 1786 3525 1789 3536
rect 1914 3533 1948 3536
rect 1978 3533 2004 3536
rect 2306 3533 2332 3536
rect 2370 3533 2388 3536
rect 2466 3533 2484 3536
rect 2514 3533 2532 3536
rect 2570 3533 2604 3536
rect 2628 3533 2645 3536
rect 2650 3533 2660 3536
rect 2698 3533 2732 3536
rect 2756 3533 2765 3536
rect 2820 3533 2852 3536
rect 2890 3533 2908 3536
rect 2988 3533 2997 3536
rect 3042 3533 3060 3536
rect 3098 3533 3108 3536
rect 3146 3533 3188 3536
rect 3300 3533 3317 3536
rect 3332 3533 3356 3536
rect 3380 3533 3389 3536
rect 3530 3533 3548 3536
rect 3572 3533 3604 3536
rect 3618 3533 3652 3536
rect 3676 3533 3709 3536
rect 3778 3533 3788 3536
rect 3812 3533 3845 3536
rect 3906 3533 3916 3536
rect 1804 3523 1813 3526
rect 1858 3523 1876 3526
rect 2050 3523 2076 3526
rect 2148 3523 2173 3526
rect 2218 3523 2236 3526
rect 2386 3523 2396 3526
rect 2482 3523 2492 3526
rect 2514 3523 2540 3526
rect 2602 3523 2612 3526
rect 2626 3523 2668 3526
rect 2706 3523 2740 3526
rect 2754 3523 2796 3526
rect 2916 3523 2949 3526
rect 3010 3523 3020 3526
rect 3068 3523 3101 3526
rect 2756 3513 2781 3516
rect 3314 3515 3317 3533
rect 3372 3523 3381 3526
rect 3386 3523 3404 3526
rect 3538 3523 3556 3526
rect 3330 3513 3356 3516
rect 3572 3513 3581 3516
rect 3618 3515 3621 3533
rect 3668 3523 3677 3526
rect 3786 3523 3796 3526
rect 3868 3523 3901 3526
rect 3938 3523 3956 3526
rect 3986 3523 3996 3526
rect 3634 3513 3652 3516
rect 3812 3513 3852 3516
rect 14 3467 4211 3473
rect 2522 3423 2532 3426
rect 2644 3423 2661 3426
rect 114 3413 124 3416
rect 138 3413 156 3416
rect 530 3413 540 3416
rect 132 3403 149 3406
rect 180 3403 189 3406
rect 306 3403 332 3406
rect 348 3403 365 3406
rect 570 3403 573 3414
rect 644 3413 669 3416
rect 802 3413 820 3416
rect 914 3413 932 3416
rect 988 3413 1069 3416
rect 1116 3413 1133 3416
rect 1148 3413 1157 3416
rect 1218 3413 1228 3416
rect 1292 3413 1333 3416
rect 1420 3413 1445 3416
rect 1530 3406 1533 3414
rect 1538 3413 1564 3416
rect 1594 3413 1604 3416
rect 1610 3413 1620 3416
rect 1676 3413 1685 3416
rect 1722 3413 1748 3416
rect 1786 3413 1796 3416
rect 1834 3413 1852 3416
rect 1964 3413 1981 3416
rect 2074 3413 2092 3416
rect 2130 3413 2140 3416
rect 2212 3413 2221 3416
rect 2244 3413 2285 3416
rect 2330 3413 2357 3416
rect 2442 3413 2452 3416
rect 2484 3413 2493 3416
rect 2508 3413 2533 3416
rect 2548 3413 2572 3416
rect 2586 3413 2604 3416
rect 2618 3413 2629 3416
rect 2676 3413 2708 3416
rect 2722 3413 2749 3416
rect 2756 3413 2765 3416
rect 2770 3413 2788 3416
rect 2794 3413 2804 3416
rect 2834 3413 2860 3416
rect 2914 3413 2932 3416
rect 2962 3413 2972 3416
rect 2986 3413 3012 3416
rect 3044 3413 3061 3416
rect 756 3403 765 3406
rect 788 3403 828 3406
rect 850 3403 860 3406
rect 1084 3403 1101 3406
rect 1108 3403 1117 3406
rect 1122 3403 1140 3406
rect 1300 3403 1356 3406
rect 1492 3403 1501 3406
rect 1530 3403 1549 3406
rect 1610 3403 1628 3406
rect 1644 3403 1653 3406
rect 1658 3403 1668 3406
rect 1890 3403 1916 3406
rect 2250 3403 2292 3406
rect 2324 3403 2349 3406
rect 2354 3405 2357 3413
rect 2394 3403 2412 3406
rect 2516 3403 2525 3406
rect 2618 3405 2621 3413
rect 2684 3403 2693 3406
rect 2722 3405 2725 3413
rect 2738 3403 2748 3406
rect 2794 3405 2797 3413
rect 3106 3406 3109 3425
rect 3114 3423 3140 3426
rect 3290 3423 3316 3426
rect 3330 3423 3348 3426
rect 3644 3423 3653 3426
rect 3196 3413 3205 3416
rect 3266 3413 3276 3416
rect 3282 3413 3324 3416
rect 3394 3413 3405 3416
rect 3484 3413 3501 3416
rect 3642 3413 3700 3416
rect 3746 3413 3764 3416
rect 3810 3413 3820 3416
rect 3874 3413 3892 3416
rect 2988 3403 3005 3406
rect 3020 3403 3029 3406
rect 3050 3403 3092 3406
rect 3106 3403 3140 3406
rect 3284 3403 3293 3406
rect 3332 3403 3348 3406
rect 3372 3403 3397 3406
rect 3402 3405 3405 3413
rect 3898 3406 3901 3425
rect 3946 3413 3965 3416
rect 3492 3403 3501 3406
rect 3506 3403 3524 3406
rect 3610 3403 3620 3406
rect 3682 3403 3692 3406
rect 3730 3403 3756 3406
rect 3794 3403 3812 3406
rect 3858 3403 3884 3406
rect 3898 3403 3916 3406
rect 3940 3403 3957 3406
rect 3962 3405 3965 3413
rect 4002 3413 4036 3416
rect 4066 3413 4076 3416
rect 4082 3413 4100 3416
rect 4002 3406 4005 3413
rect 3996 3403 4005 3406
rect 4010 3403 4028 3406
rect 4084 3403 4093 3406
rect 4108 3403 4133 3406
rect 986 3393 1076 3396
rect 1090 3393 1100 3396
rect 1338 3393 1341 3403
rect 38 3367 4187 3373
rect 180 3333 189 3336
rect 108 3323 133 3326
rect 178 3323 188 3326
rect 218 3325 221 3336
rect 236 3333 245 3336
rect 268 3333 277 3336
rect 796 3333 829 3336
rect 866 3333 892 3336
rect 1140 3333 1180 3336
rect 1370 3333 1380 3336
rect 1524 3333 1533 3336
rect 1548 3333 1557 3336
rect 1580 3333 1629 3336
rect 1770 3333 1780 3336
rect 292 3323 301 3326
rect 420 3323 429 3326
rect 700 3323 725 3326
rect 818 3323 828 3326
rect 860 3323 877 3326
rect 938 3323 964 3326
rect 1092 3323 1109 3326
rect 1204 3323 1213 3326
rect 1218 3323 1236 3326
rect 1292 3323 1317 3326
rect 1362 3323 1372 3326
rect 1444 3323 1469 3326
rect 1530 3323 1540 3326
rect 1546 3323 1556 3326
rect 1594 3323 1636 3326
rect 1682 3323 1692 3326
rect 1730 3323 1756 3326
rect 1802 3325 1805 3336
rect 1810 3333 1820 3336
rect 1954 3333 1996 3336
rect 2124 3333 2133 3336
rect 2300 3333 2324 3336
rect 2546 3334 2564 3336
rect 1828 3323 1837 3326
rect 1954 3323 1957 3333
rect 2188 3323 2213 3326
rect 2258 3323 2276 3326
rect 2348 3323 2372 3326
rect 2428 3323 2453 3326
rect 2490 3323 2493 3334
rect 2546 3333 2565 3334
rect 2594 3333 2604 3336
rect 2618 3333 2628 3336
rect 2540 3323 2549 3326
rect 2562 3323 2565 3333
rect 2722 3326 2725 3334
rect 2804 3333 2812 3336
rect 2858 3326 2861 3334
rect 2900 3333 2908 3336
rect 3058 3333 3068 3336
rect 3258 3333 3268 3336
rect 3058 3326 3061 3333
rect 2572 3323 2581 3326
rect 2594 3323 2612 3326
rect 2650 3323 2677 3326
rect 2716 3323 2725 3326
rect 2764 3323 2788 3326
rect 2858 3323 2869 3326
rect 3052 3323 3061 3326
rect 3092 3323 3101 3326
rect 3140 3323 3165 3326
rect 3202 3323 3220 3326
rect 3250 3323 3276 3326
rect 3298 3323 3301 3334
rect 3410 3326 3413 3334
rect 3618 3333 3644 3336
rect 3668 3333 3693 3336
rect 3348 3323 3373 3326
rect 3404 3323 3413 3326
rect 3420 3323 3436 3326
rect 3602 3323 3612 3326
rect 2548 3313 2557 3316
rect 2594 3315 2597 3323
rect 2650 3315 2653 3323
rect 2674 3315 2677 3323
rect 2748 3313 2757 3316
rect 3618 3315 3621 3333
rect 3698 3326 3701 3334
rect 3660 3323 3669 3326
rect 3690 3323 3701 3326
rect 3738 3323 3741 3334
rect 3906 3326 3909 3334
rect 3996 3333 4005 3336
rect 3898 3323 3909 3326
rect 3626 3313 3644 3316
rect 14 3267 4211 3273
rect 2674 3223 2684 3226
rect 2746 3216 2749 3225
rect 2908 3223 2916 3226
rect 4092 3223 4100 3226
rect 108 3213 133 3216
rect 178 3213 188 3216
rect 418 3213 444 3216
rect 482 3213 500 3216
rect 506 3213 532 3216
rect 612 3213 637 3216
rect 674 3213 692 3216
rect 740 3213 804 3216
rect 836 3213 845 3216
rect 850 3213 868 3216
rect 908 3213 925 3216
rect 940 3213 965 3216
rect 980 3213 1005 3216
rect 1034 3213 1052 3216
rect 1116 3213 1141 3216
rect 1178 3213 1188 3216
rect 1306 3213 1316 3216
rect 180 3203 189 3206
rect 362 3203 372 3206
rect 388 3203 436 3206
rect 508 3203 533 3206
rect 556 3203 573 3206
rect 700 3203 709 3206
rect 786 3203 812 3206
rect 834 3203 860 3206
rect 922 3203 932 3206
rect 972 3203 989 3206
rect 1010 3203 1020 3206
rect 1060 3203 1069 3206
rect 1108 3203 1148 3206
rect 1178 3205 1181 3213
rect 1292 3203 1317 3206
rect 1346 3203 1349 3214
rect 1418 3213 1444 3216
rect 1548 3213 1580 3216
rect 1610 3213 1620 3216
rect 1652 3213 1661 3216
rect 1668 3213 1677 3216
rect 1714 3213 1740 3216
rect 1778 3213 1788 3216
rect 1834 3213 1844 3216
rect 1874 3213 1900 3216
rect 2018 3213 2044 3216
rect 2156 3213 2181 3216
rect 2212 3213 2221 3216
rect 1834 3206 1837 3213
rect 1482 3203 1492 3206
rect 1514 3203 1524 3206
rect 1556 3203 1565 3206
rect 1604 3203 1613 3206
rect 1650 3203 1660 3206
rect 1812 3203 1837 3206
rect 2218 3205 2221 3213
rect 2266 3205 2269 3216
rect 2324 3213 2341 3216
rect 2612 3213 2637 3216
rect 2722 3206 2725 3214
rect 2730 3213 2740 3216
rect 2746 3213 2773 3216
rect 2828 3213 2853 3216
rect 2890 3213 2900 3216
rect 2930 3213 2940 3216
rect 2978 3213 2996 3216
rect 3068 3213 3085 3216
rect 3124 3213 3133 3216
rect 3162 3213 3172 3216
rect 3244 3213 3261 3216
rect 3330 3213 3340 3216
rect 3444 3213 3453 3216
rect 3484 3213 3501 3216
rect 3514 3213 3532 3216
rect 3572 3213 3612 3216
rect 3668 3213 3692 3216
rect 2700 3203 2716 3206
rect 2722 3203 2732 3206
rect 2746 3203 2756 3206
rect 2930 3205 2933 3213
rect 3130 3205 3133 3213
rect 3258 3206 3261 3213
rect 3258 3203 3268 3206
rect 3450 3205 3453 3213
rect 3466 3203 3476 3206
rect 3716 3203 3733 3206
rect 3738 3205 3741 3216
rect 3818 3213 3844 3216
rect 3930 3213 3964 3216
rect 4066 3213 4084 3216
rect 4066 3203 4076 3206
rect 4116 3203 4149 3206
rect 874 3193 892 3196
rect 914 3193 924 3196
rect 938 3193 964 3196
rect 978 3193 1012 3196
rect 1610 3183 1613 3203
rect 38 3167 4187 3173
rect 914 3143 924 3146
rect 2826 3143 2836 3146
rect 180 3133 189 3136
rect 364 3133 381 3136
rect 386 3133 396 3136
rect 530 3133 540 3136
rect 682 3133 700 3136
rect 738 3133 756 3136
rect 788 3133 797 3136
rect 908 3133 917 3136
rect 1068 3133 1085 3136
rect 1090 3133 1100 3136
rect 1116 3133 1164 3136
rect 1196 3133 1213 3136
rect 1314 3133 1324 3136
rect 794 3126 797 3133
rect 108 3123 133 3126
rect 372 3123 389 3126
rect 468 3123 485 3126
rect 604 3123 629 3126
rect 666 3123 676 3126
rect 738 3123 764 3126
rect 794 3123 804 3126
rect 850 3123 860 3126
rect 940 3123 949 3126
rect 988 3123 1005 3126
rect 1346 3125 1349 3136
rect 1354 3133 1372 3136
rect 1612 3133 1621 3136
rect 1650 3133 1660 3136
rect 2196 3133 2205 3136
rect 2330 3126 2333 3135
rect 2378 3133 2396 3136
rect 2412 3133 2429 3136
rect 2660 3133 2708 3136
rect 2962 3133 2980 3136
rect 2994 3133 3012 3136
rect 3060 3133 3084 3136
rect 3114 3133 3132 3136
rect 3244 3133 3253 3136
rect 3380 3133 3389 3136
rect 3788 3133 3797 3136
rect 2426 3126 2429 3133
rect 1418 3123 1444 3126
rect 1578 3123 1588 3126
rect 1668 3123 1685 3126
rect 1722 3123 1748 3126
rect 1794 3123 1812 3126
rect 1842 3123 1868 3126
rect 1954 3123 1972 3126
rect 2114 3123 2124 3126
rect 2172 3123 2180 3126
rect 2260 3123 2285 3126
rect 2330 3123 2348 3126
rect 2426 3123 2444 3126
rect 2474 3123 2500 3126
rect 2538 3123 2548 3126
rect 2578 3123 2604 3126
rect 2706 3123 2716 3126
rect 3010 3123 3013 3133
rect 3266 3126 3269 3133
rect 3108 3123 3133 3126
rect 3258 3123 3269 3126
rect 3524 3123 3549 3126
rect 3620 3123 3645 3126
rect 3842 3123 3852 3126
rect 3900 3123 3909 3126
rect 3996 3123 4021 3126
rect 3258 3093 3261 3123
rect 14 3067 4211 3073
rect 2746 3023 2756 3026
rect 2810 3023 2820 3026
rect 3244 3023 3261 3026
rect 4026 3016 4029 3036
rect 108 3013 133 3016
rect 170 3013 212 3016
rect 186 3003 204 3006
rect 250 3003 253 3014
rect 284 3013 293 3016
rect 436 3013 461 3016
rect 276 3003 301 3006
rect 508 3003 517 3006
rect 564 3003 573 3006
rect 610 3003 613 3014
rect 684 3013 709 3016
rect 740 3013 749 3016
rect 954 3013 964 3016
rect 1116 3013 1125 3016
rect 1244 3013 1253 3016
rect 1308 3013 1317 3016
rect 1322 3013 1340 3016
rect 1386 3013 1396 3016
rect 1434 3013 1460 3016
rect 1508 3013 1517 3016
rect 1578 3013 1588 3016
rect 1674 3013 1700 3016
rect 1778 3013 1788 3016
rect 1858 3013 1876 3016
rect 1978 3013 1988 3016
rect 2060 3013 2077 3016
rect 2156 3013 2181 3016
rect 2274 3013 2285 3016
rect 2338 3013 2348 3016
rect 2354 3013 2381 3016
rect 2578 3013 2588 3016
rect 2716 3013 2725 3016
rect 2740 3013 2764 3016
rect 2804 3013 2828 3016
rect 2852 3013 2861 3016
rect 2868 3013 2877 3016
rect 2908 3013 2917 3016
rect 2932 3013 2949 3016
rect 3034 3013 3060 3016
rect 3098 3013 3132 3016
rect 3170 3013 3180 3016
rect 636 3003 645 3006
rect 796 3003 805 3006
rect 858 3003 876 3006
rect 1012 3003 1021 3006
rect 1066 3003 1092 3006
rect 1108 3003 1156 3006
rect 1188 3003 1229 3006
rect 1250 3003 1284 3006
rect 1306 3003 1348 3006
rect 1370 3003 1388 3006
rect 1556 3003 1573 3006
rect 1578 2996 1581 3013
rect 1586 3003 1596 3006
rect 1618 3003 1628 3006
rect 1738 3003 1748 3006
rect 1770 3003 1780 3006
rect 1826 3003 1836 3006
rect 1858 3003 1884 3006
rect 1906 3003 1916 3006
rect 2268 3003 2277 3006
rect 2282 3005 2285 3013
rect 2316 3003 2325 3006
rect 2378 3005 2381 3013
rect 2722 3003 2732 3006
rect 2772 3003 2781 3006
rect 2938 3003 2948 3006
rect 2994 3003 3012 3006
rect 3050 3003 3068 3006
rect 3084 3003 3125 3006
rect 3156 3003 3173 3006
rect 3250 3003 3276 3006
rect 3298 3003 3301 3014
rect 3306 3013 3340 3016
rect 3372 3013 3381 3016
rect 3402 3013 3412 3016
rect 3314 3003 3348 3006
rect 3370 3003 3420 3006
rect 1122 2993 1149 2996
rect 1570 2993 1581 2996
rect 3426 2996 3429 3016
rect 3434 3013 3468 3016
rect 3498 3006 3501 3014
rect 3506 3013 3516 3016
rect 3658 3013 3668 3016
rect 3898 3013 3916 3016
rect 4026 3013 4037 3016
rect 4034 3007 4037 3013
rect 3466 3003 3476 3006
rect 3498 3003 3509 3006
rect 3644 3003 3653 3006
rect 4020 3003 4029 3006
rect 3426 2995 3437 2996
rect 3428 2993 3437 2995
rect 38 2967 4187 2973
rect 850 2943 860 2946
rect 3244 2943 3261 2946
rect 3850 2943 3860 2946
rect 140 2933 149 2936
rect 180 2933 189 2936
rect 306 2933 324 2936
rect 346 2933 356 2936
rect 626 2933 636 2936
rect 642 2933 652 2936
rect 714 2933 741 2936
rect 842 2933 868 2936
rect 138 2923 156 2926
rect 188 2923 205 2926
rect 348 2923 357 2926
rect 492 2923 501 2926
rect 540 2923 557 2926
rect 650 2923 660 2926
rect 708 2923 733 2926
rect 738 2923 748 2926
rect 794 2923 804 2926
rect 882 2923 892 2926
rect 932 2923 949 2926
rect 988 2923 997 2926
rect 1092 2923 1109 2926
rect 1114 2925 1117 2936
rect 1146 2925 1149 2936
rect 1324 2933 1333 2936
rect 1586 2933 1596 2936
rect 1618 2933 1628 2936
rect 1834 2933 1844 2936
rect 2290 2933 2300 2936
rect 2842 2933 2852 2936
rect 2890 2933 2900 2936
rect 3010 2926 3013 2935
rect 3194 2933 3228 2936
rect 3316 2933 3333 2936
rect 1188 2923 1197 2926
rect 1276 2923 1285 2926
rect 1316 2923 1325 2926
rect 1418 2923 1444 2926
rect 1506 2923 1516 2926
rect 1546 2923 1556 2926
rect 1620 2923 1629 2926
rect 1674 2923 1700 2926
rect 1778 2923 1796 2926
rect 2212 2923 2237 2926
rect 2268 2923 2277 2926
rect 2284 2923 2301 2926
rect 2762 2923 2788 2926
rect 2844 2923 2860 2926
rect 2866 2923 2884 2926
rect 2898 2923 2908 2926
rect 2980 2923 3013 2926
rect 3020 2923 3029 2926
rect 3202 2923 3220 2926
rect 3250 2923 3276 2926
rect 3298 2923 3308 2926
rect 3322 2923 3340 2926
rect 3370 2925 3373 2936
rect 3386 2933 3404 2936
rect 3378 2923 3396 2926
rect 3530 2925 3533 2936
rect 3562 2933 3572 2936
rect 3594 2925 3597 2936
rect 3634 2933 3644 2936
rect 3876 2933 3916 2936
rect 3938 2933 3956 2936
rect 3970 2933 3980 2936
rect 4018 2933 4036 2936
rect 3714 2923 3732 2926
rect 3738 2923 3748 2926
rect 3794 2923 3804 2926
rect 3850 2923 3860 2926
rect 3932 2923 3949 2926
rect 3954 2923 3964 2926
rect 4004 2923 4013 2926
rect 4060 2923 4077 2926
rect 2892 2913 2901 2916
rect 3188 2913 3213 2916
rect 3490 2913 3500 2916
rect 3738 2915 3741 2923
rect 4066 2913 4084 2916
rect 2922 2903 2940 2906
rect 3044 2903 3053 2906
rect 3484 2903 3509 2906
rect 14 2867 4211 2873
rect 2994 2833 3036 2836
rect 3506 2826 3509 2836
rect 108 2813 133 2816
rect 218 2803 221 2814
rect 260 2813 285 2816
rect 330 2813 340 2816
rect 332 2803 341 2806
rect 370 2803 373 2814
rect 506 2805 509 2816
rect 548 2813 573 2816
rect 610 2803 620 2806
rect 642 2803 645 2814
rect 658 2805 661 2816
rect 780 2813 797 2816
rect 802 2813 820 2816
rect 884 2813 901 2816
rect 940 2813 965 2816
rect 970 2813 988 2816
rect 1034 2813 1060 2816
rect 700 2803 740 2806
rect 762 2803 772 2806
rect 786 2803 828 2806
rect 844 2803 861 2806
rect 866 2803 876 2806
rect 898 2803 901 2813
rect 1146 2806 1149 2826
rect 2386 2816 2389 2825
rect 2860 2823 2877 2826
rect 2938 2823 2964 2826
rect 2988 2823 3013 2826
rect 3420 2823 3437 2826
rect 3506 2823 3516 2826
rect 2938 2816 2941 2823
rect 3562 2816 3565 2825
rect 3978 2823 3988 2826
rect 4068 2823 4084 2826
rect 1154 2813 1164 2816
rect 1234 2813 1260 2816
rect 1354 2813 1380 2816
rect 1426 2813 1436 2816
rect 1498 2813 1516 2816
rect 1354 2806 1357 2813
rect 1028 2803 1061 2806
rect 1090 2803 1116 2806
rect 1132 2803 1141 2806
rect 1146 2803 1156 2806
rect 1170 2803 1188 2806
rect 1298 2803 1324 2806
rect 1340 2803 1357 2806
rect 1500 2803 1517 2806
rect 1554 2805 1557 2816
rect 1666 2813 1684 2816
rect 1884 2813 1893 2816
rect 1898 2813 1908 2816
rect 1938 2813 1956 2816
rect 1996 2813 2005 2816
rect 2052 2813 2061 2816
rect 2092 2813 2101 2816
rect 2108 2813 2117 2816
rect 2170 2813 2196 2816
rect 2268 2813 2293 2816
rect 2058 2806 2061 2813
rect 1620 2803 1636 2806
rect 1668 2803 1677 2806
rect 1788 2803 1797 2806
rect 1820 2803 1844 2806
rect 2058 2803 2068 2806
rect 914 2793 924 2796
rect 2114 2795 2117 2813
rect 2330 2807 2333 2816
rect 2364 2813 2373 2816
rect 2386 2813 2396 2816
rect 2442 2813 2452 2816
rect 2594 2813 2604 2816
rect 2676 2813 2685 2816
rect 2932 2813 2941 2816
rect 2370 2807 2373 2813
rect 3178 2807 3181 2816
rect 3220 2813 3229 2816
rect 3346 2813 3356 2816
rect 3386 2813 3404 2816
rect 3418 2807 3421 2816
rect 3442 2813 3452 2816
rect 3466 2813 3492 2816
rect 3498 2813 3524 2816
rect 3538 2813 3548 2816
rect 3562 2813 3580 2816
rect 3602 2813 3645 2816
rect 3748 2813 3757 2816
rect 3786 2806 3789 2814
rect 3794 2813 3820 2816
rect 3906 2806 3909 2814
rect 4018 2813 4036 2816
rect 4074 2813 4092 2816
rect 2346 2803 2356 2806
rect 2404 2803 2413 2806
rect 2900 2803 2917 2806
rect 2924 2803 2957 2806
rect 3154 2803 3180 2806
rect 3378 2803 3396 2806
rect 3588 2803 3613 2806
rect 3634 2803 3644 2806
rect 3674 2803 3684 2806
rect 3740 2803 3765 2806
rect 3786 2803 3805 2806
rect 3844 2803 3853 2806
rect 3874 2803 3892 2806
rect 3906 2803 3916 2806
rect 3972 2803 3981 2806
rect 4100 2803 4133 2806
rect 3706 2793 3724 2796
rect 4130 2793 4133 2803
rect 38 2767 4187 2773
rect 1002 2753 1029 2756
rect 802 2743 820 2746
rect 946 2743 980 2746
rect 2964 2743 2972 2746
rect 3490 2736 3493 2756
rect 108 2723 133 2726
rect 178 2723 181 2734
rect 218 2733 237 2736
rect 316 2733 333 2736
rect 362 2733 372 2736
rect 572 2733 597 2736
rect 740 2733 765 2736
rect 818 2733 828 2736
rect 218 2725 221 2733
rect 234 2725 237 2733
rect 268 2723 277 2726
rect 412 2723 421 2726
rect 500 2723 525 2726
rect 570 2723 596 2726
rect 668 2723 693 2726
rect 738 2723 764 2726
rect 834 2725 837 2736
rect 988 2733 1013 2736
rect 1060 2733 1069 2736
rect 1106 2733 1148 2736
rect 1106 2726 1109 2733
rect 884 2723 901 2726
rect 996 2723 1029 2726
rect 1100 2723 1109 2726
rect 1170 2725 1173 2736
rect 1202 2733 1228 2736
rect 1260 2733 1293 2736
rect 1314 2733 1340 2736
rect 1754 2733 1780 2736
rect 2066 2733 2084 2736
rect 2314 2733 2332 2736
rect 2338 2733 2348 2736
rect 2770 2733 2812 2736
rect 2884 2733 2893 2736
rect 2900 2733 2909 2736
rect 2956 2733 2973 2736
rect 2986 2733 3020 2736
rect 3300 2733 3317 2736
rect 3330 2733 3340 2736
rect 3452 2733 3461 2736
rect 3490 2733 3500 2736
rect 3612 2733 3645 2736
rect 3914 2733 3924 2736
rect 3938 2733 3964 2736
rect 4002 2733 4028 2736
rect 1308 2723 1325 2726
rect 1364 2723 1380 2726
rect 1420 2723 1429 2726
rect 1634 2723 1644 2726
rect 1682 2723 1692 2726
rect 1698 2723 1708 2726
rect 1890 2723 1900 2726
rect 2092 2723 2116 2726
rect 2154 2723 2172 2726
rect 2308 2723 2325 2726
rect 2340 2723 2349 2726
rect 2356 2723 2380 2726
rect 2474 2723 2492 2726
rect 2530 2723 2533 2733
rect 2546 2723 2556 2726
rect 2748 2723 2757 2726
rect 2764 2723 2805 2726
rect 1754 2713 1781 2716
rect 1970 2713 1996 2716
rect 2396 2713 2404 2716
rect 2826 2713 2836 2716
rect 2842 2706 2845 2725
rect 2866 2723 2876 2726
rect 2882 2723 2892 2726
rect 2940 2723 2948 2726
rect 2988 2723 3045 2726
rect 3178 2723 3181 2733
rect 3188 2723 3205 2726
rect 3258 2723 3261 2733
rect 3338 2726 3341 2733
rect 3266 2723 3292 2726
rect 3298 2723 3341 2726
rect 3498 2723 3501 2733
rect 3650 2723 3660 2726
rect 3940 2723 3949 2726
rect 3980 2723 4013 2726
rect 4018 2723 4036 2726
rect 2860 2713 2869 2716
rect 3042 2713 3052 2716
rect 3076 2713 3117 2716
rect 3196 2713 3205 2716
rect 3274 2713 3284 2716
rect 4018 2713 4021 2723
rect 2826 2703 2845 2706
rect 3034 2703 3068 2706
rect 3082 2703 3140 2706
rect 14 2667 4211 2673
rect 1892 2633 1925 2636
rect 1940 2633 1965 2636
rect 2026 2633 2044 2636
rect 610 2623 621 2626
rect 610 2616 613 2623
rect 116 2613 124 2616
rect 154 2605 157 2616
rect 554 2613 572 2616
rect 604 2613 613 2616
rect 618 2613 636 2616
rect 666 2613 700 2616
rect 780 2613 829 2616
rect 924 2613 949 2616
rect 978 2613 988 2616
rect 1010 2606 1013 2626
rect 1842 2623 1852 2626
rect 1100 2613 1125 2616
rect 1156 2613 1165 2616
rect 1250 2613 1292 2616
rect 1322 2613 1348 2616
rect 1386 2613 1396 2616
rect 1418 2613 1428 2616
rect 354 2603 364 2606
rect 386 2603 396 2606
rect 556 2603 573 2606
rect 724 2603 757 2606
rect 762 2603 772 2606
rect 786 2603 828 2606
rect 860 2603 901 2606
rect 1005 2603 1013 2606
rect 1044 2603 1061 2606
rect 1210 2603 1220 2606
rect 1250 2605 1253 2613
rect 1418 2606 1421 2613
rect 1412 2603 1421 2606
rect 1498 2605 1501 2616
rect 1756 2613 1773 2616
rect 2010 2613 2020 2616
rect 2098 2613 2125 2616
rect 2196 2613 2221 2616
rect 2298 2613 2316 2616
rect 2098 2606 2101 2613
rect 2346 2607 2349 2616
rect 2666 2613 2684 2616
rect 2858 2613 2900 2616
rect 3100 2613 3125 2616
rect 3194 2613 3220 2616
rect 3284 2613 3293 2616
rect 3410 2613 3420 2616
rect 3538 2613 3556 2616
rect 3786 2613 3804 2616
rect 4140 2613 4149 2616
rect 1644 2603 1661 2606
rect 2058 2603 2084 2606
rect 2090 2603 2101 2606
rect 2122 2603 2132 2606
rect 2162 2603 2172 2606
rect 2210 2603 2228 2606
rect 2258 2603 2268 2606
rect 730 2593 764 2596
rect 866 2593 908 2596
rect 2394 2595 2397 2606
rect 2404 2603 2413 2606
rect 2860 2603 2869 2606
rect 3524 2603 3533 2606
rect 3660 2603 3685 2606
rect 4148 2603 4221 2606
rect 38 2567 4187 2573
rect 730 2543 764 2546
rect 1018 2536 1021 2546
rect 634 2533 644 2536
rect 666 2533 692 2536
rect 724 2533 741 2536
rect 746 2533 772 2536
rect 836 2533 853 2536
rect 996 2533 1021 2536
rect 1106 2533 1116 2536
rect 1266 2533 1276 2536
rect 1292 2533 1309 2536
rect 1322 2533 1340 2536
rect 1362 2533 1372 2536
rect 1402 2533 1428 2536
rect 1490 2533 1508 2536
rect 634 2526 637 2533
rect 108 2523 117 2526
rect 324 2523 349 2526
rect 428 2523 437 2526
rect 532 2523 549 2526
rect 588 2523 597 2526
rect 620 2523 637 2526
rect 660 2523 693 2526
rect 780 2523 813 2526
rect 884 2523 901 2526
rect 954 2523 972 2526
rect 1005 2523 1029 2526
rect 1124 2523 1141 2526
rect 1242 2523 1268 2526
rect 1300 2523 1309 2526
rect 1388 2523 1413 2526
rect 1450 2523 1468 2526
rect 1562 2523 1565 2534
rect 1594 2533 1612 2536
rect 1628 2533 1677 2536
rect 1578 2523 1604 2526
rect 1690 2523 1693 2534
rect 1706 2533 1748 2536
rect 1764 2533 1797 2536
rect 1706 2523 1740 2526
rect 1850 2523 1876 2526
rect 1962 2523 1972 2526
rect 2052 2523 2077 2526
rect 2114 2525 2117 2536
rect 2146 2533 2172 2536
rect 2186 2533 2204 2536
rect 2218 2533 2228 2536
rect 2274 2533 2292 2536
rect 2322 2533 2332 2536
rect 2370 2534 2380 2536
rect 2370 2533 2381 2534
rect 2402 2533 2412 2536
rect 2442 2533 2468 2536
rect 2482 2533 2500 2536
rect 2522 2533 2532 2536
rect 2554 2533 2580 2536
rect 2602 2533 2629 2536
rect 2666 2533 2684 2536
rect 2378 2526 2381 2533
rect 2882 2526 2885 2534
rect 3052 2533 3060 2536
rect 3100 2533 3109 2536
rect 3138 2533 3149 2536
rect 3178 2533 3188 2536
rect 3380 2533 3388 2536
rect 3708 2533 3716 2536
rect 3802 2533 3812 2536
rect 2154 2523 2180 2526
rect 2212 2523 2221 2526
rect 2252 2523 2277 2526
rect 2316 2523 2325 2526
rect 2356 2523 2381 2526
rect 2394 2523 2404 2526
rect 2540 2523 2549 2526
rect 2604 2523 2628 2526
rect 2882 2523 2893 2526
rect 2914 2523 2924 2526
rect 2980 2523 2989 2526
rect 2996 2523 3005 2526
rect 3098 2523 3108 2526
rect 3138 2525 3141 2533
rect 3914 2526 3917 2534
rect 3970 2533 3980 2536
rect 4002 2533 4012 2536
rect 3180 2523 3189 2526
rect 3268 2523 3285 2526
rect 3324 2523 3333 2526
rect 3356 2523 3381 2526
rect 3684 2523 3709 2526
rect 3836 2523 3845 2526
rect 3908 2523 3917 2526
rect 3962 2523 3972 2526
rect 4004 2523 4013 2526
rect 14 2467 4211 2473
rect 2642 2443 2685 2446
rect 2012 2433 2061 2436
rect 1212 2423 1261 2426
rect 2018 2423 2028 2426
rect 2090 2423 2109 2426
rect 3026 2416 3029 2425
rect 3138 2416 3141 2425
rect 132 2413 141 2416
rect 180 2413 189 2416
rect 282 2406 285 2416
rect 172 2403 197 2406
rect 236 2403 245 2406
rect 268 2403 308 2406
rect 338 2405 341 2416
rect 346 2413 356 2416
rect 378 2413 388 2416
rect 434 2413 444 2416
rect 506 2413 540 2416
rect 666 2413 692 2416
rect 722 2413 765 2416
rect 820 2413 829 2416
rect 908 2413 925 2416
rect 962 2406 965 2414
rect 1058 2413 1076 2416
rect 1122 2413 1196 2416
rect 1348 2413 1357 2416
rect 1682 2413 1700 2416
rect 1738 2413 1748 2416
rect 364 2403 389 2406
rect 412 2403 429 2406
rect 458 2403 468 2406
rect 484 2403 532 2406
rect 564 2403 581 2406
rect 660 2403 677 2406
rect 754 2403 764 2406
rect 900 2403 965 2406
rect 988 2403 1005 2406
rect 1066 2403 1084 2406
rect 1100 2403 1117 2406
rect 1138 2403 1188 2406
rect 1212 2403 1269 2406
rect 1276 2403 1293 2406
rect 1298 2403 1324 2406
rect 1442 2403 1452 2406
rect 1580 2403 1589 2406
rect 1594 2403 1612 2406
rect 1676 2403 1693 2406
rect 1730 2403 1756 2406
rect 1778 2403 1781 2414
rect 1866 2413 1884 2416
rect 1948 2413 1965 2416
rect 2084 2413 2109 2416
rect 2172 2413 2189 2416
rect 2202 2413 2228 2416
rect 2258 2413 2284 2416
rect 2340 2413 2357 2416
rect 2402 2413 2420 2416
rect 2556 2413 2581 2416
rect 2106 2406 2109 2413
rect 2202 2406 2205 2413
rect 1866 2403 1892 2406
rect 1908 2403 1925 2406
rect 1930 2403 1940 2406
rect 2050 2403 2068 2406
rect 2106 2403 2117 2406
rect 2122 2403 2148 2406
rect 2164 2403 2205 2406
rect 2578 2406 2581 2413
rect 2626 2407 2629 2416
rect 2634 2413 2701 2416
rect 2698 2407 2701 2413
rect 2738 2413 2788 2416
rect 2834 2413 2844 2416
rect 2738 2406 2741 2413
rect 3002 2407 3005 2416
rect 3012 2413 3029 2416
rect 3074 2413 3084 2416
rect 3138 2413 3156 2416
rect 3218 2407 3221 2416
rect 3252 2413 3261 2416
rect 3418 2407 3421 2416
rect 3538 2407 3541 2436
rect 3562 2416 3565 2425
rect 3618 2416 3621 2425
rect 3548 2413 3565 2416
rect 3604 2413 3621 2416
rect 3690 2407 3693 2416
rect 3732 2413 3757 2416
rect 3826 2413 3836 2416
rect 3842 2413 3852 2416
rect 3890 2406 3893 2414
rect 3916 2413 3933 2416
rect 4098 2413 4116 2416
rect 2578 2403 2596 2406
rect 2732 2403 2741 2406
rect 3162 2403 3172 2406
rect 3850 2403 3860 2406
rect 3882 2403 3893 2406
rect 3922 2403 3940 2406
rect 1922 2396 1925 2403
rect 882 2393 892 2396
rect 1218 2393 1268 2396
rect 1922 2393 1933 2396
rect 2578 2393 2581 2403
rect 2106 2383 2125 2386
rect 38 2367 4187 2373
rect 922 2343 980 2346
rect 1258 2343 1277 2346
rect 2610 2343 2637 2346
rect 1274 2336 1277 2343
rect 202 2325 205 2336
rect 220 2333 245 2336
rect 274 2333 292 2336
rect 340 2333 349 2336
rect 378 2333 388 2336
rect 628 2333 669 2336
rect 732 2333 773 2336
rect 786 2333 796 2336
rect 818 2333 853 2336
rect 866 2333 892 2336
rect 916 2333 933 2336
rect 954 2333 988 2336
rect 1034 2333 1068 2336
rect 1106 2333 1172 2336
rect 1196 2333 1269 2336
rect 1274 2333 1284 2336
rect 1306 2326 1309 2335
rect 1362 2333 1372 2336
rect 1434 2333 1444 2336
rect 1500 2333 1525 2336
rect 1540 2333 1565 2336
rect 1836 2333 1877 2336
rect 276 2323 285 2326
rect 322 2323 332 2326
rect 338 2323 348 2326
rect 380 2323 396 2326
rect 556 2323 581 2326
rect 620 2323 629 2326
rect 658 2323 668 2326
rect 754 2323 788 2326
rect 826 2323 869 2326
rect 874 2323 900 2326
rect 996 2323 1061 2326
rect 1066 2323 1076 2326
rect 1090 2323 1165 2326
rect 1188 2323 1221 2326
rect 1306 2323 1380 2326
rect 1386 2323 1412 2326
rect 1466 2323 1484 2326
rect 1514 2323 1532 2326
rect 1538 2323 1564 2326
rect 1596 2323 1621 2326
rect 1660 2323 1669 2326
rect 1764 2323 1781 2326
rect 1866 2323 1876 2326
rect 1906 2325 1909 2336
rect 1956 2333 1965 2336
rect 2322 2333 2340 2336
rect 2356 2333 2420 2336
rect 2452 2333 2461 2336
rect 2586 2333 2613 2336
rect 2650 2333 2660 2336
rect 2692 2333 2749 2336
rect 2754 2333 2772 2336
rect 2818 2333 2828 2336
rect 3770 2333 3788 2336
rect 3812 2333 3829 2336
rect 3948 2333 3957 2336
rect 1962 2323 1972 2326
rect 2066 2323 2092 2326
rect 2250 2323 2268 2326
rect 2444 2323 2477 2326
rect 2506 2323 2556 2326
rect 2698 2323 2764 2326
rect 2842 2323 2845 2333
rect 2890 2323 2916 2326
rect 2970 2323 2980 2326
rect 3026 2323 3036 2326
rect 3058 2323 3068 2326
rect 3108 2323 3125 2326
rect 3258 2323 3284 2326
rect 3322 2323 3332 2326
rect 3362 2323 3388 2326
rect 3458 2323 3484 2326
rect 3522 2323 3540 2326
rect 3684 2323 3709 2326
rect 3804 2323 3813 2326
rect 3954 2323 3964 2326
rect 3994 2323 4020 2326
rect 4090 2323 4116 2326
rect 916 2313 973 2316
rect 1092 2313 1157 2316
rect 1210 2313 1284 2316
rect 1866 2313 1869 2323
rect 2066 2313 2085 2316
rect 834 2286 837 2296
rect 834 2283 853 2286
rect 14 2267 4211 2273
rect 882 2253 909 2256
rect 722 2216 725 2226
rect 108 2213 117 2216
rect 204 2213 213 2216
rect 260 2213 269 2216
rect 316 2213 325 2216
rect 420 2213 429 2216
rect 476 2213 493 2216
rect 578 2213 596 2216
rect 610 2213 636 2216
rect 378 2203 396 2206
rect 418 2203 428 2206
rect 442 2203 460 2206
rect 482 2203 500 2206
rect 522 2203 532 2206
rect 604 2203 637 2206
rect 666 2203 669 2214
rect 674 2205 677 2216
rect 684 2213 701 2216
rect 722 2213 733 2216
rect 740 2213 757 2216
rect 796 2213 837 2216
rect 730 2205 733 2213
rect 842 2206 845 2214
rect 876 2213 901 2216
rect 906 2206 909 2253
rect 2682 2216 2685 2226
rect 2714 2216 2717 2236
rect 788 2203 845 2206
rect 868 2203 909 2206
rect 938 2203 941 2214
rect 1028 2213 1037 2216
rect 1082 2213 1108 2216
rect 1332 2213 1349 2216
rect 1402 2213 1420 2216
rect 1492 2213 1517 2216
rect 1548 2213 1581 2216
rect 1642 2213 1660 2216
rect 1738 2213 1748 2216
rect 1914 2213 1948 2216
rect 2042 2213 2076 2216
rect 2148 2213 2204 2216
rect 2300 2213 2325 2216
rect 2436 2213 2461 2216
rect 2498 2213 2524 2216
rect 2586 2213 2596 2216
rect 2676 2213 2701 2216
rect 2714 2213 2724 2216
rect 970 2203 1020 2206
rect 1346 2205 1349 2213
rect 2314 2206 2317 2213
rect 1570 2203 1596 2206
rect 1626 2203 1668 2206
rect 1690 2203 1700 2206
rect 1714 2203 1756 2206
rect 1778 2203 1812 2206
rect 1850 2203 1876 2206
rect 1892 2203 1917 2206
rect 1938 2203 1956 2206
rect 1978 2203 2020 2206
rect 2084 2203 2117 2206
rect 2250 2203 2276 2206
rect 2314 2203 2364 2206
rect 2380 2203 2397 2206
rect 2418 2203 2428 2206
rect 2562 2203 2588 2206
rect 2602 2203 2652 2206
rect 2674 2203 2732 2206
rect 2754 2203 2757 2214
rect 2762 2205 2765 2216
rect 2810 2213 2836 2216
rect 3066 2213 3084 2216
rect 3140 2213 3149 2216
rect 3196 2213 3205 2216
rect 3308 2213 3325 2216
rect 3202 2205 3205 2213
rect 3322 2205 3325 2213
rect 3362 2203 3365 2214
rect 3412 2213 3437 2216
rect 3490 2203 3493 2214
rect 3618 2203 3621 2214
rect 3756 2213 3765 2216
rect 3812 2213 3837 2216
rect 3868 2213 3877 2216
rect 3924 2213 3933 2216
rect 4116 2213 4125 2216
rect 3762 2205 3765 2213
rect 3874 2205 3877 2213
rect 4122 2205 4125 2213
rect 746 2193 780 2196
rect 978 2193 997 2196
rect 38 2167 4187 2173
rect 874 2143 916 2146
rect 2442 2143 2476 2146
rect 2682 2143 2708 2146
rect 3202 2136 3205 2146
rect 132 2133 149 2136
rect 180 2133 204 2136
rect 290 2133 300 2136
rect 362 2133 396 2136
rect 626 2133 660 2136
rect 676 2133 685 2136
rect 826 2133 836 2136
rect 860 2133 869 2136
rect 924 2133 989 2136
rect 1012 2133 1037 2136
rect 1050 2133 1076 2136
rect 1154 2133 1164 2136
rect 1188 2133 1245 2136
rect 826 2126 829 2133
rect 114 2123 124 2126
rect 138 2123 156 2126
rect 188 2123 197 2126
rect 202 2123 212 2126
rect 298 2123 308 2126
rect 356 2123 381 2126
rect 556 2123 581 2126
rect 612 2123 637 2126
rect 642 2123 652 2126
rect 812 2123 829 2126
rect 834 2123 844 2126
rect 866 2123 909 2126
rect 932 2123 981 2126
rect 986 2125 989 2133
rect 1250 2126 1253 2135
rect 1284 2133 1348 2136
rect 1380 2133 1389 2136
rect 1516 2133 1557 2136
rect 1572 2133 1605 2136
rect 1020 2123 1053 2126
rect 1066 2123 1084 2126
rect 1180 2123 1213 2126
rect 1226 2123 1253 2126
rect 1594 2123 1604 2126
rect 1634 2125 1637 2136
rect 2114 2133 2124 2136
rect 2154 2133 2172 2136
rect 2330 2133 2340 2136
rect 2402 2133 2412 2136
rect 2428 2133 2469 2136
rect 2490 2133 2524 2136
rect 1706 2123 1716 2126
rect 1946 2123 1972 2126
rect 2100 2123 2109 2126
rect 2148 2123 2165 2126
rect 2180 2123 2189 2126
rect 2226 2123 2252 2126
rect 2290 2123 2300 2126
rect 2338 2123 2348 2126
rect 2466 2123 2469 2133
rect 2594 2126 2597 2136
rect 2626 2133 2668 2136
rect 2716 2133 2749 2136
rect 2844 2133 2869 2136
rect 2882 2133 2892 2136
rect 2956 2133 2988 2136
rect 3052 2133 3061 2136
rect 3108 2133 3125 2136
rect 3202 2133 3220 2136
rect 3266 2133 3284 2136
rect 3330 2126 3333 2134
rect 3466 2133 3476 2136
rect 3522 2126 3525 2134
rect 3554 2126 3557 2134
rect 3716 2133 3724 2136
rect 2554 2125 2597 2126
rect 2554 2123 2596 2125
rect 2628 2123 2645 2126
rect 2676 2123 2693 2126
rect 2786 2123 2820 2126
rect 2858 2123 2917 2126
rect 2948 2123 2973 2126
rect 2978 2123 2996 2126
rect 3026 2123 3044 2126
rect 3218 2123 3228 2126
rect 3258 2123 3292 2126
rect 3330 2123 3356 2126
rect 3386 2123 3412 2126
rect 3522 2123 3541 2126
rect 3554 2123 3573 2126
rect 3682 2123 3692 2126
rect 3722 2123 3732 2126
rect 3770 2125 3773 2136
rect 3796 2133 3813 2136
rect 4002 2133 4012 2136
rect 3804 2123 3812 2126
rect 3850 2123 3860 2126
rect 3890 2123 3924 2126
rect 3954 2123 3972 2126
rect 3978 2123 4020 2126
rect 860 2113 901 2116
rect 1100 2113 1125 2116
rect 2730 2113 2756 2116
rect 2780 2113 2789 2116
rect 3172 2113 3181 2116
rect 3196 2113 3205 2116
rect 3562 2113 3596 2116
rect 3754 2113 3764 2116
rect 14 2067 4211 2073
rect 1972 2033 1997 2036
rect 3114 2033 3156 2036
rect 724 2023 757 2026
rect 1162 2023 1188 2026
rect 1914 2023 1964 2026
rect 1988 2023 2005 2026
rect 2994 2023 3028 2026
rect 3052 2023 3084 2026
rect 3108 2023 3133 2026
rect 3164 2023 3181 2026
rect 3434 2023 3452 2026
rect 3780 2023 3797 2026
rect 2002 2016 2005 2023
rect 108 2013 117 2016
rect 394 2013 421 2016
rect 426 2013 436 2016
rect 468 2013 485 2016
rect 554 2013 580 2016
rect 652 2013 693 2016
rect 738 2013 772 2016
rect 418 2006 421 2013
rect 858 2006 861 2014
rect 180 2003 189 2006
rect 194 2003 204 2006
rect 338 2003 356 2006
rect 388 2003 413 2006
rect 418 2003 444 2006
rect 466 2003 508 2006
rect 746 2003 780 2006
rect 802 2003 861 2006
rect 884 2003 925 2006
rect 970 2003 973 2014
rect 1004 2013 1077 2016
rect 1204 2013 1213 2016
rect 1314 2013 1364 2016
rect 1370 2013 1380 2016
rect 1410 2013 1436 2016
rect 1492 2013 1500 2016
rect 1556 2013 1565 2016
rect 1722 2013 1748 2016
rect 1812 2013 1884 2016
rect 2002 2013 2020 2016
rect 2076 2013 2085 2016
rect 996 2003 1013 2006
rect 1018 2003 1084 2006
rect 1108 2003 1117 2006
rect 1122 2003 1188 2006
rect 1212 2003 1277 2006
rect 1316 2003 1357 2006
rect 1370 2005 1373 2013
rect 1658 2003 1684 2006
rect 1770 2003 1788 2006
rect 1826 2003 1876 2006
rect 1908 2003 1933 2006
rect 2028 2003 2045 2006
rect 2090 2003 2108 2006
rect 2210 2003 2220 2006
rect 2252 2003 2261 2006
rect 2274 2003 2277 2014
rect 2468 2013 2477 2016
rect 2538 2013 2548 2016
rect 2474 2005 2477 2013
rect 2524 2003 2549 2006
rect 2556 2003 2565 2006
rect 2602 2005 2605 2016
rect 2690 2013 2700 2016
rect 2764 2013 2821 2016
rect 2972 2013 2997 2016
rect 2930 2003 2948 2006
rect 3042 2003 3045 2014
rect 3244 2013 3253 2016
rect 3266 2013 3276 2016
rect 3412 2013 3421 2016
rect 3204 2003 3213 2006
rect 3236 2003 3261 2006
rect 3418 2005 3421 2013
rect 3498 2003 3501 2014
rect 3538 2005 3541 2016
rect 3668 2013 3693 2016
rect 3786 2013 3812 2016
rect 3850 2013 3860 2016
rect 3980 2013 3989 2016
rect 4002 2013 4012 2016
rect 3690 2005 3693 2013
rect 3802 2003 3820 2006
rect 3836 2003 3845 2006
rect 3986 2005 3989 2013
rect 626 1993 636 1996
rect 1658 1993 1677 1996
rect 38 1967 4187 1973
rect 722 1943 756 1946
rect 770 1943 796 1946
rect 826 1943 852 1946
rect 180 1933 189 1936
rect 458 1933 484 1936
rect 516 1933 525 1936
rect 652 1933 677 1936
rect 764 1933 797 1936
rect 804 1933 837 1936
rect 866 1933 884 1936
rect 900 1933 957 1936
rect 980 1933 1029 1936
rect 1034 1933 1052 1936
rect 1250 1926 1253 1934
rect 1282 1933 1292 1936
rect 108 1923 125 1926
rect 260 1923 269 1926
rect 356 1923 365 1926
rect 444 1923 461 1926
rect 564 1923 589 1926
rect 626 1923 644 1926
rect 658 1923 676 1926
rect 708 1923 725 1926
rect 772 1923 789 1926
rect 812 1923 853 1926
rect 988 1923 1005 1926
rect 1084 1923 1101 1926
rect 1180 1923 1189 1926
rect 1236 1923 1253 1926
rect 1260 1923 1285 1926
rect 1322 1923 1325 1934
rect 1330 1933 1356 1936
rect 1402 1926 1405 1934
rect 1524 1933 1533 1936
rect 1620 1933 1629 1936
rect 1666 1933 1676 1936
rect 1708 1933 1749 1936
rect 1900 1933 1909 1936
rect 1994 1933 2004 1936
rect 2370 1926 2373 1934
rect 2396 1933 2429 1936
rect 2554 1926 2557 1934
rect 2580 1933 2621 1936
rect 2650 1926 2653 1934
rect 2772 1933 2781 1936
rect 2826 1933 2844 1936
rect 2884 1933 2933 1936
rect 2972 1933 2981 1936
rect 3010 1926 3013 1934
rect 3314 1926 3317 1934
rect 3386 1933 3404 1936
rect 3420 1933 3429 1936
rect 3540 1933 3557 1936
rect 3580 1933 3589 1936
rect 3762 1926 3765 1934
rect 3778 1933 3796 1936
rect 3812 1933 3829 1936
rect 3868 1933 3877 1936
rect 4020 1933 4037 1936
rect 3778 1926 3781 1933
rect 1386 1923 1396 1926
rect 1402 1923 1412 1926
rect 1442 1923 1468 1926
rect 1580 1923 1604 1926
rect 1700 1923 1709 1926
rect 1874 1923 1884 1926
rect 1994 1923 2012 1926
rect 2292 1923 2301 1926
rect 2348 1923 2373 1926
rect 2524 1923 2557 1926
rect 2602 1923 2621 1926
rect 2650 1923 2668 1926
rect 2892 1923 2925 1926
rect 2970 1923 3004 1926
rect 3010 1923 3036 1926
rect 3066 1923 3092 1926
rect 1994 1916 1997 1923
rect 1938 1913 1948 1916
rect 1972 1913 1997 1916
rect 2044 1913 2053 1916
rect 2058 1913 2076 1916
rect 2602 1913 2628 1916
rect 2812 1913 2829 1916
rect 3138 1913 3148 1916
rect 2050 1906 2053 1913
rect 3162 1906 3165 1925
rect 3244 1923 3269 1926
rect 3300 1923 3317 1926
rect 3324 1923 3349 1926
rect 3506 1923 3516 1926
rect 3546 1923 3572 1926
rect 3692 1923 3717 1926
rect 3748 1923 3765 1926
rect 3772 1923 3781 1926
rect 3978 1923 3996 1926
rect 4026 1923 4044 1926
rect 3172 1913 3205 1916
rect 3458 1913 3476 1916
rect 1956 1903 1989 1906
rect 2050 1903 2061 1906
rect 2066 1903 2092 1906
rect 3162 1903 3189 1906
rect 14 1867 4211 1873
rect 858 1853 909 1856
rect 2690 1853 2709 1856
rect 2730 1833 2804 1836
rect 2874 1833 2885 1836
rect 772 1823 805 1826
rect 836 1823 901 1826
rect 1066 1823 1116 1826
rect 1162 1823 1189 1826
rect 2788 1823 2797 1826
rect 2818 1823 2860 1826
rect 108 1813 117 1816
rect 170 1813 188 1816
rect 202 1813 212 1816
rect 244 1813 253 1816
rect 266 1813 284 1816
rect 290 1813 316 1816
rect 362 1813 380 1816
rect 386 1813 404 1816
rect 492 1813 509 1816
rect 556 1813 581 1816
rect 626 1813 636 1816
rect 658 1813 668 1816
rect 700 1813 725 1816
rect 794 1813 820 1816
rect 196 1803 213 1806
rect 236 1803 261 1806
rect 292 1803 317 1806
rect 388 1803 405 1806
rect 442 1803 468 1806
rect 644 1803 669 1806
rect 706 1803 748 1806
rect 772 1803 789 1806
rect 794 1803 812 1806
rect 836 1803 853 1806
rect 914 1803 917 1814
rect 996 1813 1021 1816
rect 1052 1813 1061 1816
rect 1132 1813 1173 1816
rect 1220 1813 1261 1816
rect 1300 1813 1317 1816
rect 1410 1813 1444 1816
rect 1514 1813 1548 1816
rect 1634 1813 1644 1816
rect 1722 1813 1756 1816
rect 1844 1813 1853 1816
rect 1962 1813 1988 1816
rect 2148 1813 2157 1816
rect 2250 1813 2260 1816
rect 2298 1813 2308 1816
rect 2314 1813 2324 1816
rect 2356 1813 2365 1816
rect 2474 1813 2524 1816
rect 2874 1815 2877 1833
rect 2884 1823 2893 1826
rect 3266 1823 3292 1826
rect 3316 1823 3341 1826
rect 1514 1806 1517 1813
rect 1066 1803 1116 1806
rect 1140 1803 1189 1806
rect 1234 1803 1261 1806
rect 1362 1803 1372 1806
rect 1404 1803 1413 1806
rect 1452 1803 1485 1806
rect 1508 1803 1517 1806
rect 1572 1803 1581 1806
rect 1700 1803 1749 1806
rect 1754 1803 1764 1806
rect 1780 1803 1797 1806
rect 1836 1803 1869 1806
rect 1898 1803 1916 1806
rect 2052 1803 2077 1806
rect 2090 1803 2100 1806
rect 2114 1803 2124 1806
rect 2140 1803 2188 1806
rect 2212 1803 2221 1806
rect 2276 1803 2293 1806
rect 2316 1803 2325 1806
rect 2386 1803 2404 1806
rect 2428 1803 2453 1806
rect 2514 1803 2532 1806
rect 2548 1803 2636 1806
rect 2658 1803 2661 1814
rect 2666 1803 2716 1806
rect 2794 1803 2797 1814
rect 2922 1813 2932 1816
rect 2938 1813 2956 1816
rect 2986 1813 3012 1816
rect 3084 1813 3109 1816
rect 3140 1813 3157 1816
rect 3162 1813 3172 1816
rect 3330 1813 3356 1816
rect 2938 1805 2941 1813
rect 3380 1803 3389 1806
rect 3562 1803 3565 1814
rect 3610 1813 3636 1816
rect 3756 1803 3773 1806
rect 3812 1803 3845 1806
rect 3890 1803 3908 1806
rect 3930 1803 3933 1814
rect 3978 1813 3996 1816
rect 3948 1803 3973 1806
rect 1066 1793 1085 1796
rect 1410 1793 1413 1803
rect 1810 1793 1828 1796
rect 2026 1793 2044 1796
rect 38 1767 4187 1773
rect 1714 1743 1724 1746
rect 1738 1743 1780 1746
rect 1930 1736 1933 1746
rect 1986 1743 2012 1746
rect 2114 1743 2133 1746
rect 3130 1743 3165 1746
rect 3834 1743 3845 1746
rect 3938 1743 3949 1746
rect 3834 1736 3837 1743
rect 228 1733 237 1736
rect 380 1733 389 1736
rect 570 1726 573 1735
rect 818 1733 828 1736
rect 844 1733 876 1736
rect 1066 1733 1076 1736
rect 1092 1733 1141 1736
rect 1178 1733 1212 1736
rect 1268 1733 1293 1736
rect 1348 1733 1357 1736
rect 1412 1733 1429 1736
rect 1586 1733 1628 1736
rect 1642 1733 1668 1736
rect 1692 1733 1709 1736
rect 1732 1733 1781 1736
rect 1794 1733 1828 1736
rect 1858 1733 1892 1736
rect 1908 1733 1956 1736
rect 1980 1733 2005 1736
rect 2020 1733 2045 1736
rect 2066 1733 2076 1736
rect 2092 1733 2125 1736
rect 2130 1733 2140 1736
rect 2276 1733 2317 1736
rect 2346 1733 2373 1736
rect 2500 1733 2517 1736
rect 2522 1733 2540 1736
rect 2556 1733 2588 1736
rect 2668 1733 2701 1736
rect 2948 1733 3012 1736
rect 3044 1733 3077 1736
rect 3154 1733 3172 1736
rect 3194 1733 3228 1736
rect 3242 1733 3260 1736
rect 3290 1733 3308 1736
rect 3388 1733 3397 1736
rect 3428 1733 3437 1736
rect 116 1723 141 1726
rect 186 1723 220 1726
rect 226 1723 236 1726
rect 308 1723 333 1726
rect 532 1723 573 1726
rect 692 1723 709 1726
rect 754 1723 796 1726
rect 906 1723 964 1726
rect 1026 1723 1068 1726
rect 1138 1723 1164 1726
rect 1330 1723 1340 1726
rect 1346 1723 1372 1726
rect 1378 1723 1404 1726
rect 1530 1723 1540 1726
rect 1588 1723 1605 1726
rect 1658 1723 1676 1726
rect 1740 1723 1773 1726
rect 1802 1723 1836 1726
rect 1866 1723 1884 1726
rect 1916 1723 1933 1726
rect 2028 1723 2061 1726
rect 2100 1723 2109 1726
rect 2148 1723 2157 1726
rect 2194 1723 2220 1726
rect 2258 1723 2268 1726
rect 2306 1723 2316 1726
rect 2348 1723 2365 1726
rect 900 1713 957 1716
rect 1692 1713 1717 1716
rect 1852 1713 1869 1716
rect 1874 1703 1877 1723
rect 2370 1716 2373 1733
rect 3290 1726 3293 1733
rect 3762 1726 3765 1735
rect 3778 1733 3788 1736
rect 3820 1733 3837 1736
rect 3842 1733 3860 1736
rect 2412 1723 2437 1726
rect 2474 1723 2492 1726
rect 2498 1723 2532 1726
rect 2586 1723 2596 1726
rect 2634 1723 2652 1726
rect 2698 1723 2716 1726
rect 1980 1713 1989 1716
rect 2362 1713 2373 1716
rect 2746 1713 2756 1716
rect 2770 1706 2773 1725
rect 2786 1723 2805 1726
rect 2940 1723 2965 1726
rect 2994 1723 3020 1726
rect 3050 1723 3100 1726
rect 3130 1723 3180 1726
rect 3276 1723 3293 1726
rect 3330 1723 3364 1726
rect 3402 1723 3420 1726
rect 3700 1723 3725 1726
rect 3756 1723 3765 1726
rect 3772 1723 3781 1726
rect 3812 1723 3868 1726
rect 2802 1716 2805 1723
rect 3938 1716 3941 1743
rect 3946 1733 3964 1736
rect 3996 1733 4021 1736
rect 4122 1723 4140 1726
rect 2780 1713 2797 1716
rect 2802 1713 2820 1716
rect 3434 1713 3444 1716
rect 3938 1713 3949 1716
rect 2770 1703 2805 1706
rect 2828 1703 2837 1706
rect 14 1667 4211 1673
rect 1164 1623 1173 1626
rect 1772 1623 1789 1626
rect 2130 1623 2156 1626
rect 2452 1623 2461 1626
rect 3250 1623 3260 1626
rect 3522 1623 3612 1626
rect 3636 1623 3669 1626
rect 108 1613 117 1616
rect 372 1613 389 1616
rect 442 1613 460 1616
rect 548 1613 573 1616
rect 626 1613 660 1616
rect 180 1603 189 1606
rect 332 1603 341 1606
rect 380 1603 412 1606
rect 428 1603 468 1606
rect 484 1603 509 1606
rect 620 1603 661 1606
rect 690 1603 693 1614
rect 770 1613 796 1616
rect 828 1613 853 1616
rect 882 1613 892 1616
rect 972 1613 997 1616
rect 1028 1613 1069 1616
rect 1084 1613 1117 1616
rect 1138 1613 1148 1616
rect 1162 1613 1212 1616
rect 1274 1613 1284 1616
rect 1476 1613 1501 1616
rect 740 1603 757 1606
rect 820 1603 877 1606
rect 890 1603 900 1606
rect 916 1603 933 1606
rect 946 1603 964 1606
rect 1020 1603 1029 1606
rect 1092 1603 1109 1606
rect 1130 1603 1140 1606
rect 1178 1603 1204 1606
rect 1266 1603 1276 1606
rect 1538 1603 1541 1614
rect 1572 1613 1612 1616
rect 1644 1613 1677 1616
rect 1714 1613 1756 1616
rect 1820 1613 1836 1616
rect 1868 1613 1893 1616
rect 2036 1613 2053 1616
rect 1578 1603 1620 1606
rect 1730 1603 1748 1606
rect 1778 1603 1804 1606
rect 1876 1603 1901 1606
rect 1924 1603 1941 1606
rect 2050 1605 2053 1613
rect 2122 1606 2125 1614
rect 2172 1613 2189 1616
rect 2228 1613 2253 1616
rect 2324 1613 2349 1616
rect 2386 1613 2396 1616
rect 2402 1613 2436 1616
rect 2450 1613 2485 1616
rect 2588 1613 2605 1616
rect 2692 1613 2709 1616
rect 2746 1613 2772 1616
rect 2898 1613 2924 1616
rect 3092 1613 3109 1616
rect 3172 1613 3213 1616
rect 3420 1613 3429 1616
rect 3458 1613 3484 1616
rect 3642 1613 3684 1616
rect 3714 1613 3732 1616
rect 3796 1613 3813 1616
rect 3852 1613 3861 1616
rect 3868 1613 3885 1616
rect 3890 1613 3908 1616
rect 2076 1603 2085 1606
rect 2122 1603 2156 1606
rect 2404 1603 2421 1606
rect 2450 1605 2453 1613
rect 2602 1606 2605 1613
rect 2466 1603 2500 1606
rect 2516 1603 2549 1606
rect 2602 1603 2628 1606
rect 2650 1603 2684 1606
rect 2948 1603 2997 1606
rect 3106 1605 3109 1613
rect 3130 1603 3148 1606
rect 3164 1603 3205 1606
rect 3244 1603 3253 1606
rect 3426 1605 3429 1613
rect 3508 1603 3533 1606
rect 3858 1605 3861 1613
rect 3874 1606 3877 1613
rect 3874 1603 3916 1606
rect 3938 1603 3941 1614
rect 4132 1613 4141 1616
rect 3946 1603 3972 1606
rect 4138 1605 4141 1613
rect 706 1593 732 1596
rect 978 1593 1012 1596
rect 1650 1593 1692 1596
rect 2090 1593 2108 1596
rect 38 1567 4187 1573
rect 754 1543 764 1546
rect 922 1543 940 1546
rect 180 1533 213 1536
rect 218 1533 228 1536
rect 404 1533 437 1536
rect 490 1533 500 1536
rect 610 1533 620 1536
rect 642 1533 652 1536
rect 682 1533 716 1536
rect 740 1533 749 1536
rect 812 1533 821 1536
rect 842 1533 852 1536
rect 108 1523 117 1526
rect 194 1523 220 1526
rect 258 1523 268 1526
rect 332 1523 357 1526
rect 410 1523 436 1526
rect 468 1523 485 1526
rect 538 1523 548 1526
rect 602 1523 612 1526
rect 660 1523 677 1526
rect 706 1523 724 1526
rect 780 1523 789 1526
rect 826 1523 844 1526
rect 882 1525 885 1536
rect 908 1533 941 1536
rect 948 1533 965 1536
rect 1066 1533 1092 1536
rect 1116 1533 1165 1536
rect 1194 1526 1197 1535
rect 1228 1533 1245 1536
rect 1362 1526 1365 1535
rect 1378 1533 1396 1536
rect 1428 1533 1437 1536
rect 1548 1533 1557 1536
rect 1562 1533 1580 1536
rect 1596 1533 1621 1536
rect 1634 1533 1644 1536
rect 1668 1533 1693 1536
rect 1794 1533 1812 1536
rect 1866 1533 1876 1536
rect 1900 1533 1909 1536
rect 1922 1533 1932 1536
rect 2060 1533 2069 1536
rect 2082 1533 2092 1536
rect 2116 1533 2133 1536
rect 2156 1533 2181 1536
rect 2212 1533 2229 1536
rect 2234 1533 2252 1536
rect 2282 1533 2308 1536
rect 2332 1533 2341 1536
rect 2346 1533 2364 1536
rect 2388 1533 2413 1536
rect 2452 1533 2461 1536
rect 2516 1533 2541 1536
rect 2572 1533 2597 1536
rect 2628 1533 2653 1536
rect 2690 1533 2716 1536
rect 2746 1533 2756 1536
rect 2818 1533 2852 1536
rect 1562 1526 1565 1533
rect 3010 1526 3013 1534
rect 3074 1533 3100 1536
rect 916 1523 933 1526
rect 956 1523 965 1526
rect 1004 1523 1013 1526
rect 1108 1523 1117 1526
rect 1154 1516 1157 1526
rect 1194 1523 1261 1526
rect 1300 1523 1317 1526
rect 1356 1523 1365 1526
rect 1420 1523 1429 1526
rect 1476 1523 1501 1526
rect 1546 1523 1565 1526
rect 1634 1523 1652 1526
rect 1722 1523 1772 1526
rect 1828 1523 1844 1526
rect 1898 1523 1940 1526
rect 1956 1523 1973 1526
rect 1996 1523 2044 1526
rect 2066 1523 2100 1526
rect 2130 1523 2140 1526
rect 2162 1523 2196 1526
rect 2210 1523 2260 1526
rect 2274 1523 2316 1526
rect 2330 1523 2372 1526
rect 2402 1523 2436 1526
rect 2450 1523 2500 1526
rect 2514 1523 2556 1526
rect 1970 1516 1973 1523
rect 740 1513 757 1516
rect 812 1513 837 1516
rect 1122 1513 1172 1516
rect 1668 1513 1693 1516
rect 1866 1513 1876 1516
rect 1970 1513 1980 1516
rect 2212 1513 2229 1516
rect 2572 1513 2604 1516
rect 2634 1513 2660 1516
rect 2674 1506 2677 1525
rect 2876 1523 2885 1526
rect 2996 1523 3013 1526
rect 2684 1513 2717 1516
rect 3026 1513 3044 1516
rect 3058 1506 3061 1525
rect 3116 1523 3124 1526
rect 3146 1525 3149 1536
rect 3172 1533 3181 1536
rect 3220 1533 3229 1536
rect 3380 1533 3397 1536
rect 3466 1533 3540 1536
rect 3562 1533 3580 1536
rect 3644 1533 3661 1536
rect 3708 1533 3717 1536
rect 3964 1533 3981 1536
rect 3242 1523 3252 1526
rect 3282 1523 3308 1526
rect 3418 1523 3444 1526
rect 3466 1523 3588 1526
rect 3626 1523 3636 1526
rect 3642 1523 3684 1526
rect 3770 1523 3796 1526
rect 3834 1523 3844 1526
rect 3874 1523 3900 1526
rect 3986 1523 3989 1534
rect 4122 1526 4125 1534
rect 4116 1523 4125 1526
rect 3068 1513 3077 1516
rect 2674 1503 2701 1506
rect 3058 1503 3093 1506
rect 14 1467 4211 1473
rect 2786 1433 2797 1436
rect 764 1423 797 1426
rect 108 1413 133 1416
rect 164 1413 189 1416
rect 194 1413 204 1416
rect 236 1413 253 1416
rect 292 1413 317 1416
rect 362 1413 396 1416
rect 428 1413 445 1416
rect 540 1413 581 1416
rect 738 1413 748 1416
rect 820 1413 829 1416
rect 884 1413 909 1416
rect 946 1413 972 1416
rect 1034 1413 1037 1424
rect 1090 1423 1116 1426
rect 1722 1423 1732 1426
rect 1812 1423 1821 1426
rect 1188 1413 1213 1416
rect 1300 1413 1349 1416
rect 1388 1413 1429 1416
rect 1524 1413 1541 1416
rect 1572 1413 1581 1416
rect 1700 1413 1725 1416
rect 186 1406 189 1413
rect 186 1403 212 1406
rect 228 1403 237 1406
rect 364 1403 397 1406
rect 578 1405 581 1413
rect 612 1403 629 1406
rect 764 1403 773 1406
rect 802 1403 812 1406
rect 954 1403 964 1406
rect 978 1403 1012 1406
rect 1082 1403 1116 1406
rect 1140 1403 1149 1406
rect 1314 1403 1364 1406
rect 1396 1403 1429 1406
rect 1538 1405 1541 1413
rect 1818 1406 1821 1423
rect 2770 1423 2781 1426
rect 1860 1413 1877 1416
rect 1964 1413 1989 1416
rect 2020 1413 2029 1416
rect 2076 1413 2093 1416
rect 2132 1413 2141 1416
rect 2148 1413 2165 1416
rect 2170 1413 2196 1416
rect 2340 1413 2349 1416
rect 2372 1413 2428 1416
rect 2458 1413 2492 1416
rect 2498 1413 2509 1416
rect 2514 1413 2540 1416
rect 2570 1413 2588 1416
rect 2652 1413 2677 1416
rect 2708 1413 2717 1416
rect 2724 1413 2733 1416
rect 1682 1403 1692 1406
rect 1706 1403 1732 1406
rect 1762 1403 1788 1406
rect 1818 1403 1844 1406
rect 2026 1405 2029 1413
rect 2138 1405 2141 1413
rect 2178 1403 2188 1406
rect 2220 1403 2229 1406
rect 2346 1405 2349 1413
rect 2506 1406 2509 1413
rect 2394 1403 2420 1406
rect 2506 1403 2532 1406
rect 2596 1403 2613 1406
rect 2714 1405 2717 1413
rect 2770 1406 2773 1423
rect 2786 1413 2789 1433
rect 2794 1413 2812 1416
rect 2866 1413 2876 1416
rect 2996 1413 3005 1416
rect 3012 1413 3021 1416
rect 3060 1413 3069 1416
rect 3116 1413 3125 1416
rect 3138 1413 3172 1416
rect 3202 1413 3228 1416
rect 3234 1413 3292 1416
rect 3298 1413 3348 1416
rect 3378 1413 3396 1416
rect 3460 1413 3485 1416
rect 3516 1413 3525 1416
rect 3602 1413 3620 1416
rect 3626 1413 3644 1416
rect 3698 1413 3732 1416
rect 3770 1413 3805 1416
rect 3842 1413 3884 1416
rect 3930 1413 3940 1416
rect 3994 1413 4012 1416
rect 4042 1413 4084 1416
rect 2764 1403 2773 1406
rect 2778 1403 2804 1406
rect 2818 1403 2868 1406
rect 3002 1405 3005 1413
rect 3122 1405 3125 1413
rect 3146 1403 3164 1406
rect 3236 1403 3245 1406
rect 3330 1403 3340 1406
rect 3378 1403 3388 1406
rect 3522 1405 3525 1413
rect 3628 1403 3637 1406
rect 3684 1403 3717 1406
rect 3756 1403 3789 1406
rect 3844 1403 3869 1406
rect 3964 1403 3981 1406
rect 4036 1403 4069 1406
rect 4092 1403 4117 1406
rect 786 1393 804 1396
rect 2770 1386 2773 1403
rect 4114 1393 4117 1403
rect 2770 1383 2789 1386
rect 38 1367 4187 1373
rect 650 1353 677 1356
rect 754 1353 789 1356
rect 2914 1353 2941 1356
rect 642 1343 684 1346
rect 180 1333 213 1336
rect 308 1333 341 1336
rect 402 1333 428 1336
rect 444 1333 469 1336
rect 628 1333 685 1336
rect 714 1333 724 1336
rect 740 1333 804 1336
rect 834 1333 900 1336
rect 108 1323 133 1326
rect 194 1323 212 1326
rect 244 1323 269 1326
rect 274 1323 284 1326
rect 316 1323 341 1326
rect 386 1323 420 1326
rect 490 1323 516 1326
rect 578 1323 604 1326
rect 636 1323 645 1326
rect 700 1323 709 1326
rect 786 1323 812 1326
rect 826 1323 892 1326
rect 922 1325 925 1336
rect 930 1333 996 1336
rect 1020 1333 1029 1336
rect 1034 1333 1108 1336
rect 1132 1333 1141 1336
rect 1154 1326 1157 1335
rect 1274 1333 1308 1336
rect 1340 1333 1373 1336
rect 1490 1326 1493 1335
rect 1554 1333 1572 1336
rect 1794 1333 1804 1336
rect 1818 1333 1836 1336
rect 1874 1333 1892 1336
rect 1940 1333 1973 1336
rect 2012 1333 2052 1336
rect 2276 1333 2317 1336
rect 2322 1326 2325 1335
rect 2356 1333 2365 1336
rect 2396 1333 2405 1336
rect 2556 1333 2565 1336
rect 3010 1333 3020 1336
rect 1012 1323 1109 1326
rect 1130 1323 1148 1326
rect 1154 1323 1180 1326
rect 1210 1323 1236 1326
rect 1332 1323 1349 1326
rect 1468 1323 1493 1326
rect 1506 1323 1532 1326
rect 1546 1323 1589 1326
rect 1628 1323 1653 1326
rect 1700 1323 1709 1326
rect 1756 1323 1773 1326
rect 1812 1323 1837 1326
rect 1874 1323 1900 1326
rect 1954 1323 1988 1326
rect 2076 1323 2132 1326
rect 2170 1323 2204 1326
rect 2234 1323 2268 1326
rect 2314 1323 2325 1326
rect 2362 1323 2388 1326
rect 2514 1323 2532 1326
rect 2700 1323 2725 1326
rect 2756 1323 2765 1326
rect 2770 1323 2780 1326
rect 2842 1323 2860 1326
rect 2986 1323 3028 1326
rect 3058 1325 3061 1336
rect 3090 1333 3124 1336
rect 3140 1333 3205 1336
rect 3508 1333 3533 1336
rect 3796 1333 3805 1336
rect 3906 1326 3909 1335
rect 3092 1323 3116 1326
rect 3162 1323 3181 1326
rect 3410 1323 3436 1326
rect 3516 1323 3541 1326
rect 3620 1323 3629 1326
rect 3746 1323 3772 1326
rect 3900 1323 3909 1326
rect 3922 1325 3925 1336
rect 3954 1325 3957 1336
rect 3978 1333 3988 1336
rect 4132 1333 4149 1336
rect 828 1313 877 1316
rect 1026 1313 1108 1316
rect 1770 1313 1773 1323
rect 2314 1313 2317 1323
rect 2842 1313 2845 1323
rect 14 1267 4211 1273
rect 106 1216 109 1226
rect 1012 1223 1069 1226
rect 106 1213 124 1216
rect 156 1213 173 1216
rect 196 1213 205 1216
rect 500 1213 517 1216
rect 588 1213 605 1216
rect 706 1213 748 1216
rect 804 1213 829 1216
rect 202 1206 205 1213
rect 148 1203 173 1206
rect 202 1203 213 1206
rect 236 1203 261 1206
rect 514 1205 517 1213
rect 906 1206 909 1216
rect 932 1213 981 1216
rect 1138 1213 1188 1216
rect 1220 1213 1245 1216
rect 1420 1213 1429 1216
rect 1442 1213 1484 1216
rect 1490 1213 1508 1216
rect 1522 1213 1556 1216
rect 1604 1213 1621 1216
rect 1660 1213 1685 1216
rect 1842 1213 1852 1216
rect 2002 1213 2020 1216
rect 2212 1213 2221 1216
rect 2434 1213 2444 1216
rect 730 1203 740 1206
rect 876 1203 909 1206
rect 930 1203 988 1206
rect 1098 1203 1108 1206
rect 1132 1203 1173 1206
rect 1234 1203 1292 1206
rect 1330 1203 1396 1206
rect 1428 1203 1461 1206
rect 1516 1203 1549 1206
rect 1674 1203 1684 1206
rect 1716 1203 1748 1206
rect 2058 1203 2068 1206
rect 2100 1203 2117 1206
rect 2218 1205 2221 1213
rect 2474 1206 2477 1226
rect 2482 1213 2492 1216
rect 2612 1213 2621 1216
rect 2676 1213 2701 1216
rect 2732 1213 2749 1216
rect 2756 1213 2781 1216
rect 2842 1213 2860 1216
rect 2426 1203 2436 1206
rect 2468 1203 2477 1206
rect 2500 1203 2517 1206
rect 2618 1205 2621 1213
rect 2746 1205 2749 1213
rect 2818 1203 2845 1206
rect 2890 1203 2893 1214
rect 3162 1213 3196 1216
rect 3340 1213 3349 1216
rect 3370 1213 3388 1216
rect 3508 1213 3533 1216
rect 3546 1213 3556 1216
rect 3586 1213 3612 1216
rect 3642 1213 3668 1216
rect 3698 1213 3708 1216
rect 3852 1213 3861 1216
rect 3908 1213 3933 1216
rect 3964 1213 3973 1216
rect 3994 1213 4012 1216
rect 4092 1213 4101 1216
rect 3346 1205 3349 1213
rect 3530 1205 3533 1213
rect 3620 1203 3637 1206
rect 3858 1205 3861 1213
rect 3970 1205 3973 1213
rect 890 1193 916 1196
rect 38 1167 4187 1173
rect 1818 1143 1844 1146
rect 2194 1143 2228 1146
rect 492 1133 517 1136
rect 540 1133 565 1136
rect 570 1133 580 1136
rect 1060 1133 1077 1136
rect 1226 1126 1229 1134
rect 1458 1126 1461 1134
rect 1548 1133 1557 1136
rect 1554 1126 1557 1133
rect 1754 1126 1757 1134
rect 1812 1133 1845 1136
rect 1852 1133 1861 1136
rect 2084 1133 2109 1136
rect 2130 1133 2156 1136
rect 2188 1133 2197 1136
rect 2236 1133 2245 1136
rect 2298 1133 2316 1136
rect 2674 1133 2708 1136
rect 2818 1133 2828 1136
rect 2844 1133 2853 1136
rect 108 1123 117 1126
rect 204 1123 213 1126
rect 300 1123 325 1126
rect 362 1123 372 1126
rect 412 1123 437 1126
rect 474 1123 484 1126
rect 490 1123 516 1126
rect 618 1123 628 1126
rect 692 1123 709 1126
rect 802 1123 812 1126
rect 884 1123 901 1126
rect 994 1123 1004 1126
rect 1068 1123 1085 1126
rect 1226 1123 1252 1126
rect 1396 1123 1413 1126
rect 1452 1123 1461 1126
rect 1498 1123 1524 1126
rect 1554 1123 1564 1126
rect 1692 1123 1717 1126
rect 1748 1123 1757 1126
rect 1948 1123 1973 1126
rect 2004 1123 2029 1126
rect 2124 1123 2149 1126
rect 2244 1123 2261 1126
rect 2300 1123 2317 1126
rect 2362 1123 2388 1126
rect 2532 1123 2541 1126
rect 2578 1123 2604 1126
rect 2732 1123 2765 1126
rect 2866 1123 2869 1134
rect 3066 1133 3092 1136
rect 3114 1133 3140 1136
rect 2930 1123 2956 1126
rect 2988 1123 2997 1126
rect 3002 1123 3012 1126
rect 3026 1123 3044 1126
rect 3074 1123 3133 1126
rect 3170 1123 3173 1134
rect 3218 1123 3221 1134
rect 3260 1133 3293 1136
rect 3322 1133 3340 1136
rect 3268 1123 3285 1126
rect 3362 1125 3365 1136
rect 3474 1133 3492 1136
rect 3508 1133 3541 1136
rect 3874 1133 3892 1136
rect 3914 1133 3948 1136
rect 3370 1123 3380 1126
rect 3410 1123 3436 1126
rect 3580 1123 3589 1126
rect 3772 1123 3797 1126
rect 3828 1123 3837 1126
rect 3882 1123 3900 1126
rect 3978 1123 3981 1134
rect 1812 1113 1837 1116
rect 2738 1113 2772 1116
rect 2796 1113 2813 1116
rect 2924 1113 2949 1116
rect 3178 1113 3188 1116
rect 3522 1113 3541 1116
rect 2780 1103 2789 1106
rect 14 1067 4211 1073
rect 1130 1023 1180 1026
rect 1242 1016 1245 1036
rect 2268 1023 2277 1026
rect 108 1013 125 1016
rect 218 1003 221 1014
rect 362 1013 372 1016
rect 460 1013 485 1016
rect 530 1013 540 1016
rect 570 1006 573 1014
rect 578 1006 581 1014
rect 322 1003 332 1006
rect 348 1003 364 1006
rect 532 1003 541 1006
rect 570 1003 581 1006
rect 610 1003 613 1014
rect 650 1006 653 1016
rect 668 1013 693 1016
rect 708 1013 725 1016
rect 772 1013 789 1016
rect 802 1013 812 1016
rect 842 1013 860 1016
rect 898 1013 924 1016
rect 972 1013 997 1016
rect 1034 1013 1044 1016
rect 1202 1013 1229 1016
rect 1236 1013 1245 1016
rect 1252 1013 1277 1016
rect 1332 1013 1357 1016
rect 1508 1013 1517 1016
rect 1618 1013 1628 1016
rect 1634 1013 1660 1016
rect 644 1003 653 1006
rect 660 1003 669 1006
rect 690 1005 693 1013
rect 716 1003 733 1006
rect 764 1003 773 1006
rect 786 1003 804 1006
rect 818 1003 868 1006
rect 884 1003 901 1006
rect 906 1003 916 1006
rect 930 1003 964 1006
rect 978 1003 1012 1006
rect 1106 1003 1116 1006
rect 1204 1003 1221 1006
rect 1226 1005 1229 1013
rect 1746 1006 1749 1014
rect 1826 1013 1852 1016
rect 1922 1013 1964 1016
rect 2028 1013 2053 1016
rect 2148 1013 2165 1016
rect 2210 1013 2252 1016
rect 1266 1003 1308 1006
rect 1522 1003 1556 1006
rect 1636 1003 1653 1006
rect 1706 1003 1724 1006
rect 1746 1003 1757 1006
rect 1780 1003 1789 1006
rect 1924 1003 1949 1006
rect 1972 1003 1989 1006
rect 2100 1003 2109 1006
rect 2170 1003 2180 1006
rect 2196 1003 2244 1006
rect 2266 1005 2269 1016
rect 2282 1013 2292 1016
rect 2354 1013 2364 1016
rect 2546 1006 2549 1016
rect 2588 1013 2605 1016
rect 2650 1013 2684 1016
rect 2756 1013 2765 1016
rect 2802 1013 2820 1016
rect 2900 1013 2925 1016
rect 2956 1013 2965 1016
rect 2972 1013 2981 1016
rect 3074 1013 3100 1016
rect 3172 1013 3197 1016
rect 2316 1003 2349 1006
rect 2410 1003 2420 1006
rect 2436 1003 2469 1006
rect 2532 1003 2564 1006
rect 2596 1003 2613 1006
rect 2692 1003 2717 1006
rect 2962 1005 2965 1013
rect 3234 1006 3237 1016
rect 3242 1013 3260 1016
rect 3292 1013 3309 1016
rect 3410 1013 3428 1016
rect 3458 1013 3484 1016
rect 3522 1013 3540 1016
rect 3546 1013 3580 1016
rect 3716 1013 3725 1016
rect 3868 1013 3877 1016
rect 3924 1013 3949 1016
rect 3980 1013 3989 1016
rect 4132 1013 4141 1016
rect 2994 1003 3004 1006
rect 3234 1003 3268 1006
rect 3284 1003 3317 1006
rect 3404 1003 3421 1006
rect 3548 1003 3565 1006
rect 3604 1003 3613 1006
rect 3722 1005 3725 1013
rect 3874 1005 3877 1013
rect 3986 1005 3989 1013
rect 4138 1005 4141 1013
rect 786 996 789 1003
rect 778 993 789 996
rect 898 996 901 1003
rect 898 993 909 996
rect 1522 993 1541 996
rect 38 967 4187 973
rect 722 943 740 946
rect 762 943 796 946
rect 962 943 980 946
rect 108 923 133 926
rect 186 925 189 936
rect 218 925 221 936
rect 266 933 292 936
rect 308 933 340 936
rect 428 933 477 936
rect 530 933 540 936
rect 594 933 604 936
rect 748 933 797 936
rect 804 933 813 936
rect 884 933 901 936
rect 906 933 932 936
rect 1010 933 1020 936
rect 1044 933 1069 936
rect 1074 933 1084 936
rect 898 926 901 933
rect 1114 926 1117 935
rect 1180 933 1197 936
rect 1354 933 1372 936
rect 1404 933 1429 936
rect 1444 933 1453 936
rect 1674 933 1724 936
rect 1794 933 1820 936
rect 1836 933 1861 936
rect 1994 933 2004 936
rect 2074 933 2084 936
rect 2098 933 2116 936
rect 2474 926 2477 935
rect 2500 933 2509 936
rect 2532 933 2565 936
rect 2602 933 2636 936
rect 2772 933 2781 936
rect 2820 933 2829 936
rect 2844 933 2861 936
rect 3004 933 3013 936
rect 3194 926 3197 935
rect 3380 933 3397 936
rect 3484 933 3493 936
rect 3650 933 3661 936
rect 3706 933 3724 936
rect 3770 933 3788 936
rect 3826 933 3860 936
rect 3876 933 3917 936
rect 3932 933 3973 936
rect 3978 933 4004 936
rect 4092 933 4125 936
rect 3650 926 3653 933
rect 316 923 341 926
rect 386 923 420 926
rect 426 923 476 926
rect 508 923 525 926
rect 538 923 548 926
rect 612 923 621 926
rect 716 923 725 926
rect 756 923 797 926
rect 812 923 853 926
rect 898 923 933 926
rect 1092 923 1117 926
rect 1130 923 1172 926
rect 1234 923 1260 926
rect 1290 923 1316 926
rect 1410 923 1436 926
rect 1508 923 1517 926
rect 1612 923 1637 926
rect 1668 923 1709 926
rect 1788 923 1805 926
rect 1900 923 1917 926
rect 2098 923 2124 926
rect 2316 923 2325 926
rect 2412 923 2437 926
rect 2468 923 2477 926
rect 2514 923 2524 926
rect 2604 923 2637 926
rect 2682 923 2708 926
rect 2818 923 2836 926
rect 2850 923 2868 926
rect 2898 923 2924 926
rect 3018 923 3028 926
rect 3068 923 3085 926
rect 3188 923 3197 926
rect 3210 923 3228 926
rect 3274 923 3284 926
rect 3402 923 3412 926
rect 3442 923 3476 926
rect 1132 913 1149 916
rect 2500 913 2509 916
rect 3594 913 3604 916
rect 3618 906 3621 925
rect 3644 923 3653 926
rect 3692 923 3716 926
rect 3748 923 3757 926
rect 3762 923 3796 926
rect 3834 923 3852 926
rect 3890 923 3924 926
rect 3970 923 3973 933
rect 4002 923 4012 926
rect 4042 923 4084 926
rect 4122 923 4125 933
rect 3754 916 3757 923
rect 3754 913 3773 916
rect 3618 903 3629 906
rect 14 867 4211 873
rect 988 823 1013 826
rect 1730 816 1733 826
rect 2690 823 2700 826
rect 2756 823 2765 826
rect 108 813 133 816
rect 204 813 221 816
rect 226 813 244 816
rect 276 813 309 816
rect 380 813 389 816
rect 476 813 501 816
rect 554 813 564 816
rect 652 813 677 816
rect 714 813 732 816
rect 738 813 756 816
rect 802 813 836 816
rect 884 813 893 816
rect 932 813 949 816
rect 1036 813 1084 816
rect 1274 813 1292 816
rect 1298 813 1324 816
rect 1380 813 1397 816
rect 1444 813 1469 816
rect 1538 813 1548 816
rect 1628 813 1637 816
rect 1730 813 1748 816
rect 1812 813 1821 816
rect 1892 813 1909 816
rect 1932 813 1941 816
rect 2012 813 2037 816
rect 2068 813 2077 816
rect 2122 813 2132 816
rect 2162 813 2172 816
rect 2284 813 2293 816
rect 2370 813 2380 816
rect 2508 813 2517 816
rect 2604 813 2612 816
rect 2644 813 2661 816
rect 2668 813 2693 816
rect 268 803 308 806
rect 548 803 565 806
rect 588 803 605 806
rect 740 803 757 806
rect 780 803 828 806
rect 852 803 869 806
rect 876 803 917 806
rect 930 803 964 806
rect 988 803 997 806
rect 1010 803 1020 806
rect 1044 803 1077 806
rect 1234 803 1244 806
rect 1276 803 1285 806
rect 1300 803 1317 806
rect 1338 803 1356 806
rect 1388 803 1405 806
rect 1516 803 1549 806
rect 1572 803 1589 806
rect 1690 803 1700 806
rect 1722 803 1740 806
rect 1884 803 1917 806
rect 1930 803 1948 806
rect 2074 805 2077 813
rect 2180 803 2189 806
rect 2290 805 2293 813
rect 2410 803 2420 806
rect 2436 803 2469 806
rect 2570 803 2580 806
rect 2596 803 2605 806
rect 2642 803 2660 806
rect 2746 803 2749 814
rect 2874 803 2877 814
rect 2908 813 2917 816
rect 2964 813 2997 816
rect 3034 813 3060 816
rect 3090 813 3116 816
rect 3154 813 3164 816
rect 3202 813 3220 816
rect 3282 813 3308 816
rect 3378 813 3404 816
rect 3572 813 3597 816
rect 3628 813 3653 816
rect 3850 813 3868 816
rect 2900 803 2933 806
rect 2972 803 2989 806
rect 3836 803 3861 806
rect 4140 803 4149 806
rect 890 793 916 796
rect 1890 793 1916 796
rect 2466 793 2469 803
rect 38 767 4187 773
rect 1178 736 1181 746
rect 3866 736 3869 756
rect 396 733 413 736
rect 108 723 125 726
rect 204 723 229 726
rect 266 723 276 726
rect 324 723 349 726
rect 394 723 412 726
rect 444 723 468 726
rect 498 725 501 736
rect 546 733 556 736
rect 588 733 597 736
rect 756 733 789 736
rect 586 723 596 726
rect 628 723 637 726
rect 684 723 709 726
rect 770 723 788 726
rect 818 725 821 736
rect 826 733 836 736
rect 860 733 877 736
rect 900 733 924 736
rect 954 733 980 736
rect 1002 726 1005 735
rect 1042 733 1052 736
rect 1090 733 1108 736
rect 1172 733 1181 736
rect 1220 733 1229 736
rect 1540 733 1557 736
rect 1586 733 1612 736
rect 1636 733 1645 736
rect 1674 733 1692 736
rect 1820 733 1829 736
rect 1852 733 1869 736
rect 1922 733 1940 736
rect 1964 733 1989 736
rect 2028 733 2045 736
rect 1042 726 1045 733
rect 1002 723 1013 726
rect 1034 723 1045 726
rect 1082 723 1116 726
rect 1164 723 1181 726
rect 1370 723 1388 726
rect 1460 723 1485 726
rect 1522 723 1532 726
rect 1546 723 1556 726
rect 1588 723 1620 726
rect 1628 723 1637 726
rect 1700 723 1709 726
rect 1746 723 1772 726
rect 1812 723 1821 726
rect 1860 723 1884 726
rect 1922 716 1925 733
rect 2466 726 2469 735
rect 2492 733 2501 736
rect 2508 733 2517 736
rect 1956 723 1989 726
rect 2034 723 2076 726
rect 2306 723 2324 726
rect 2460 723 2469 726
rect 2498 725 2501 733
rect 2586 723 2596 726
rect 2634 723 2652 726
rect 2722 723 2748 726
rect 2786 725 2789 736
rect 2818 725 2821 736
rect 2946 726 2949 735
rect 2868 723 2893 726
rect 2924 723 2949 726
rect 2994 725 2997 736
rect 3050 726 3053 735
rect 3316 733 3333 736
rect 3378 733 3396 736
rect 3634 726 3637 735
rect 3692 733 3701 736
rect 3866 733 3876 736
rect 3908 733 3933 736
rect 3050 723 3060 726
rect 3090 723 3116 726
rect 3188 723 3197 726
rect 3250 723 3292 726
rect 3426 723 3444 726
rect 3474 723 3500 726
rect 3572 723 3597 726
rect 3628 723 3637 726
rect 3644 723 3661 726
rect 3698 723 3724 726
rect 3852 723 3869 726
rect 3874 723 3884 726
rect 860 713 869 716
rect 948 713 973 716
rect 1042 713 1052 716
rect 1916 713 1925 716
rect 1986 713 1989 723
rect 2058 713 2061 723
rect 3372 713 3389 716
rect 14 667 4211 673
rect 866 626 869 636
rect 860 623 869 626
rect 1042 623 1052 626
rect 1892 623 1909 626
rect 1938 623 1972 626
rect 138 613 156 616
rect 228 613 253 616
rect 298 613 316 616
rect 348 613 372 616
rect 420 613 445 616
rect 482 613 492 616
rect 612 613 621 616
rect 658 613 684 616
rect 730 613 740 616
rect 828 613 837 616
rect 858 613 877 616
rect 946 613 972 616
rect 1194 613 1220 616
rect 1276 613 1301 616
rect 1332 613 1341 616
rect 1444 613 1469 616
rect 1556 613 1565 616
rect 1698 613 1716 616
rect 1788 613 1805 616
rect 1844 613 1869 616
rect 874 606 877 613
rect 132 603 149 606
rect 180 603 189 606
rect 300 603 317 606
rect 354 603 364 606
rect 498 603 508 606
rect 546 603 564 606
rect 770 603 780 606
rect 826 603 836 606
rect 860 603 869 606
rect 874 603 884 606
rect 1010 603 1052 606
rect 1076 603 1085 606
rect 1186 603 1212 606
rect 1338 605 1341 613
rect 1516 603 1525 606
rect 1548 603 1564 606
rect 1866 605 1869 613
rect 1994 613 2020 616
rect 2082 613 2092 616
rect 2122 613 2148 616
rect 2186 613 2220 616
rect 2260 613 2293 616
rect 2314 613 2340 616
rect 1892 603 1917 606
rect 1924 603 1933 606
rect 1938 603 1972 606
rect 1994 605 1997 613
rect 2002 603 2012 606
rect 2042 603 2052 606
rect 2266 603 2292 606
rect 2322 603 2332 606
rect 2356 603 2373 606
rect 2394 603 2397 614
rect 2428 613 2445 616
rect 2578 606 2581 614
rect 2586 606 2589 614
rect 2620 613 2629 616
rect 2660 613 2668 616
rect 2748 613 2773 616
rect 2804 613 2813 616
rect 2852 613 2869 616
rect 2900 613 2917 616
rect 3012 613 3021 616
rect 3042 613 3052 616
rect 3058 613 3068 616
rect 3098 613 3124 616
rect 3196 613 3213 616
rect 3252 613 3261 616
rect 3274 613 3284 616
rect 3330 613 3340 616
rect 3378 613 3388 616
rect 3564 613 3589 616
rect 3620 613 3629 616
rect 3636 613 3661 616
rect 3706 613 3724 616
rect 3938 613 3964 616
rect 4132 613 4141 616
rect 2420 603 2452 606
rect 2476 603 2501 606
rect 2540 603 2556 606
rect 2578 603 2589 606
rect 2618 603 2628 606
rect 2810 605 2813 613
rect 2866 603 2892 606
rect 2906 603 2924 606
rect 3020 603 3037 606
rect 3058 605 3061 613
rect 3258 605 3261 613
rect 3308 603 3333 606
rect 3348 603 3373 606
rect 3418 603 3444 606
rect 3626 605 3629 613
rect 3714 603 3732 606
rect 4138 605 4141 613
rect 1930 596 1933 603
rect 794 593 812 596
rect 1898 593 1916 596
rect 1930 593 1965 596
rect 38 567 4187 573
rect 954 543 980 546
rect 1906 543 1916 546
rect 108 523 133 526
rect 170 525 173 536
rect 196 533 212 536
rect 226 533 244 536
rect 276 533 316 536
rect 332 533 341 536
rect 460 533 477 536
rect 514 533 532 536
rect 564 533 581 536
rect 586 533 604 536
rect 626 533 644 536
rect 586 526 589 533
rect 268 523 277 526
rect 388 523 413 526
rect 458 523 476 526
rect 562 523 589 526
rect 690 523 716 526
rect 858 525 861 536
rect 884 533 893 536
rect 898 533 908 536
rect 970 533 988 536
rect 1330 526 1333 535
rect 1508 533 1533 536
rect 1604 533 1621 536
rect 1666 533 1692 536
rect 1716 533 1725 536
rect 1852 533 1876 536
rect 1900 533 1917 536
rect 1924 533 1933 536
rect 2162 526 2165 535
rect 2298 526 2301 535
rect 2476 533 2485 536
rect 2508 533 2525 536
rect 2532 533 2581 536
rect 2636 533 2645 536
rect 2684 533 2693 536
rect 2756 533 2773 536
rect 3130 533 3156 536
rect 3172 533 3197 536
rect 2770 526 2773 533
rect 3306 526 3309 535
rect 3466 526 3469 535
rect 916 523 925 526
rect 996 523 1005 526
rect 1268 523 1293 526
rect 1324 523 1333 526
rect 1436 523 1461 526
rect 1506 523 1532 526
rect 1610 523 1636 526
rect 1668 523 1677 526
rect 1708 523 1725 526
rect 1860 523 1869 526
rect 1874 523 1884 526
rect 2010 523 2028 526
rect 2100 523 2125 526
rect 2156 523 2165 526
rect 2292 523 2301 526
rect 2314 523 2324 526
rect 2482 523 2492 526
rect 2596 523 2605 526
rect 2714 523 2740 526
rect 2770 523 2796 526
rect 3130 523 3148 526
rect 3180 523 3205 526
rect 3244 523 3269 526
rect 3300 523 3309 526
rect 3356 523 3365 526
rect 3460 523 3469 526
rect 3666 525 3669 536
rect 3810 526 3813 535
rect 3804 523 3813 526
rect 3826 523 3836 526
rect 3850 525 3853 536
rect 3876 533 3893 536
rect 4050 526 4053 535
rect 4092 533 4149 536
rect 4044 523 4053 526
rect 4066 523 4084 526
rect 4146 523 4149 533
rect 948 513 973 516
rect 1900 513 1909 516
rect 3052 513 3077 516
rect 3578 513 3596 516
rect 3620 513 3629 516
rect 14 467 4211 473
rect 1900 423 1909 426
rect 2380 423 2389 426
rect 2802 423 2828 426
rect 3212 423 3229 426
rect 260 413 285 416
rect 322 413 332 416
rect 388 413 413 416
rect 186 403 196 406
rect 460 403 469 406
rect 498 403 501 414
rect 588 413 597 416
rect 642 413 668 416
rect 722 406 725 414
rect 748 413 757 416
rect 812 413 821 416
rect 922 413 932 416
rect 970 413 980 416
rect 1156 413 1181 416
rect 1212 413 1221 416
rect 1268 413 1293 416
rect 1324 413 1333 416
rect 1372 413 1396 416
rect 1476 413 1501 416
rect 516 403 533 406
rect 722 403 732 406
rect 772 403 781 406
rect 860 403 869 406
rect 1218 405 1221 413
rect 1330 405 1333 413
rect 1548 403 1557 406
rect 1618 403 1628 406
rect 1650 403 1653 414
rect 1690 413 1716 416
rect 1788 413 1805 416
rect 1852 413 1861 416
rect 1874 413 1884 416
rect 2020 413 2037 416
rect 2076 413 2085 416
rect 2236 413 2261 416
rect 2292 413 2309 416
rect 2316 413 2357 416
rect 2466 413 2492 416
rect 2602 413 2628 416
rect 2716 413 2725 416
rect 2756 413 2780 416
rect 2892 413 2917 416
rect 2948 413 2965 416
rect 2996 413 3005 416
rect 3066 413 3076 416
rect 3082 413 3092 416
rect 3122 413 3148 416
rect 3362 413 3380 416
rect 3508 413 3525 416
rect 3788 413 3805 416
rect 3850 413 3876 416
rect 3906 413 3932 416
rect 3994 413 4004 416
rect 4140 413 4149 416
rect 1860 403 1869 406
rect 1900 403 1917 406
rect 1924 403 1933 406
rect 1938 403 1948 406
rect 1972 403 1981 406
rect 2082 405 2085 413
rect 2098 403 2108 406
rect 2306 405 2309 413
rect 2354 405 2357 413
rect 3066 406 3069 413
rect 2380 403 2389 406
rect 2556 403 2565 406
rect 2714 403 2724 406
rect 2954 403 2972 406
rect 3010 403 3036 406
rect 3052 403 3069 406
rect 3082 405 3085 413
rect 3260 403 3269 406
rect 3284 403 3309 406
rect 3354 403 3372 406
rect 3522 405 3525 413
rect 3802 405 3805 413
rect 3970 403 3996 406
rect 1906 393 1916 396
rect 38 367 4187 373
rect 148 333 181 336
rect 204 333 213 336
rect 218 333 228 336
rect 106 323 124 326
rect 130 323 140 326
rect 170 323 180 326
rect 252 323 276 326
rect 418 325 421 336
rect 444 333 453 336
rect 554 333 564 336
rect 492 323 509 326
rect 594 325 597 336
rect 1028 333 1037 336
rect 1074 333 1084 336
rect 1108 333 1117 336
rect 1122 326 1125 335
rect 1154 326 1157 335
rect 1314 326 1317 335
rect 1066 323 1092 326
rect 1106 323 1125 326
rect 1146 323 1157 326
rect 1252 323 1277 326
rect 1308 323 1317 326
rect 1402 326 1405 335
rect 1532 333 1549 336
rect 1578 333 1588 336
rect 1620 333 1637 336
rect 1858 333 1868 336
rect 1924 333 1933 336
rect 1940 333 1949 336
rect 1634 326 1637 333
rect 1986 326 1989 335
rect 2290 326 2293 335
rect 1402 323 1413 326
rect 1460 323 1485 326
rect 1530 323 1548 326
rect 1586 323 1596 326
rect 1634 323 1652 326
rect 1746 323 1756 326
rect 1796 323 1821 326
rect 1978 323 1989 326
rect 2058 323 2068 326
rect 2130 323 2156 326
rect 2228 323 2253 326
rect 2284 323 2293 326
rect 2300 323 2309 326
rect 2346 323 2349 335
rect 2410 326 2413 335
rect 2418 333 2428 336
rect 2370 323 2389 326
rect 2410 323 2429 326
rect 2508 323 2533 326
rect 2570 323 2580 326
rect 2586 325 2589 336
rect 2602 333 2612 336
rect 2684 333 2693 336
rect 2946 326 2949 335
rect 3042 333 3060 336
rect 3076 333 3093 336
rect 2682 323 2692 326
rect 2786 323 2812 326
rect 2884 323 2909 326
rect 2940 323 2949 326
rect 3090 326 3093 333
rect 3106 326 3109 335
rect 3604 333 3613 336
rect 3090 323 3100 326
rect 3106 323 3124 326
rect 3154 323 3180 326
rect 3252 323 3277 326
rect 3498 323 3508 326
rect 3554 323 3564 326
rect 3596 323 3605 326
rect 1068 313 1077 316
rect 1108 313 1117 316
rect 2370 315 2373 323
rect 3618 316 3621 336
rect 3802 326 3805 335
rect 3876 333 3901 336
rect 4042 326 4045 335
rect 3796 323 3805 326
rect 3842 323 3852 326
rect 4036 323 4045 326
rect 2378 313 2388 316
rect 3482 313 3492 316
rect 3514 313 3524 316
rect 3618 313 3628 316
rect 14 267 4211 273
rect 1050 216 1053 226
rect 2034 216 2037 225
rect 108 213 133 216
rect 244 213 252 216
rect 314 213 340 216
rect 372 213 381 216
rect 442 213 452 216
rect 484 213 493 216
rect 506 213 516 216
rect 634 213 652 216
rect 756 213 765 216
rect 802 213 812 216
rect 850 213 860 216
rect 914 213 924 216
rect 1044 213 1053 216
rect 1084 213 1093 216
rect 1188 213 1197 216
rect 1332 213 1357 216
rect 1388 213 1397 216
rect 1410 213 1436 216
rect 1450 213 1460 216
rect 1492 213 1533 216
rect 1546 213 1556 216
rect 1594 213 1612 216
rect 180 203 213 206
rect 370 203 404 206
rect 482 203 492 206
rect 540 203 549 206
rect 620 203 644 206
rect 748 203 764 206
rect 804 203 813 206
rect 836 203 852 206
rect 876 203 885 206
rect 916 203 925 206
rect 948 203 957 206
rect 1036 203 1045 206
rect 1050 203 1068 206
rect 1394 205 1397 213
rect 1674 206 1677 214
rect 1738 213 1748 216
rect 1826 213 1836 216
rect 1410 203 1428 206
rect 1452 203 1461 206
rect 1484 203 1501 206
rect 1548 203 1557 206
rect 1586 203 1604 206
rect 1636 203 1652 206
rect 1674 203 1685 206
rect 1714 203 1740 206
rect 1772 203 1788 206
rect 1828 203 1837 206
rect 1874 203 1877 214
rect 1954 213 1964 216
rect 2034 213 2045 216
rect 2114 213 2124 216
rect 2154 213 2164 216
rect 2284 213 2293 216
rect 2306 213 2316 216
rect 2346 213 2365 216
rect 2444 213 2452 216
rect 2484 213 2493 216
rect 2548 213 2565 216
rect 2604 213 2612 216
rect 2644 213 2661 216
rect 2676 213 2685 216
rect 2690 213 2700 216
rect 2794 213 2820 216
rect 2908 213 2925 216
rect 2970 213 2988 216
rect 3018 213 3044 216
rect 3074 213 3084 216
rect 3114 213 3140 216
rect 3178 213 3196 216
rect 3274 213 3284 216
rect 3322 213 3348 216
rect 3378 213 3396 216
rect 3428 213 3453 216
rect 3458 213 3468 216
rect 3500 213 3525 216
rect 3610 213 3620 216
rect 3652 213 3661 216
rect 3738 213 3748 216
rect 3796 213 3804 216
rect 3890 213 3908 216
rect 3970 213 3980 216
rect 3994 213 4020 216
rect 4050 213 4076 216
rect 4082 213 4092 216
rect 1900 203 1917 206
rect 1946 203 1956 206
rect 1980 203 1989 206
rect 1996 203 2005 206
rect 2042 205 2045 213
rect 2068 203 2077 206
rect 2290 205 2293 213
rect 2362 205 2365 213
rect 2922 206 2925 213
rect 3450 206 3453 213
rect 4146 206 4149 216
rect 2404 203 2413 206
rect 2442 203 2460 206
rect 2482 203 2492 206
rect 2554 203 2580 206
rect 2596 203 2613 206
rect 2642 203 2668 206
rect 2698 203 2708 206
rect 2738 203 2748 206
rect 2922 203 2940 206
rect 2956 203 2973 206
rect 3018 203 3036 206
rect 3226 203 3236 206
rect 3252 203 3269 206
rect 3308 203 3324 206
rect 3378 203 3388 206
rect 3436 203 3445 206
rect 3450 203 3476 206
rect 3498 203 3524 206
rect 3562 203 3572 206
rect 3588 203 3605 206
rect 3660 203 3669 206
rect 3692 203 3701 206
rect 3756 203 3765 206
rect 3932 203 3940 206
rect 3988 203 4005 206
rect 4100 203 4149 206
rect 38 167 4187 173
rect 1386 126 1389 135
rect 1890 133 1908 136
rect 2018 133 2028 136
rect 2234 126 2237 135
rect 2730 133 2740 136
rect 3050 126 3053 135
rect 3194 126 3197 135
rect 3306 126 3309 135
rect 3418 126 3421 135
rect 3546 126 3549 135
rect 204 123 229 126
rect 266 123 276 126
rect 386 123 412 126
rect 498 123 516 126
rect 900 123 909 126
rect 1212 123 1221 126
rect 1372 123 1389 126
rect 1674 123 1700 126
rect 1834 123 1844 126
rect 1954 123 1980 126
rect 2074 123 2100 126
rect 2228 123 2237 126
rect 2284 123 2309 126
rect 2380 123 2397 126
rect 2682 123 2692 126
rect 2786 123 2812 126
rect 2988 123 2997 126
rect 3044 123 3053 126
rect 3124 123 3149 126
rect 3180 123 3197 126
rect 3244 123 3269 126
rect 3300 123 3309 126
rect 3412 123 3421 126
rect 3484 123 3509 126
rect 3540 123 3549 126
rect 3620 123 3629 126
rect 3836 123 3861 126
rect 14 67 4211 73
rect 38 37 4187 57
rect 14 13 4211 33
<< metal2 >>
rect 14 13 34 4127
rect 38 37 58 4103
rect 1842 4056 1845 4140
rect 1834 4053 1845 4056
rect 154 4023 173 4026
rect 82 3593 85 4006
rect 130 4003 133 4016
rect 154 3936 157 4023
rect 162 3983 165 4016
rect 170 4013 173 4023
rect 150 3933 157 3936
rect 114 3813 117 3926
rect 150 3886 153 3933
rect 146 3883 153 3886
rect 122 3793 125 3816
rect 130 3796 133 3836
rect 138 3803 141 3826
rect 146 3813 149 3883
rect 162 3833 165 3926
rect 170 3923 173 4006
rect 178 3983 181 4006
rect 186 3976 189 4016
rect 178 3973 189 3976
rect 178 3933 181 3973
rect 194 3933 197 3946
rect 162 3813 165 3826
rect 146 3796 149 3806
rect 130 3793 149 3796
rect 106 3746 109 3766
rect 106 3743 117 3746
rect 114 3696 117 3743
rect 130 3713 133 3726
rect 106 3693 117 3696
rect 106 3646 109 3693
rect 106 3643 117 3646
rect 114 3596 117 3643
rect 130 3603 133 3616
rect 106 3593 117 3596
rect 82 3143 85 3556
rect 106 3476 109 3593
rect 98 3473 109 3476
rect 98 3406 101 3473
rect 114 3413 117 3526
rect 146 3513 149 3596
rect 98 3403 109 3406
rect 106 3346 109 3403
rect 106 3343 113 3346
rect 110 3296 113 3343
rect 106 3293 113 3296
rect 106 3246 109 3293
rect 106 3243 113 3246
rect 110 3196 113 3243
rect 106 3193 113 3196
rect 82 3123 85 3136
rect 82 2606 85 3116
rect 106 2966 109 3193
rect 98 2963 109 2966
rect 98 2866 101 2963
rect 114 2946 117 3126
rect 110 2943 117 2946
rect 110 2886 113 2943
rect 110 2883 117 2886
rect 98 2863 109 2866
rect 106 2633 109 2863
rect 114 2623 117 2883
rect 90 2613 117 2616
rect 74 2586 77 2606
rect 82 2603 101 2606
rect 74 2583 85 2586
rect 66 1786 69 2566
rect 66 1783 77 1786
rect 74 1706 77 1783
rect 82 1776 85 2583
rect 106 2523 109 2606
rect 114 2593 117 2613
rect 98 2396 101 2426
rect 106 2406 109 2436
rect 114 2413 117 2526
rect 122 2463 125 3386
rect 138 3363 141 3456
rect 146 3403 149 3426
rect 130 3313 133 3326
rect 130 3213 133 3226
rect 130 3113 133 3126
rect 130 2923 133 3016
rect 146 2943 149 3356
rect 154 3106 157 3746
rect 162 3723 165 3756
rect 170 3723 173 3796
rect 178 3763 181 3816
rect 178 3733 181 3756
rect 194 3733 197 3816
rect 202 3813 205 3826
rect 218 3813 221 4006
rect 234 3936 237 4016
rect 250 4013 253 4026
rect 290 4013 293 4026
rect 242 3993 245 4006
rect 266 3956 269 4006
rect 262 3953 269 3956
rect 234 3933 241 3936
rect 226 3813 229 3926
rect 238 3806 241 3933
rect 262 3906 265 3953
rect 290 3933 293 3946
rect 274 3913 277 3926
rect 262 3903 269 3906
rect 234 3803 241 3806
rect 218 3733 221 3766
rect 234 3743 237 3803
rect 162 3543 165 3616
rect 170 3613 173 3716
rect 186 3656 189 3726
rect 178 3653 189 3656
rect 162 3403 165 3526
rect 170 3523 173 3606
rect 178 3603 181 3653
rect 170 3413 173 3426
rect 162 3303 165 3396
rect 178 3383 181 3566
rect 194 3553 197 3716
rect 202 3703 205 3726
rect 218 3646 221 3726
rect 242 3713 245 3766
rect 250 3696 253 3816
rect 266 3763 269 3903
rect 282 3813 285 3926
rect 298 3923 301 3996
rect 282 3796 285 3806
rect 290 3803 293 3816
rect 298 3796 301 3816
rect 306 3803 309 3916
rect 322 3903 325 3926
rect 322 3813 325 3846
rect 282 3793 301 3796
rect 314 3793 317 3806
rect 258 3713 261 3726
rect 290 3723 301 3726
rect 306 3713 309 3726
rect 314 3703 317 3726
rect 322 3713 325 3736
rect 234 3693 253 3696
rect 218 3643 225 3646
rect 222 3596 225 3643
rect 218 3593 225 3596
rect 186 3543 205 3546
rect 186 3533 189 3543
rect 194 3523 197 3536
rect 202 3523 205 3543
rect 210 3533 213 3546
rect 186 3413 189 3426
rect 186 3373 189 3406
rect 170 3313 173 3326
rect 162 3213 165 3236
rect 178 3226 181 3366
rect 202 3353 205 3516
rect 218 3513 221 3593
rect 226 3423 229 3526
rect 234 3506 237 3693
rect 242 3613 245 3626
rect 242 3543 261 3546
rect 242 3523 245 3543
rect 250 3523 253 3536
rect 258 3533 261 3543
rect 234 3503 241 3506
rect 186 3343 205 3346
rect 186 3333 189 3343
rect 194 3303 197 3336
rect 202 3323 205 3343
rect 170 3213 173 3226
rect 178 3223 189 3226
rect 162 3123 165 3196
rect 178 3126 181 3223
rect 186 3183 189 3206
rect 194 3193 197 3206
rect 202 3176 205 3216
rect 186 3173 205 3176
rect 186 3133 189 3173
rect 194 3133 197 3146
rect 170 3113 173 3126
rect 178 3123 189 3126
rect 186 3106 189 3123
rect 154 3103 161 3106
rect 158 3036 161 3103
rect 154 3033 161 3036
rect 182 3103 189 3106
rect 182 3036 185 3103
rect 182 3033 189 3036
rect 138 2923 141 2936
rect 146 2913 149 2936
rect 130 2813 133 2826
rect 130 2616 133 2726
rect 154 2683 157 3033
rect 162 2933 165 3016
rect 170 2933 173 3016
rect 186 3013 189 3033
rect 170 2913 173 2926
rect 186 2916 189 3006
rect 194 3003 197 3116
rect 202 3056 205 3126
rect 210 3113 213 3376
rect 218 3333 221 3366
rect 226 3323 229 3416
rect 238 3406 241 3503
rect 258 3483 261 3526
rect 266 3456 269 3616
rect 274 3593 277 3616
rect 282 3613 285 3626
rect 290 3563 293 3616
rect 306 3596 309 3606
rect 314 3603 317 3616
rect 322 3596 325 3616
rect 330 3613 333 3946
rect 338 3923 341 4006
rect 346 3933 349 4016
rect 394 4013 397 4026
rect 434 4013 437 4026
rect 354 3933 357 3946
rect 354 3923 365 3926
rect 370 3923 373 4006
rect 410 3973 413 4006
rect 386 3933 389 3956
rect 362 3816 365 3906
rect 386 3903 389 3926
rect 394 3913 397 3936
rect 410 3933 421 3936
rect 426 3933 429 3966
rect 434 3933 437 3986
rect 402 3903 405 3926
rect 418 3916 421 3926
rect 418 3913 429 3916
rect 346 3796 349 3816
rect 354 3803 357 3816
rect 362 3813 373 3816
rect 378 3813 381 3826
rect 418 3813 421 3826
rect 362 3796 365 3806
rect 346 3793 365 3796
rect 370 3746 373 3813
rect 394 3786 397 3806
rect 426 3796 429 3913
rect 338 3713 341 3726
rect 346 3723 349 3746
rect 354 3743 373 3746
rect 386 3783 397 3786
rect 422 3793 429 3796
rect 354 3696 357 3743
rect 346 3693 357 3696
rect 346 3636 349 3693
rect 346 3633 357 3636
rect 354 3613 357 3633
rect 362 3616 365 3736
rect 386 3733 389 3783
rect 370 3713 373 3726
rect 410 3713 413 3726
rect 362 3613 389 3616
rect 306 3593 325 3596
rect 330 3593 333 3606
rect 338 3566 341 3606
rect 378 3593 381 3606
rect 394 3603 397 3616
rect 402 3593 405 3606
rect 330 3563 341 3566
rect 274 3513 277 3526
rect 290 3496 293 3536
rect 314 3513 317 3526
rect 234 3403 241 3406
rect 250 3453 269 3456
rect 286 3493 293 3496
rect 234 3323 237 3403
rect 250 3373 253 3453
rect 286 3436 289 3493
rect 330 3486 333 3563
rect 362 3523 373 3526
rect 378 3496 381 3576
rect 410 3573 413 3666
rect 422 3566 425 3793
rect 386 3523 389 3536
rect 394 3533 397 3566
rect 422 3563 429 3566
rect 402 3523 405 3556
rect 410 3503 413 3536
rect 418 3533 421 3546
rect 426 3523 429 3563
rect 434 3513 437 3926
rect 450 3883 453 3936
rect 466 3933 469 3956
rect 490 3953 493 4016
rect 514 4013 517 4026
rect 554 4013 557 4026
rect 506 3966 509 4006
rect 506 3963 517 3966
rect 498 3933 501 3946
rect 458 3913 461 3926
rect 466 3923 477 3926
rect 506 3923 509 3936
rect 514 3923 517 3963
rect 458 3813 477 3816
rect 474 3803 477 3813
rect 482 3803 485 3836
rect 490 3813 493 3826
rect 506 3813 509 3916
rect 498 3783 501 3806
rect 506 3803 517 3806
rect 530 3793 533 4006
rect 554 3933 557 3956
rect 610 3953 613 4016
rect 634 3993 637 4006
rect 594 3943 613 3946
rect 594 3933 597 3943
rect 554 3893 557 3926
rect 562 3813 565 3926
rect 474 3733 477 3756
rect 474 3706 477 3726
rect 466 3703 477 3706
rect 466 3636 469 3703
rect 466 3633 477 3636
rect 442 3553 445 3626
rect 450 3573 453 3606
rect 450 3533 453 3546
rect 458 3533 461 3616
rect 474 3593 477 3633
rect 482 3613 485 3726
rect 490 3723 493 3736
rect 506 3733 509 3746
rect 498 3623 501 3726
rect 514 3713 517 3736
rect 522 3613 525 3726
rect 530 3663 533 3736
rect 538 3733 541 3746
rect 546 3713 549 3726
rect 570 3696 573 3896
rect 578 3843 581 3926
rect 602 3876 605 3936
rect 610 3923 613 3943
rect 594 3873 605 3876
rect 566 3693 573 3696
rect 466 3533 469 3586
rect 450 3523 461 3526
rect 362 3493 381 3496
rect 242 3343 261 3346
rect 242 3333 245 3343
rect 242 3316 245 3326
rect 250 3323 253 3336
rect 258 3323 261 3343
rect 266 3326 269 3436
rect 286 3433 293 3436
rect 282 3376 285 3416
rect 290 3413 293 3433
rect 298 3413 301 3486
rect 330 3483 341 3486
rect 338 3453 341 3483
rect 330 3416 333 3436
rect 314 3406 317 3416
rect 322 3413 333 3416
rect 290 3383 293 3406
rect 274 3373 285 3376
rect 274 3333 277 3373
rect 266 3323 277 3326
rect 242 3313 261 3316
rect 218 3213 221 3246
rect 226 3213 229 3226
rect 234 3203 237 3236
rect 242 3183 245 3216
rect 250 3173 253 3206
rect 258 3203 261 3313
rect 282 3263 285 3336
rect 298 3333 301 3406
rect 306 3383 309 3406
rect 314 3403 325 3406
rect 218 3093 221 3126
rect 234 3123 237 3136
rect 202 3053 221 3056
rect 218 3003 221 3053
rect 226 3013 229 3106
rect 258 3103 261 3126
rect 234 3003 237 3026
rect 202 2923 205 2966
rect 218 2933 221 2946
rect 186 2913 197 2916
rect 194 2896 197 2913
rect 194 2893 205 2896
rect 162 2793 165 2816
rect 170 2813 173 2826
rect 186 2813 189 2866
rect 202 2836 205 2893
rect 194 2833 205 2836
rect 170 2803 181 2806
rect 162 2723 165 2736
rect 194 2733 197 2833
rect 202 2803 205 2816
rect 218 2813 221 2926
rect 242 2923 245 3016
rect 250 2963 253 3036
rect 266 3013 269 3026
rect 258 2983 261 3006
rect 274 2993 277 3216
rect 298 3213 301 3326
rect 306 3313 309 3326
rect 322 3213 325 3403
rect 330 3363 333 3413
rect 338 3403 341 3416
rect 354 3413 357 3446
rect 362 3413 365 3493
rect 458 3456 461 3523
rect 482 3486 485 3606
rect 498 3593 501 3606
rect 498 3496 501 3556
rect 506 3503 509 3536
rect 514 3523 517 3536
rect 498 3493 509 3496
rect 482 3483 493 3486
rect 450 3453 461 3456
rect 362 3363 365 3406
rect 370 3346 373 3406
rect 378 3373 381 3416
rect 386 3403 389 3426
rect 394 3386 397 3446
rect 410 3403 413 3416
rect 390 3383 397 3386
rect 362 3343 373 3346
rect 346 3313 349 3326
rect 362 3266 365 3343
rect 390 3326 393 3383
rect 390 3323 397 3326
rect 402 3323 405 3366
rect 410 3333 413 3376
rect 434 3346 437 3416
rect 450 3376 453 3453
rect 490 3413 493 3483
rect 506 3413 509 3493
rect 530 3446 533 3646
rect 566 3606 569 3693
rect 578 3613 581 3736
rect 586 3733 589 3746
rect 586 3703 589 3726
rect 566 3603 573 3606
rect 554 3523 557 3536
rect 530 3443 541 3446
rect 498 3393 501 3406
rect 450 3373 461 3376
rect 514 3373 517 3406
rect 522 3393 525 3416
rect 530 3413 533 3436
rect 426 3343 437 3346
rect 426 3323 429 3343
rect 442 3336 445 3346
rect 434 3333 445 3336
rect 394 3306 397 3323
rect 394 3303 405 3306
rect 362 3263 373 3266
rect 354 3213 357 3226
rect 362 3213 365 3246
rect 298 3166 301 3206
rect 298 3163 305 3166
rect 302 3086 305 3163
rect 314 3123 317 3146
rect 362 3136 365 3206
rect 370 3203 373 3263
rect 378 3213 381 3266
rect 402 3236 405 3303
rect 394 3233 405 3236
rect 386 3203 389 3226
rect 322 3113 325 3136
rect 346 3133 365 3136
rect 298 3083 305 3086
rect 298 3026 301 3083
rect 330 3066 333 3126
rect 338 3093 341 3126
rect 330 3063 341 3066
rect 282 3023 301 3026
rect 282 2986 285 3023
rect 290 3003 293 3016
rect 338 3013 341 3063
rect 282 2983 289 2986
rect 210 2793 213 2806
rect 202 2733 213 2736
rect 218 2733 221 2806
rect 234 2783 237 2806
rect 258 2796 261 2946
rect 286 2886 289 2983
rect 298 2923 301 3006
rect 314 2993 317 3006
rect 306 2896 309 2986
rect 346 2983 349 3133
rect 354 3113 357 3126
rect 370 3056 373 3126
rect 378 3106 381 3146
rect 386 3133 389 3156
rect 394 3126 397 3233
rect 386 3123 397 3126
rect 402 3113 405 3126
rect 378 3103 389 3106
rect 354 3053 373 3056
rect 330 2943 349 2946
rect 282 2883 289 2886
rect 298 2893 309 2896
rect 282 2836 285 2883
rect 298 2856 301 2893
rect 314 2863 317 2926
rect 330 2923 333 2943
rect 338 2923 341 2936
rect 346 2933 349 2943
rect 298 2853 305 2856
rect 250 2793 261 2796
rect 274 2833 285 2836
rect 170 2656 173 2726
rect 178 2713 181 2726
rect 186 2693 189 2726
rect 170 2653 197 2656
rect 130 2613 149 2616
rect 154 2613 157 2626
rect 138 2603 149 2606
rect 170 2603 173 2616
rect 194 2613 197 2653
rect 202 2623 205 2726
rect 210 2663 213 2733
rect 226 2716 229 2776
rect 250 2756 253 2793
rect 222 2713 229 2716
rect 234 2753 253 2756
rect 222 2656 225 2713
rect 218 2653 225 2656
rect 138 2563 141 2603
rect 170 2533 173 2596
rect 202 2533 205 2616
rect 218 2576 221 2653
rect 234 2603 237 2753
rect 242 2706 245 2746
rect 258 2733 261 2786
rect 274 2773 277 2833
rect 282 2813 285 2826
rect 250 2713 253 2726
rect 242 2703 253 2706
rect 266 2703 269 2766
rect 274 2733 285 2736
rect 274 2713 277 2726
rect 242 2596 245 2686
rect 250 2613 253 2703
rect 282 2666 285 2726
rect 290 2713 293 2776
rect 302 2756 305 2853
rect 314 2813 317 2836
rect 322 2813 325 2826
rect 330 2813 333 2856
rect 298 2753 305 2756
rect 298 2723 301 2753
rect 306 2723 309 2736
rect 282 2663 293 2666
rect 290 2613 293 2663
rect 314 2623 317 2736
rect 322 2713 325 2806
rect 338 2796 341 2806
rect 346 2803 349 2836
rect 354 2823 357 3053
rect 386 3036 389 3103
rect 410 3063 413 3136
rect 418 3123 421 3216
rect 442 3213 445 3326
rect 450 3243 453 3336
rect 458 3213 461 3373
rect 466 3233 469 3336
rect 474 3323 477 3336
rect 482 3313 485 3326
rect 450 3183 453 3206
rect 466 3193 469 3206
rect 426 3133 429 3146
rect 378 3033 389 3036
rect 378 3016 381 3033
rect 378 3013 397 3016
rect 410 3003 413 3016
rect 362 2913 365 2926
rect 378 2886 381 2996
rect 402 2913 405 2926
rect 378 2883 389 2886
rect 354 2796 357 2816
rect 370 2813 373 2826
rect 338 2793 357 2796
rect 362 2783 365 2806
rect 370 2763 373 2806
rect 386 2756 389 2883
rect 330 2733 333 2756
rect 370 2753 389 2756
rect 346 2743 365 2746
rect 330 2703 333 2726
rect 338 2606 341 2736
rect 346 2723 349 2743
rect 354 2723 357 2736
rect 362 2733 365 2743
rect 362 2713 365 2726
rect 346 2613 349 2626
rect 354 2613 357 2696
rect 370 2633 373 2753
rect 378 2723 381 2736
rect 386 2733 389 2746
rect 402 2733 405 2766
rect 410 2733 413 2816
rect 418 2773 421 2966
rect 442 2883 445 3156
rect 482 3123 485 3216
rect 474 3056 477 3116
rect 490 3103 493 3256
rect 498 3166 501 3346
rect 522 3336 525 3386
rect 530 3363 533 3406
rect 538 3383 541 3443
rect 546 3366 549 3416
rect 554 3413 557 3506
rect 570 3483 573 3603
rect 562 3403 565 3446
rect 538 3363 549 3366
rect 570 3396 573 3406
rect 578 3403 581 3416
rect 586 3396 589 3486
rect 594 3413 597 3873
rect 618 3813 621 3936
rect 642 3933 645 3956
rect 650 3943 669 3946
rect 626 3893 629 3926
rect 650 3923 653 3943
rect 658 3873 661 3936
rect 666 3933 669 3943
rect 666 3863 669 3926
rect 674 3923 677 4016
rect 714 3953 717 4016
rect 690 3923 693 3936
rect 698 3893 701 3926
rect 706 3873 709 3936
rect 730 3933 733 4016
rect 746 3943 765 3946
rect 714 3913 717 3926
rect 730 3923 741 3926
rect 746 3923 749 3943
rect 626 3813 629 3826
rect 666 3813 669 3826
rect 602 3803 621 3806
rect 602 3723 605 3803
rect 642 3786 645 3806
rect 634 3783 645 3786
rect 618 3733 621 3746
rect 618 3693 621 3726
rect 634 3643 637 3783
rect 722 3733 725 3816
rect 658 3706 661 3726
rect 714 3706 717 3726
rect 658 3703 669 3706
rect 602 3493 605 3636
rect 610 3443 613 3526
rect 618 3503 621 3606
rect 626 3533 629 3606
rect 634 3596 637 3616
rect 642 3603 645 3616
rect 650 3613 653 3696
rect 666 3646 669 3703
rect 706 3703 717 3706
rect 706 3656 709 3703
rect 730 3686 733 3896
rect 754 3893 757 3936
rect 762 3933 765 3943
rect 762 3843 765 3926
rect 770 3906 773 3926
rect 778 3923 781 4016
rect 850 4013 853 4026
rect 858 4006 861 4016
rect 890 4013 893 4026
rect 810 3993 813 4006
rect 834 3976 837 4006
rect 850 4003 861 4006
rect 834 3973 845 3976
rect 786 3933 789 3966
rect 770 3903 777 3906
rect 786 3903 789 3926
rect 802 3916 805 3936
rect 818 3926 821 3946
rect 826 3933 829 3956
rect 798 3913 805 3916
rect 810 3913 813 3926
rect 818 3923 829 3926
rect 754 3813 757 3826
rect 738 3763 741 3806
rect 762 3803 765 3816
rect 774 3796 777 3903
rect 798 3846 801 3913
rect 810 3876 813 3896
rect 810 3873 817 3876
rect 798 3843 805 3846
rect 794 3813 797 3826
rect 802 3813 805 3843
rect 770 3793 777 3796
rect 738 3733 741 3756
rect 722 3683 733 3686
rect 658 3643 669 3646
rect 658 3613 661 3643
rect 650 3596 653 3606
rect 674 3603 677 3626
rect 682 3613 685 3656
rect 706 3653 717 3656
rect 634 3593 653 3596
rect 690 3583 693 3606
rect 698 3553 701 3616
rect 706 3603 709 3636
rect 714 3603 717 3653
rect 634 3543 653 3546
rect 634 3523 637 3543
rect 642 3523 645 3536
rect 650 3533 653 3543
rect 722 3533 725 3683
rect 746 3646 749 3726
rect 762 3656 765 3726
rect 770 3723 773 3793
rect 786 3733 789 3746
rect 738 3643 749 3646
rect 754 3653 765 3656
rect 730 3553 733 3606
rect 650 3483 653 3526
rect 642 3406 645 3426
rect 666 3413 669 3526
rect 698 3413 701 3526
rect 738 3496 741 3643
rect 754 3536 757 3653
rect 762 3593 765 3606
rect 770 3596 773 3616
rect 778 3603 781 3646
rect 794 3633 797 3806
rect 802 3723 805 3766
rect 814 3756 817 3873
rect 826 3853 829 3923
rect 834 3893 837 3936
rect 842 3923 845 3973
rect 850 3933 853 4003
rect 858 3933 861 3976
rect 850 3923 861 3926
rect 866 3903 869 3926
rect 842 3793 845 3806
rect 810 3753 817 3756
rect 810 3643 813 3753
rect 818 3683 821 3736
rect 842 3733 845 3746
rect 858 3733 861 3816
rect 826 3713 829 3726
rect 866 3646 869 3826
rect 874 3793 877 3996
rect 882 3933 885 3956
rect 914 3933 917 4006
rect 938 3993 941 4006
rect 954 4003 957 4016
rect 922 3943 941 3946
rect 890 3913 893 3926
rect 898 3923 909 3926
rect 922 3923 925 3943
rect 930 3893 933 3936
rect 938 3933 941 3943
rect 946 3943 965 3946
rect 978 3943 981 3956
rect 946 3933 949 3943
rect 938 3863 941 3926
rect 962 3923 965 3936
rect 970 3823 973 3936
rect 994 3933 997 4016
rect 1042 3993 1045 4006
rect 1002 3893 1005 3926
rect 898 3776 901 3796
rect 898 3773 905 3776
rect 874 3743 893 3746
rect 874 3723 877 3743
rect 882 3703 885 3736
rect 890 3733 893 3743
rect 890 3693 893 3726
rect 902 3686 905 3773
rect 914 3723 917 3816
rect 954 3813 973 3816
rect 938 3793 941 3806
rect 954 3803 957 3813
rect 954 3783 957 3796
rect 922 3743 925 3756
rect 970 3753 973 3806
rect 978 3793 981 3876
rect 1010 3833 1013 3936
rect 1034 3933 1037 3946
rect 1042 3943 1061 3946
rect 1018 3913 1021 3926
rect 1026 3873 1029 3926
rect 1042 3923 1045 3943
rect 1050 3923 1053 3936
rect 1058 3933 1061 3943
rect 1066 3903 1069 3926
rect 1074 3856 1077 4006
rect 1090 3926 1093 3966
rect 1098 3933 1101 4016
rect 1154 3996 1157 4016
rect 1178 4013 1181 4026
rect 1218 4013 1221 4026
rect 1146 3993 1157 3996
rect 1170 3993 1173 4006
rect 1106 3933 1109 3946
rect 1090 3923 1109 3926
rect 1074 3853 1081 3856
rect 986 3763 989 3806
rect 994 3793 997 3816
rect 898 3683 905 3686
rect 898 3666 901 3683
rect 826 3626 829 3646
rect 858 3643 869 3646
rect 890 3663 901 3666
rect 786 3613 789 3626
rect 802 3613 805 3626
rect 822 3623 829 3626
rect 786 3596 789 3606
rect 770 3593 789 3596
rect 810 3593 813 3616
rect 822 3576 825 3623
rect 842 3613 845 3626
rect 822 3573 829 3576
rect 778 3543 797 3546
rect 754 3533 765 3536
rect 730 3493 741 3496
rect 570 3393 589 3396
rect 522 3333 533 3336
rect 522 3313 525 3326
rect 530 3296 533 3333
rect 514 3293 533 3296
rect 506 3203 509 3216
rect 498 3163 509 3166
rect 474 3053 481 3056
rect 458 3013 461 3026
rect 478 2976 481 3053
rect 490 2993 493 3016
rect 498 3013 501 3026
rect 506 2986 509 3163
rect 514 3153 517 3293
rect 530 3213 533 3266
rect 522 3176 525 3196
rect 530 3186 533 3206
rect 538 3193 541 3363
rect 570 3356 573 3393
rect 566 3353 573 3356
rect 546 3213 549 3326
rect 566 3286 569 3353
rect 618 3343 621 3406
rect 642 3403 653 3406
rect 706 3403 709 3446
rect 634 3333 637 3396
rect 650 3356 653 3403
rect 714 3393 717 3416
rect 722 3383 725 3406
rect 730 3366 733 3493
rect 746 3423 749 3526
rect 738 3403 741 3416
rect 730 3363 741 3366
rect 642 3353 653 3356
rect 642 3326 645 3353
rect 562 3283 569 3286
rect 530 3183 549 3186
rect 522 3173 533 3176
rect 530 3136 533 3173
rect 514 3133 533 3136
rect 514 3106 517 3133
rect 522 3113 525 3126
rect 514 3103 525 3106
rect 530 3103 533 3126
rect 514 3013 517 3096
rect 514 2996 517 3006
rect 522 3003 525 3103
rect 530 2996 533 3016
rect 514 2993 533 2996
rect 538 2993 541 3126
rect 546 3123 549 3183
rect 554 3113 557 3146
rect 546 3013 549 3026
rect 562 3023 565 3283
rect 578 3256 581 3326
rect 570 3253 581 3256
rect 618 3323 645 3326
rect 570 3203 573 3253
rect 586 3203 589 3236
rect 618 3226 621 3323
rect 658 3303 661 3336
rect 674 3236 677 3336
rect 674 3233 693 3236
rect 618 3223 625 3226
rect 610 3186 613 3216
rect 606 3183 613 3186
rect 578 3133 581 3156
rect 606 3116 609 3183
rect 622 3176 625 3223
rect 634 3213 637 3226
rect 666 3193 669 3216
rect 674 3213 677 3226
rect 690 3216 693 3233
rect 686 3213 693 3216
rect 618 3173 625 3176
rect 606 3113 613 3116
rect 610 3093 613 3113
rect 506 2983 517 2986
rect 474 2973 481 2976
rect 466 2933 469 2956
rect 474 2926 477 2973
rect 482 2933 485 2956
rect 498 2933 501 2946
rect 450 2923 461 2926
rect 474 2923 485 2926
rect 458 2903 461 2923
rect 418 2733 421 2756
rect 426 2733 429 2836
rect 378 2713 389 2716
rect 394 2713 397 2726
rect 242 2593 249 2596
rect 266 2593 269 2606
rect 338 2603 357 2606
rect 370 2596 373 2616
rect 378 2603 381 2616
rect 386 2613 389 2713
rect 418 2703 421 2726
rect 434 2713 437 2776
rect 442 2733 445 2756
rect 450 2703 453 2806
rect 466 2786 469 2816
rect 474 2793 477 2806
rect 458 2783 469 2786
rect 458 2723 461 2783
rect 482 2773 485 2923
rect 490 2803 493 2846
rect 498 2813 501 2926
rect 506 2813 509 2906
rect 514 2833 517 2983
rect 554 2923 557 3016
rect 506 2776 509 2796
rect 502 2773 509 2776
rect 474 2676 477 2746
rect 502 2696 505 2773
rect 502 2693 509 2696
rect 474 2673 485 2676
rect 506 2673 509 2693
rect 402 2613 405 2626
rect 386 2596 389 2606
rect 218 2573 237 2576
rect 106 2403 125 2406
rect 98 2393 109 2396
rect 106 2323 109 2393
rect 130 2386 133 2516
rect 162 2446 165 2526
rect 186 2503 189 2526
rect 162 2443 173 2446
rect 138 2413 141 2426
rect 122 2383 133 2386
rect 122 2286 125 2383
rect 138 2363 141 2406
rect 146 2393 149 2416
rect 154 2403 157 2416
rect 162 2413 165 2436
rect 170 2413 173 2443
rect 186 2413 189 2466
rect 202 2426 205 2526
rect 202 2423 213 2426
rect 122 2283 129 2286
rect 106 1946 109 2126
rect 114 2123 117 2216
rect 126 2176 129 2283
rect 154 2226 157 2336
rect 162 2323 165 2346
rect 170 2233 173 2396
rect 178 2333 181 2346
rect 186 2323 189 2366
rect 194 2313 197 2416
rect 210 2356 213 2423
rect 226 2413 229 2526
rect 202 2353 213 2356
rect 202 2336 205 2353
rect 202 2333 213 2336
rect 234 2326 237 2573
rect 246 2496 249 2593
rect 298 2533 301 2596
rect 370 2593 389 2596
rect 242 2493 249 2496
rect 242 2413 245 2493
rect 242 2396 245 2406
rect 250 2403 253 2476
rect 258 2396 261 2416
rect 242 2393 261 2396
rect 274 2356 277 2416
rect 282 2413 285 2526
rect 314 2376 317 2436
rect 322 2403 325 2456
rect 298 2373 317 2376
rect 274 2353 285 2356
rect 242 2343 261 2346
rect 242 2333 245 2343
rect 150 2223 157 2226
rect 126 2173 133 2176
rect 130 2056 133 2173
rect 150 2156 153 2223
rect 150 2153 157 2156
rect 138 2123 141 2136
rect 146 2113 149 2136
rect 126 2053 133 2056
rect 114 2013 117 2026
rect 126 1946 129 2053
rect 106 1943 113 1946
rect 126 1943 133 1946
rect 110 1896 113 1943
rect 122 1913 125 1926
rect 106 1893 113 1896
rect 82 1773 93 1776
rect 90 1733 93 1773
rect 106 1746 109 1893
rect 130 1856 133 1943
rect 146 1923 149 1946
rect 126 1853 133 1856
rect 114 1813 117 1826
rect 126 1776 129 1853
rect 126 1773 133 1776
rect 106 1743 121 1746
rect 74 1703 85 1706
rect 82 1236 85 1703
rect 118 1646 121 1743
rect 118 1643 125 1646
rect 114 1613 117 1626
rect 114 1523 117 1536
rect 122 1506 125 1643
rect 114 1503 125 1506
rect 114 1406 117 1503
rect 130 1456 133 1773
rect 154 1766 157 2153
rect 162 2133 165 2216
rect 178 2193 181 2206
rect 170 2113 173 2126
rect 162 1993 165 2016
rect 170 2013 173 2026
rect 178 1996 181 2136
rect 194 2133 197 2196
rect 194 2113 197 2126
rect 202 2103 205 2236
rect 210 2213 213 2326
rect 234 2323 245 2326
rect 218 2193 221 2316
rect 242 2303 245 2323
rect 250 2313 253 2336
rect 258 2323 261 2343
rect 218 2133 221 2146
rect 226 2126 229 2256
rect 266 2203 269 2336
rect 274 2333 277 2346
rect 282 2323 285 2353
rect 298 2253 301 2373
rect 306 2333 309 2366
rect 330 2356 333 2416
rect 338 2413 341 2426
rect 346 2413 349 2526
rect 378 2426 381 2526
rect 402 2426 405 2596
rect 418 2593 421 2636
rect 442 2613 445 2626
rect 482 2553 485 2673
rect 490 2613 501 2616
rect 506 2603 509 2666
rect 514 2613 517 2776
rect 522 2743 525 2886
rect 522 2713 525 2726
rect 538 2663 541 2786
rect 546 2623 549 2836
rect 554 2776 557 2886
rect 562 2783 565 3016
rect 570 3013 573 3056
rect 570 2996 573 3006
rect 578 3003 581 3016
rect 586 2996 589 3016
rect 570 2993 589 2996
rect 594 2923 597 3006
rect 602 2946 605 3026
rect 610 2963 613 3046
rect 618 3033 621 3173
rect 686 3156 689 3213
rect 686 3153 693 3156
rect 666 3133 677 3136
rect 626 3113 629 3126
rect 618 3003 621 3016
rect 626 3013 629 3106
rect 634 2996 637 3036
rect 642 3013 645 3026
rect 658 3013 661 3126
rect 666 3113 669 3126
rect 674 3103 677 3133
rect 682 3123 685 3136
rect 690 3076 693 3153
rect 686 3073 693 3076
rect 686 3006 689 3073
rect 618 2993 637 2996
rect 642 2993 645 3006
rect 602 2943 613 2946
rect 602 2913 605 2936
rect 610 2863 613 2943
rect 618 2873 621 2993
rect 658 2983 661 3006
rect 686 3003 693 3006
rect 690 2983 693 3003
rect 626 2943 629 2956
rect 698 2946 701 3356
rect 722 3323 725 3336
rect 738 3273 741 3363
rect 746 3333 749 3416
rect 754 3323 757 3416
rect 762 3413 765 3533
rect 778 3513 781 3543
rect 786 3523 789 3536
rect 794 3523 797 3543
rect 826 3536 829 3573
rect 842 3543 845 3566
rect 858 3536 861 3643
rect 874 3543 877 3576
rect 890 3563 893 3663
rect 906 3583 909 3596
rect 762 3396 765 3406
rect 770 3403 773 3416
rect 778 3396 781 3416
rect 794 3413 797 3466
rect 802 3413 805 3506
rect 818 3453 821 3536
rect 826 3533 837 3536
rect 826 3446 829 3526
rect 810 3443 829 3446
rect 762 3393 781 3396
rect 762 3313 765 3336
rect 706 3213 709 3226
rect 706 3196 709 3206
rect 714 3203 717 3216
rect 722 3196 725 3216
rect 706 3193 725 3196
rect 714 3133 717 3156
rect 730 3133 733 3206
rect 738 3133 741 3146
rect 706 3113 709 3126
rect 722 3103 725 3126
rect 738 3113 741 3126
rect 746 3086 749 3176
rect 730 3083 749 3086
rect 730 3066 733 3083
rect 726 3063 733 3066
rect 706 3003 709 3016
rect 726 3006 729 3063
rect 726 3003 733 3006
rect 570 2813 573 2836
rect 586 2793 589 2856
rect 626 2853 629 2936
rect 642 2933 645 2946
rect 666 2943 693 2946
rect 698 2943 709 2946
rect 666 2933 669 2943
rect 674 2933 685 2936
rect 634 2923 645 2926
rect 650 2913 653 2926
rect 674 2923 693 2926
rect 690 2896 693 2923
rect 682 2893 693 2896
rect 602 2793 605 2816
rect 610 2813 613 2826
rect 626 2813 629 2826
rect 642 2813 645 2866
rect 682 2836 685 2893
rect 650 2813 653 2836
rect 682 2833 693 2836
rect 658 2813 661 2826
rect 554 2773 573 2776
rect 554 2703 557 2726
rect 562 2713 565 2726
rect 570 2723 573 2773
rect 610 2766 613 2806
rect 634 2793 637 2806
rect 642 2766 645 2806
rect 666 2793 669 2806
rect 674 2803 677 2816
rect 682 2783 685 2806
rect 602 2763 613 2766
rect 626 2763 645 2766
rect 594 2693 597 2736
rect 522 2593 525 2606
rect 530 2583 533 2616
rect 538 2603 541 2616
rect 506 2533 509 2556
rect 378 2423 397 2426
rect 402 2423 413 2426
rect 378 2386 381 2416
rect 386 2393 389 2406
rect 394 2403 397 2423
rect 402 2393 405 2416
rect 378 2383 397 2386
rect 314 2353 333 2356
rect 290 2193 293 2206
rect 234 2133 245 2136
rect 218 2123 229 2126
rect 186 2003 189 2026
rect 194 2013 197 2036
rect 210 2013 213 2026
rect 194 1996 197 2006
rect 178 1993 197 1996
rect 218 1993 221 2006
rect 162 1903 165 1926
rect 170 1913 173 1926
rect 162 1813 165 1836
rect 170 1813 173 1826
rect 154 1763 161 1766
rect 138 1713 141 1726
rect 158 1686 161 1763
rect 170 1703 173 1726
rect 154 1683 161 1686
rect 154 1626 157 1683
rect 150 1623 157 1626
rect 150 1516 153 1623
rect 162 1583 165 1616
rect 170 1613 173 1626
rect 162 1523 165 1546
rect 178 1536 181 1986
rect 186 1933 189 1946
rect 194 1933 197 1993
rect 226 1956 229 2106
rect 242 2096 245 2126
rect 234 2093 245 2096
rect 234 1983 237 2093
rect 250 2086 253 2136
rect 258 2113 261 2166
rect 266 2133 269 2146
rect 274 2143 293 2146
rect 274 2123 277 2143
rect 282 2123 285 2136
rect 290 2133 293 2143
rect 242 2083 253 2086
rect 290 2083 293 2126
rect 242 2013 245 2083
rect 218 1953 229 1956
rect 186 1913 189 1926
rect 194 1923 205 1926
rect 210 1903 213 1946
rect 218 1896 221 1953
rect 234 1933 237 1956
rect 202 1893 221 1896
rect 202 1783 205 1893
rect 210 1796 213 1806
rect 218 1803 221 1836
rect 226 1796 229 1816
rect 210 1793 229 1796
rect 186 1713 189 1726
rect 226 1706 229 1786
rect 250 1763 253 1816
rect 234 1743 253 1746
rect 234 1733 237 1743
rect 218 1703 229 1706
rect 242 1703 245 1736
rect 250 1723 253 1743
rect 186 1613 189 1636
rect 202 1613 213 1616
rect 186 1593 189 1606
rect 194 1573 197 1606
rect 210 1583 213 1606
rect 178 1533 185 1536
rect 150 1513 157 1516
rect 130 1453 149 1456
rect 130 1413 133 1426
rect 114 1403 125 1406
rect 78 1233 85 1236
rect 78 1176 81 1233
rect 98 1226 101 1246
rect 90 1203 93 1226
rect 98 1223 109 1226
rect 122 1216 125 1403
rect 130 1313 133 1326
rect 78 1173 85 1176
rect 82 1133 85 1173
rect 98 1143 101 1216
rect 118 1213 125 1216
rect 138 1213 141 1226
rect 118 1146 121 1213
rect 130 1203 141 1206
rect 118 1143 125 1146
rect 114 1113 117 1126
rect 122 1096 125 1143
rect 114 1093 125 1096
rect 82 943 85 1006
rect 114 986 117 1093
rect 122 1013 125 1026
rect 114 983 121 986
rect 82 733 85 936
rect 106 676 109 976
rect 118 746 121 983
rect 130 966 133 1166
rect 146 973 149 1453
rect 154 1106 157 1513
rect 170 1426 173 1526
rect 162 1423 173 1426
rect 182 1416 185 1533
rect 178 1413 185 1416
rect 162 1303 165 1326
rect 170 1313 173 1326
rect 170 1213 173 1256
rect 162 1123 165 1206
rect 170 1193 173 1206
rect 178 1163 181 1413
rect 194 1243 197 1566
rect 218 1563 221 1703
rect 258 1656 261 1966
rect 266 1813 269 1926
rect 274 1913 277 1956
rect 282 1783 285 2036
rect 298 2013 301 2126
rect 314 2103 317 2353
rect 322 2333 325 2346
rect 322 2306 325 2326
rect 338 2323 341 2376
rect 346 2343 365 2346
rect 346 2333 349 2343
rect 354 2313 357 2336
rect 362 2323 365 2343
rect 322 2303 333 2306
rect 330 2236 333 2303
rect 370 2296 373 2346
rect 322 2233 333 2236
rect 362 2293 373 2296
rect 362 2236 365 2293
rect 362 2233 373 2236
rect 322 2213 325 2233
rect 370 2213 373 2233
rect 322 2176 325 2196
rect 322 2173 333 2176
rect 330 2096 333 2173
rect 346 2113 349 2136
rect 362 2133 365 2146
rect 378 2133 381 2336
rect 386 2213 389 2306
rect 394 2263 397 2383
rect 410 2233 413 2423
rect 418 2413 421 2426
rect 434 2413 437 2526
rect 426 2393 429 2406
rect 450 2403 453 2416
rect 458 2413 461 2466
rect 466 2413 477 2416
rect 434 2306 437 2326
rect 458 2313 461 2406
rect 482 2403 485 2526
rect 546 2523 549 2616
rect 490 2403 493 2416
rect 434 2303 445 2306
rect 402 2196 405 2216
rect 410 2203 413 2226
rect 418 2196 421 2206
rect 402 2193 421 2196
rect 378 2103 381 2126
rect 322 2093 333 2096
rect 322 1986 325 2093
rect 386 2033 389 2176
rect 426 2156 429 2266
rect 442 2256 445 2303
rect 434 2253 445 2256
rect 434 2213 437 2253
rect 442 2176 445 2236
rect 474 2216 477 2236
rect 490 2223 493 2326
rect 498 2323 501 2506
rect 554 2426 557 2686
rect 570 2596 573 2606
rect 578 2603 581 2616
rect 586 2596 589 2616
rect 602 2613 605 2763
rect 610 2693 613 2726
rect 618 2703 621 2736
rect 626 2686 629 2763
rect 674 2756 677 2776
rect 690 2773 693 2833
rect 698 2766 701 2936
rect 670 2753 677 2756
rect 682 2763 701 2766
rect 618 2683 629 2686
rect 570 2593 589 2596
rect 594 2523 597 2606
rect 602 2533 605 2556
rect 554 2423 573 2426
rect 506 2283 509 2416
rect 546 2403 549 2416
rect 554 2346 557 2416
rect 554 2343 561 2346
rect 514 2216 517 2336
rect 418 2153 429 2156
rect 434 2173 445 2176
rect 466 2213 477 2216
rect 490 2213 517 2216
rect 338 1993 341 2006
rect 322 1983 333 1986
rect 314 1886 317 1936
rect 314 1883 325 1886
rect 290 1813 293 1826
rect 266 1683 269 1726
rect 282 1666 285 1756
rect 306 1753 309 1826
rect 314 1796 317 1806
rect 322 1803 325 1883
rect 330 1823 333 1983
rect 362 1936 365 2016
rect 370 1983 373 2006
rect 378 1976 381 2016
rect 394 1996 397 2136
rect 402 2113 405 2126
rect 410 2003 413 2146
rect 418 2083 421 2153
rect 434 2133 437 2173
rect 466 2156 469 2213
rect 466 2153 473 2156
rect 458 2103 461 2126
rect 394 1993 401 1996
rect 378 1973 389 1976
rect 362 1933 373 1936
rect 362 1906 365 1926
rect 358 1903 365 1906
rect 358 1836 361 1903
rect 358 1833 365 1836
rect 330 1796 333 1816
rect 346 1813 349 1826
rect 314 1793 333 1796
rect 338 1793 341 1806
rect 314 1703 317 1766
rect 322 1706 325 1786
rect 330 1713 333 1726
rect 322 1703 333 1706
rect 282 1663 309 1666
rect 258 1653 269 1656
rect 226 1603 229 1616
rect 266 1596 269 1653
rect 282 1613 285 1626
rect 258 1593 269 1596
rect 210 1516 213 1536
rect 218 1533 221 1546
rect 210 1513 221 1516
rect 234 1513 237 1526
rect 210 1403 213 1436
rect 218 1413 221 1513
rect 242 1476 245 1576
rect 258 1573 261 1593
rect 250 1503 253 1526
rect 258 1523 261 1536
rect 274 1513 277 1536
rect 234 1473 245 1476
rect 210 1343 229 1346
rect 210 1333 213 1343
rect 218 1303 221 1336
rect 226 1323 229 1343
rect 186 1203 189 1226
rect 210 1213 213 1236
rect 226 1213 229 1226
rect 234 1206 237 1473
rect 250 1403 253 1416
rect 266 1403 269 1416
rect 306 1413 309 1663
rect 322 1613 325 1626
rect 314 1413 317 1426
rect 330 1366 333 1703
rect 346 1646 349 1806
rect 354 1656 357 1816
rect 362 1813 365 1833
rect 370 1803 373 1933
rect 378 1813 381 1973
rect 398 1886 401 1993
rect 426 1953 429 2016
rect 410 1933 421 1936
rect 434 1933 437 2006
rect 442 1926 445 2086
rect 450 1996 453 2016
rect 458 2003 461 2036
rect 470 2026 473 2153
rect 482 2123 485 2206
rect 522 2203 525 2226
rect 514 2123 517 2146
rect 530 2133 533 2336
rect 558 2296 561 2343
rect 554 2293 561 2296
rect 538 2213 541 2286
rect 554 2213 557 2293
rect 546 2193 549 2206
rect 554 2203 565 2206
rect 562 2126 565 2146
rect 558 2123 565 2126
rect 470 2023 477 2026
rect 466 1996 469 2006
rect 450 1993 469 1996
rect 410 1913 413 1926
rect 418 1923 429 1926
rect 438 1923 445 1926
rect 394 1883 401 1886
rect 386 1813 389 1826
rect 362 1723 365 1746
rect 370 1713 373 1726
rect 378 1693 381 1796
rect 394 1793 397 1883
rect 402 1823 421 1826
rect 402 1803 405 1823
rect 418 1813 421 1823
rect 410 1793 413 1806
rect 426 1803 429 1916
rect 438 1866 441 1923
rect 450 1913 453 1936
rect 458 1933 461 1946
rect 474 1926 477 2023
rect 482 2013 485 2086
rect 538 2066 541 2086
rect 534 2063 541 2066
rect 514 2013 517 2026
rect 498 1933 501 1966
rect 458 1883 461 1926
rect 466 1923 477 1926
rect 490 1923 501 1926
rect 466 1866 469 1923
rect 490 1906 493 1923
rect 434 1863 441 1866
rect 458 1863 469 1866
rect 474 1903 493 1906
rect 434 1746 437 1863
rect 442 1803 445 1846
rect 458 1806 461 1863
rect 474 1813 477 1903
rect 458 1803 469 1806
rect 482 1803 485 1896
rect 386 1743 405 1746
rect 386 1733 389 1743
rect 386 1673 389 1726
rect 394 1693 397 1736
rect 402 1723 405 1743
rect 410 1733 413 1746
rect 418 1743 437 1746
rect 354 1653 373 1656
rect 346 1643 357 1646
rect 338 1603 341 1616
rect 346 1593 349 1606
rect 354 1536 357 1643
rect 370 1613 373 1653
rect 418 1626 421 1743
rect 426 1703 429 1736
rect 450 1733 453 1756
rect 466 1746 469 1803
rect 498 1746 501 1806
rect 506 1763 509 1956
rect 514 1916 517 1936
rect 522 1933 525 2036
rect 534 1966 537 2063
rect 558 2046 561 2123
rect 570 2056 573 2423
rect 578 2403 581 2446
rect 594 2413 597 2446
rect 602 2406 605 2526
rect 594 2403 605 2406
rect 578 2313 581 2326
rect 594 2276 597 2403
rect 610 2356 613 2626
rect 618 2623 621 2683
rect 618 2603 621 2616
rect 590 2273 597 2276
rect 602 2353 613 2356
rect 578 2123 581 2216
rect 590 2176 593 2273
rect 590 2173 597 2176
rect 594 2113 597 2173
rect 602 2143 605 2353
rect 610 2323 613 2346
rect 618 2306 621 2526
rect 626 2506 629 2676
rect 634 2523 637 2656
rect 642 2513 645 2746
rect 670 2666 673 2753
rect 682 2676 685 2763
rect 690 2713 693 2726
rect 706 2723 709 2943
rect 682 2673 693 2676
rect 714 2673 717 2936
rect 722 2743 725 2986
rect 730 2963 733 3003
rect 730 2923 733 2936
rect 738 2933 741 3076
rect 746 3013 749 3026
rect 754 3013 757 3306
rect 770 3303 773 3326
rect 770 3276 773 3296
rect 766 3273 773 3276
rect 766 3206 769 3273
rect 766 3203 773 3206
rect 778 3203 781 3336
rect 786 3293 789 3326
rect 810 3313 813 3443
rect 834 3426 837 3533
rect 826 3423 837 3426
rect 826 3386 829 3423
rect 834 3396 837 3416
rect 842 3403 845 3536
rect 858 3533 869 3536
rect 866 3436 869 3533
rect 858 3433 869 3436
rect 850 3413 853 3426
rect 850 3396 853 3406
rect 834 3393 853 3396
rect 826 3383 837 3386
rect 826 3333 829 3346
rect 770 3186 773 3203
rect 770 3183 781 3186
rect 770 3133 773 3166
rect 778 3113 781 3183
rect 786 3133 789 3206
rect 802 3196 805 3306
rect 818 3263 821 3326
rect 834 3216 837 3383
rect 850 3333 853 3346
rect 842 3313 845 3326
rect 798 3193 805 3196
rect 798 3136 801 3193
rect 810 3146 813 3216
rect 818 3196 821 3216
rect 826 3213 837 3216
rect 842 3213 845 3256
rect 858 3226 861 3433
rect 866 3413 869 3426
rect 874 3413 877 3446
rect 866 3313 869 3336
rect 874 3303 877 3406
rect 858 3223 865 3226
rect 826 3203 829 3213
rect 834 3196 837 3206
rect 818 3193 837 3196
rect 810 3143 817 3146
rect 798 3133 805 3136
rect 746 2993 749 3006
rect 762 2993 765 3006
rect 754 2956 757 2976
rect 770 2966 773 3106
rect 778 3003 781 3026
rect 802 3016 805 3133
rect 814 3086 817 3143
rect 814 3083 829 3086
rect 786 3003 789 3016
rect 794 3013 805 3016
rect 794 2973 797 3013
rect 802 2996 805 3006
rect 810 3003 813 3026
rect 818 2996 821 3016
rect 802 2993 821 2996
rect 750 2953 757 2956
rect 762 2963 773 2966
rect 730 2786 733 2836
rect 738 2803 741 2926
rect 750 2906 753 2953
rect 762 2913 765 2963
rect 750 2903 757 2906
rect 754 2833 757 2903
rect 778 2876 781 2966
rect 774 2873 781 2876
rect 746 2796 749 2816
rect 754 2803 757 2816
rect 762 2813 765 2856
rect 762 2796 765 2806
rect 746 2793 765 2796
rect 730 2783 741 2786
rect 670 2663 677 2666
rect 650 2613 653 2626
rect 658 2613 669 2616
rect 658 2556 661 2606
rect 654 2553 661 2556
rect 654 2506 657 2553
rect 666 2533 669 2546
rect 674 2533 677 2663
rect 690 2606 693 2673
rect 686 2603 693 2606
rect 686 2546 689 2603
rect 682 2543 689 2546
rect 626 2503 633 2506
rect 654 2503 661 2506
rect 630 2436 633 2503
rect 658 2486 661 2503
rect 682 2496 685 2543
rect 690 2513 693 2526
rect 698 2523 701 2586
rect 714 2553 717 2626
rect 722 2616 725 2726
rect 730 2713 733 2726
rect 738 2723 741 2783
rect 746 2696 749 2776
rect 774 2756 777 2873
rect 738 2693 749 2696
rect 754 2753 777 2756
rect 738 2636 741 2693
rect 754 2653 757 2753
rect 762 2743 781 2746
rect 762 2733 765 2743
rect 770 2703 773 2736
rect 778 2723 781 2743
rect 786 2736 789 2946
rect 826 2943 829 3083
rect 834 3013 837 3046
rect 842 3003 845 3146
rect 850 3123 853 3216
rect 862 3156 865 3223
rect 874 3193 877 3206
rect 858 3153 865 3156
rect 858 3073 861 3153
rect 882 3143 885 3536
rect 890 3523 893 3546
rect 898 3456 901 3576
rect 906 3543 909 3556
rect 890 3453 901 3456
rect 890 3296 893 3453
rect 906 3353 909 3536
rect 914 3506 917 3606
rect 922 3593 925 3726
rect 930 3716 933 3736
rect 930 3713 941 3716
rect 938 3656 941 3713
rect 962 3703 965 3726
rect 930 3653 941 3656
rect 922 3523 925 3586
rect 930 3573 933 3653
rect 946 3613 949 3636
rect 962 3603 965 3616
rect 962 3576 965 3596
rect 914 3503 921 3506
rect 918 3436 921 3503
rect 918 3433 925 3436
rect 914 3413 917 3426
rect 914 3326 917 3346
rect 922 3333 925 3433
rect 930 3403 933 3536
rect 938 3533 941 3546
rect 946 3523 949 3576
rect 962 3573 969 3576
rect 898 3313 901 3326
rect 906 3323 917 3326
rect 890 3293 901 3296
rect 898 3226 901 3293
rect 890 3223 901 3226
rect 890 3173 893 3223
rect 898 3136 901 3206
rect 914 3193 917 3246
rect 922 3213 925 3326
rect 938 3313 941 3326
rect 946 3276 949 3366
rect 938 3273 949 3276
rect 938 3216 941 3273
rect 938 3213 949 3216
rect 914 3143 917 3156
rect 882 3093 885 3136
rect 898 3133 909 3136
rect 898 3113 901 3126
rect 858 3013 861 3026
rect 866 3013 869 3036
rect 834 2993 845 2996
rect 850 2963 853 3006
rect 858 2953 861 3006
rect 866 2946 869 2976
rect 794 2813 797 2926
rect 826 2903 829 2936
rect 802 2813 805 2886
rect 834 2813 837 2826
rect 802 2743 805 2766
rect 786 2733 797 2736
rect 738 2633 749 2636
rect 722 2613 741 2616
rect 722 2593 733 2596
rect 706 2543 733 2546
rect 706 2533 709 2543
rect 682 2493 693 2496
rect 658 2483 677 2486
rect 626 2433 633 2436
rect 626 2406 629 2433
rect 634 2413 645 2416
rect 650 2413 653 2446
rect 626 2403 633 2406
rect 630 2346 633 2403
rect 642 2383 645 2413
rect 630 2343 637 2346
rect 626 2313 629 2326
rect 634 2306 637 2343
rect 614 2303 621 2306
rect 626 2303 637 2306
rect 614 2236 617 2303
rect 614 2233 621 2236
rect 610 2173 613 2216
rect 570 2053 577 2056
rect 558 2043 565 2046
rect 554 2013 557 2026
rect 534 1963 541 1966
rect 514 1913 521 1916
rect 518 1846 521 1913
rect 538 1906 541 1963
rect 514 1843 521 1846
rect 530 1903 541 1906
rect 466 1743 485 1746
rect 490 1743 501 1746
rect 434 1713 437 1726
rect 474 1713 477 1726
rect 402 1623 421 1626
rect 362 1583 365 1606
rect 370 1603 381 1606
rect 386 1556 389 1616
rect 402 1613 405 1623
rect 410 1613 421 1616
rect 342 1533 357 1536
rect 374 1553 389 1556
rect 342 1436 345 1533
rect 354 1513 357 1526
rect 374 1486 377 1553
rect 386 1523 389 1546
rect 394 1513 397 1526
rect 402 1506 405 1576
rect 338 1433 345 1436
rect 370 1483 377 1486
rect 394 1503 405 1506
rect 338 1386 341 1433
rect 370 1426 373 1483
rect 346 1393 349 1416
rect 354 1413 357 1426
rect 370 1423 377 1426
rect 338 1383 357 1386
rect 322 1363 333 1366
rect 290 1333 301 1336
rect 266 1293 269 1326
rect 242 1213 245 1246
rect 178 1133 181 1146
rect 210 1123 213 1206
rect 218 1203 237 1206
rect 218 1193 221 1203
rect 250 1196 253 1256
rect 274 1253 277 1326
rect 246 1193 253 1196
rect 246 1116 249 1193
rect 258 1123 261 1206
rect 274 1203 277 1216
rect 282 1213 285 1226
rect 298 1213 301 1326
rect 322 1306 325 1363
rect 338 1333 341 1346
rect 338 1313 341 1326
rect 322 1303 341 1306
rect 322 1213 325 1226
rect 298 1183 301 1206
rect 330 1176 333 1296
rect 306 1173 333 1176
rect 306 1156 309 1173
rect 338 1166 341 1303
rect 346 1203 349 1336
rect 354 1256 357 1383
rect 362 1363 365 1416
rect 374 1366 377 1423
rect 370 1363 377 1366
rect 362 1333 365 1356
rect 354 1253 365 1256
rect 302 1153 309 1156
rect 314 1163 341 1166
rect 246 1113 253 1116
rect 154 1103 161 1106
rect 158 1036 161 1103
rect 250 1046 253 1113
rect 250 1043 269 1046
rect 154 1033 161 1036
rect 130 963 149 966
rect 130 913 133 926
rect 130 813 133 826
rect 98 673 109 676
rect 114 743 121 746
rect 98 596 101 673
rect 98 593 109 596
rect 114 593 117 743
rect 146 733 149 963
rect 154 906 157 1033
rect 162 993 165 1016
rect 170 1013 173 1026
rect 186 1013 189 1026
rect 170 1003 181 1006
rect 162 923 165 936
rect 154 903 161 906
rect 158 836 161 903
rect 154 833 161 836
rect 122 706 125 726
rect 154 716 157 833
rect 170 823 173 926
rect 178 886 181 936
rect 186 933 189 946
rect 194 906 197 1006
rect 202 1003 205 1016
rect 210 993 213 1006
rect 210 936 213 956
rect 202 933 213 936
rect 218 933 221 1006
rect 234 946 237 1016
rect 234 943 245 946
rect 202 923 213 926
rect 194 903 205 906
rect 178 883 189 886
rect 178 816 181 836
rect 162 803 165 816
rect 170 813 181 816
rect 186 813 189 883
rect 178 796 181 806
rect 186 803 197 806
rect 202 796 205 903
rect 178 793 205 796
rect 178 733 181 746
rect 150 713 157 716
rect 122 703 129 706
rect 126 636 129 703
rect 150 646 153 713
rect 150 643 157 646
rect 122 633 129 636
rect 122 613 125 633
rect 138 603 141 616
rect 146 603 149 626
rect 82 203 85 576
rect 106 573 109 593
rect 130 513 133 526
rect 106 323 109 416
rect 130 333 133 406
rect 130 213 133 326
rect 154 313 157 643
rect 162 603 165 726
rect 170 613 173 626
rect 178 606 181 726
rect 202 723 205 793
rect 210 656 213 746
rect 202 653 213 656
rect 186 613 189 646
rect 162 523 165 546
rect 170 533 173 606
rect 178 603 189 606
rect 186 586 189 603
rect 186 583 197 586
rect 178 533 181 546
rect 194 533 197 583
rect 202 533 205 653
rect 218 646 221 926
rect 226 913 229 926
rect 234 923 237 936
rect 242 846 245 943
rect 250 923 253 936
rect 258 923 261 1016
rect 266 956 269 1043
rect 274 1013 277 1146
rect 302 1096 305 1153
rect 314 1106 317 1163
rect 362 1153 365 1253
rect 338 1133 365 1136
rect 322 1113 325 1126
rect 314 1103 325 1106
rect 302 1093 309 1096
rect 306 1026 309 1093
rect 302 1023 309 1026
rect 266 953 277 956
rect 266 906 269 936
rect 238 843 245 846
rect 258 903 269 906
rect 226 813 229 836
rect 238 776 241 843
rect 258 836 261 903
rect 250 833 261 836
rect 274 833 277 953
rect 302 946 305 1023
rect 282 923 285 936
rect 290 933 293 946
rect 302 943 309 946
rect 290 923 301 926
rect 306 916 309 943
rect 314 933 317 1016
rect 322 1013 325 1103
rect 322 943 325 1006
rect 290 913 309 916
rect 238 773 245 776
rect 242 743 245 773
rect 226 713 229 726
rect 218 643 229 646
rect 226 596 229 643
rect 250 633 253 833
rect 258 786 261 816
rect 258 783 269 786
rect 258 723 261 776
rect 266 733 269 783
rect 274 773 277 806
rect 290 786 293 913
rect 314 896 317 926
rect 330 923 333 1046
rect 338 1013 341 1133
rect 354 1026 357 1126
rect 362 1113 365 1126
rect 346 1023 357 1026
rect 346 1003 349 1023
rect 354 976 357 1016
rect 338 973 357 976
rect 338 913 341 973
rect 346 906 349 936
rect 354 933 357 966
rect 362 933 365 1016
rect 370 1013 373 1363
rect 378 1213 381 1346
rect 386 1333 389 1416
rect 394 1413 397 1503
rect 410 1463 413 1526
rect 418 1443 421 1556
rect 426 1526 429 1696
rect 434 1613 437 1636
rect 442 1613 445 1686
rect 450 1553 453 1666
rect 474 1613 477 1706
rect 482 1556 485 1743
rect 514 1666 517 1843
rect 530 1736 533 1903
rect 562 1886 565 2043
rect 574 1966 577 2053
rect 558 1883 565 1886
rect 570 1963 577 1966
rect 538 1746 541 1766
rect 538 1743 549 1746
rect 498 1663 517 1666
rect 522 1733 533 1736
rect 474 1553 485 1556
rect 434 1543 453 1546
rect 434 1533 437 1543
rect 442 1526 445 1536
rect 426 1523 445 1526
rect 450 1523 453 1543
rect 458 1533 461 1546
rect 394 1396 397 1406
rect 402 1403 405 1416
rect 410 1396 413 1416
rect 426 1413 429 1523
rect 466 1516 469 1526
rect 450 1513 469 1516
rect 450 1466 453 1513
rect 442 1463 453 1466
rect 394 1393 413 1396
rect 418 1393 421 1406
rect 402 1333 405 1346
rect 386 1233 389 1326
rect 386 1183 389 1216
rect 394 1203 397 1246
rect 402 1213 405 1226
rect 418 1203 421 1386
rect 434 1336 437 1446
rect 442 1386 445 1463
rect 474 1443 477 1553
rect 490 1546 493 1646
rect 482 1543 493 1546
rect 482 1523 485 1543
rect 442 1383 453 1386
rect 458 1383 461 1426
rect 434 1333 445 1336
rect 434 1243 437 1326
rect 442 1296 445 1333
rect 450 1313 453 1383
rect 442 1293 449 1296
rect 446 1236 449 1293
rect 458 1246 461 1366
rect 466 1323 469 1336
rect 474 1313 477 1336
rect 482 1323 485 1416
rect 490 1393 493 1536
rect 498 1516 501 1663
rect 506 1603 509 1656
rect 514 1533 517 1566
rect 522 1553 525 1733
rect 530 1653 533 1726
rect 546 1686 549 1743
rect 538 1683 549 1686
rect 538 1663 541 1683
rect 506 1523 517 1526
rect 498 1513 509 1516
rect 498 1363 501 1446
rect 490 1323 493 1336
rect 498 1306 501 1326
rect 490 1303 501 1306
rect 458 1243 465 1246
rect 446 1233 453 1236
rect 442 1213 445 1226
rect 386 1133 389 1146
rect 386 1026 389 1126
rect 386 1023 413 1026
rect 386 1013 389 1023
rect 378 1003 389 1006
rect 394 993 397 1006
rect 402 1003 405 1016
rect 370 933 373 956
rect 306 893 317 896
rect 322 903 349 906
rect 306 813 309 893
rect 322 816 325 903
rect 354 893 357 926
rect 362 923 373 926
rect 314 813 325 816
rect 330 813 333 856
rect 362 853 365 923
rect 386 906 389 926
rect 382 903 389 906
rect 382 836 385 903
rect 382 833 389 836
rect 282 783 293 786
rect 266 713 269 726
rect 250 613 253 626
rect 218 593 229 596
rect 162 393 165 416
rect 170 413 173 516
rect 186 446 189 526
rect 202 513 205 526
rect 178 443 189 446
rect 178 403 181 443
rect 194 416 197 426
rect 186 413 197 416
rect 186 393 189 406
rect 194 376 197 413
rect 202 403 205 416
rect 170 373 197 376
rect 162 213 165 326
rect 170 323 173 373
rect 194 353 197 373
rect 178 343 197 346
rect 178 333 181 343
rect 186 323 189 336
rect 194 323 197 343
rect 202 306 205 336
rect 210 333 213 536
rect 218 423 221 593
rect 226 533 229 546
rect 218 346 221 416
rect 218 343 229 346
rect 194 303 205 306
rect 74 123 77 186
rect 130 123 133 176
rect 170 173 173 216
rect 194 186 197 303
rect 210 213 213 326
rect 218 323 221 336
rect 226 313 229 343
rect 234 333 237 536
rect 250 466 253 596
rect 258 563 269 566
rect 258 533 261 563
rect 250 463 261 466
rect 258 396 261 463
rect 274 436 277 736
rect 282 643 285 783
rect 322 773 325 806
rect 330 803 341 806
rect 298 733 301 766
rect 354 763 357 806
rect 378 766 381 816
rect 386 813 389 833
rect 366 763 381 766
rect 346 713 349 726
rect 366 686 369 763
rect 378 703 381 726
rect 386 713 389 726
rect 362 683 369 686
rect 362 646 365 683
rect 282 593 285 616
rect 290 613 293 626
rect 298 613 301 646
rect 362 643 373 646
rect 314 596 317 606
rect 322 603 325 636
rect 330 596 333 616
rect 314 593 333 596
rect 338 593 341 606
rect 250 393 261 396
rect 270 433 277 436
rect 234 316 237 326
rect 242 323 245 336
rect 250 316 253 393
rect 270 356 273 433
rect 282 413 285 426
rect 306 406 309 536
rect 314 413 317 536
rect 338 533 341 556
rect 346 533 349 626
rect 354 553 357 636
rect 370 576 373 643
rect 394 623 397 916
rect 410 903 413 1023
rect 418 1013 421 1186
rect 434 1113 437 1126
rect 450 1043 453 1233
rect 462 1146 465 1243
rect 490 1236 493 1303
rect 490 1233 501 1236
rect 498 1213 501 1233
rect 506 1183 509 1513
rect 514 1503 517 1523
rect 522 1513 525 1526
rect 530 1433 533 1536
rect 538 1533 541 1546
rect 538 1483 541 1526
rect 522 1413 541 1416
rect 514 1316 517 1376
rect 522 1333 525 1413
rect 546 1373 549 1626
rect 558 1606 561 1883
rect 570 1643 573 1963
rect 578 1923 581 1946
rect 586 1913 589 1926
rect 602 1843 605 2126
rect 610 1926 613 1946
rect 618 1933 621 2233
rect 626 2133 629 2303
rect 642 2243 645 2356
rect 650 2313 653 2406
rect 658 2323 661 2466
rect 666 2413 669 2476
rect 674 2396 677 2483
rect 690 2426 693 2493
rect 682 2423 693 2426
rect 682 2403 685 2423
rect 706 2413 709 2526
rect 714 2503 717 2536
rect 738 2533 741 2613
rect 746 2566 749 2633
rect 754 2573 757 2606
rect 746 2563 757 2566
rect 690 2403 717 2406
rect 690 2396 693 2403
rect 674 2393 693 2396
rect 666 2353 669 2386
rect 722 2383 725 2416
rect 666 2343 685 2346
rect 666 2333 669 2343
rect 634 2196 637 2206
rect 642 2203 645 2226
rect 650 2196 653 2216
rect 674 2213 677 2336
rect 682 2323 685 2343
rect 690 2333 693 2346
rect 682 2296 685 2316
rect 682 2293 689 2296
rect 634 2193 653 2196
rect 634 2123 637 2146
rect 658 2143 661 2206
rect 666 2136 669 2206
rect 658 2133 669 2136
rect 634 2096 637 2116
rect 630 2093 637 2096
rect 630 2016 633 2093
rect 630 2013 637 2016
rect 626 1983 629 1996
rect 610 1923 621 1926
rect 626 1913 629 1926
rect 578 1813 581 1826
rect 610 1783 613 1816
rect 626 1813 629 1826
rect 634 1793 637 2013
rect 642 2003 645 2126
rect 658 2116 661 2133
rect 654 2113 661 2116
rect 654 2006 657 2113
rect 666 2103 669 2126
rect 674 2096 677 2206
rect 686 2156 689 2293
rect 698 2183 701 2326
rect 706 2293 709 2326
rect 714 2303 717 2346
rect 682 2153 689 2156
rect 682 2133 685 2153
rect 666 2093 677 2096
rect 666 2016 669 2093
rect 666 2013 673 2016
rect 654 2003 661 2006
rect 650 1966 653 1986
rect 646 1963 653 1966
rect 646 1836 649 1963
rect 658 1933 661 2003
rect 670 1966 673 2013
rect 682 1983 685 2126
rect 690 1993 693 2016
rect 698 2003 701 2146
rect 706 2093 709 2246
rect 722 2223 725 2326
rect 730 2296 733 2446
rect 738 2383 741 2496
rect 738 2313 741 2326
rect 730 2293 737 2296
rect 746 2293 749 2536
rect 754 2443 757 2563
rect 762 2413 765 2606
rect 770 2493 773 2676
rect 778 2556 781 2626
rect 786 2603 789 2696
rect 794 2683 797 2726
rect 810 2683 813 2806
rect 810 2656 813 2676
rect 802 2653 813 2656
rect 802 2596 805 2653
rect 802 2593 813 2596
rect 810 2573 813 2593
rect 778 2553 789 2556
rect 786 2466 789 2553
rect 810 2523 813 2556
rect 778 2463 789 2466
rect 754 2396 757 2406
rect 770 2403 773 2416
rect 754 2393 773 2396
rect 754 2323 757 2376
rect 770 2373 773 2393
rect 770 2313 773 2336
rect 734 2216 737 2293
rect 778 2266 781 2463
rect 794 2386 797 2406
rect 786 2383 797 2386
rect 786 2356 789 2383
rect 794 2373 805 2376
rect 786 2353 797 2356
rect 786 2333 789 2346
rect 794 2316 797 2353
rect 802 2323 805 2373
rect 810 2333 813 2376
rect 818 2333 821 2736
rect 826 2673 829 2746
rect 834 2733 837 2806
rect 826 2613 829 2636
rect 834 2583 837 2656
rect 842 2613 845 2936
rect 850 2843 853 2946
rect 858 2943 869 2946
rect 850 2813 853 2836
rect 858 2813 861 2943
rect 874 2936 877 3076
rect 906 3073 909 3133
rect 914 3123 917 3136
rect 922 3106 925 3206
rect 938 3183 941 3196
rect 946 3156 949 3213
rect 954 3206 957 3566
rect 966 3476 969 3573
rect 978 3556 981 3746
rect 1010 3743 1013 3806
rect 1018 3713 1021 3726
rect 1026 3613 1029 3626
rect 978 3553 1005 3556
rect 962 3473 969 3476
rect 962 3443 965 3473
rect 970 3393 973 3456
rect 978 3413 981 3536
rect 986 3473 989 3526
rect 1002 3453 1005 3553
rect 1034 3523 1037 3536
rect 1042 3486 1045 3756
rect 1050 3706 1053 3836
rect 1058 3813 1061 3826
rect 1078 3806 1081 3853
rect 1106 3843 1109 3923
rect 1090 3813 1093 3836
rect 1106 3813 1109 3826
rect 1074 3803 1081 3806
rect 1074 3783 1077 3803
rect 1058 3723 1061 3756
rect 1066 3713 1069 3726
rect 1050 3703 1057 3706
rect 1054 3636 1057 3703
rect 1034 3483 1045 3486
rect 1050 3633 1057 3636
rect 978 3363 981 3406
rect 986 3373 989 3396
rect 1034 3376 1037 3483
rect 1050 3426 1053 3633
rect 1058 3593 1061 3616
rect 1066 3613 1069 3626
rect 1074 3566 1077 3766
rect 1082 3733 1085 3746
rect 1082 3683 1085 3726
rect 1090 3716 1093 3736
rect 1106 3733 1109 3756
rect 1098 3723 1109 3726
rect 1114 3716 1117 3936
rect 1122 3803 1125 3926
rect 1130 3803 1133 3936
rect 1138 3886 1141 3926
rect 1146 3923 1149 3993
rect 1194 3983 1197 4006
rect 1138 3883 1149 3886
rect 1146 3836 1149 3883
rect 1138 3833 1149 3836
rect 1138 3776 1141 3833
rect 1170 3816 1173 3936
rect 1178 3913 1181 3936
rect 1186 3916 1189 3926
rect 1194 3923 1197 3936
rect 1202 3933 1205 3946
rect 1186 3913 1197 3916
rect 1202 3853 1205 3926
rect 1210 3906 1213 3936
rect 1218 3923 1221 3996
rect 1242 3933 1245 3956
rect 1274 3953 1277 4016
rect 1290 4013 1293 4026
rect 1282 3973 1285 4006
rect 1210 3903 1221 3906
rect 1218 3836 1221 3903
rect 1210 3833 1221 3836
rect 1146 3813 1173 3816
rect 1154 3793 1157 3806
rect 1130 3773 1141 3776
rect 1090 3713 1117 3716
rect 1122 3716 1125 3726
rect 1130 3716 1133 3773
rect 1162 3763 1165 3813
rect 1154 3736 1157 3746
rect 1138 3723 1141 3736
rect 1122 3713 1133 3716
rect 1090 3613 1093 3646
rect 1106 3596 1109 3606
rect 1114 3603 1117 3713
rect 1130 3636 1133 3713
rect 1130 3633 1141 3636
rect 1146 3633 1149 3736
rect 1154 3733 1165 3736
rect 1170 3733 1173 3796
rect 1162 3713 1165 3726
rect 1170 3723 1181 3726
rect 1138 3616 1141 3633
rect 1122 3596 1125 3616
rect 1138 3613 1149 3616
rect 1106 3593 1125 3596
rect 1130 3593 1133 3606
rect 1070 3563 1077 3566
rect 1070 3516 1073 3563
rect 1082 3523 1085 3556
rect 1114 3543 1133 3546
rect 1090 3523 1093 3536
rect 1070 3513 1077 3516
rect 1098 3513 1101 3526
rect 1106 3523 1109 3536
rect 1114 3533 1117 3543
rect 1074 3436 1077 3513
rect 1074 3433 1081 3436
rect 1050 3423 1061 3426
rect 1034 3373 1045 3376
rect 962 3223 965 3336
rect 986 3333 989 3356
rect 1010 3333 1013 3356
rect 962 3213 973 3216
rect 954 3203 965 3206
rect 938 3153 949 3156
rect 918 3103 925 3106
rect 866 2933 877 2936
rect 882 2933 885 3016
rect 898 3013 901 3056
rect 890 2983 893 3006
rect 906 2993 909 3016
rect 918 2976 921 3103
rect 930 3073 933 3136
rect 938 3096 941 3153
rect 946 3123 949 3146
rect 938 3093 949 3096
rect 946 3036 949 3093
rect 942 3033 949 3036
rect 918 2973 925 2976
rect 866 2836 869 2933
rect 874 2893 877 2926
rect 882 2913 885 2926
rect 866 2833 881 2836
rect 858 2793 861 2806
rect 866 2803 869 2826
rect 878 2756 881 2833
rect 878 2753 885 2756
rect 858 2733 861 2746
rect 850 2613 853 2646
rect 842 2603 853 2606
rect 826 2503 829 2526
rect 826 2403 829 2416
rect 794 2313 805 2316
rect 730 2213 737 2216
rect 730 2176 733 2213
rect 738 2193 749 2196
rect 714 2173 733 2176
rect 714 2106 717 2173
rect 730 2133 733 2156
rect 754 2123 757 2216
rect 762 2153 765 2266
rect 778 2263 785 2266
rect 770 2146 773 2256
rect 782 2176 785 2263
rect 762 2143 773 2146
rect 778 2173 785 2176
rect 714 2103 733 2106
rect 666 1963 673 1966
rect 666 1926 669 1963
rect 674 1943 693 1946
rect 674 1933 677 1943
rect 682 1926 685 1936
rect 658 1853 661 1926
rect 666 1923 685 1926
rect 690 1923 693 1943
rect 682 1896 685 1923
rect 674 1893 685 1896
rect 698 1896 701 1946
rect 706 1913 709 2016
rect 698 1893 709 1896
rect 646 1833 653 1836
rect 642 1736 645 1816
rect 578 1656 581 1726
rect 586 1663 589 1736
rect 594 1706 597 1726
rect 602 1723 605 1736
rect 634 1733 645 1736
rect 594 1703 601 1706
rect 578 1653 589 1656
rect 570 1613 573 1626
rect 558 1603 565 1606
rect 562 1543 565 1603
rect 586 1576 589 1653
rect 598 1636 601 1703
rect 634 1666 637 1733
rect 634 1663 645 1666
rect 578 1573 589 1576
rect 594 1633 601 1636
rect 554 1523 557 1536
rect 562 1533 573 1536
rect 562 1516 565 1526
rect 554 1513 565 1516
rect 530 1333 533 1366
rect 538 1333 541 1346
rect 514 1313 521 1316
rect 530 1313 533 1326
rect 518 1236 521 1313
rect 514 1233 521 1236
rect 514 1173 517 1233
rect 522 1156 525 1216
rect 530 1183 533 1206
rect 458 1143 465 1146
rect 506 1153 525 1156
rect 434 973 437 1006
rect 426 913 429 926
rect 450 913 453 996
rect 402 696 405 896
rect 434 813 437 826
rect 450 803 453 896
rect 458 856 461 1143
rect 466 1103 469 1126
rect 474 1113 477 1126
rect 466 923 469 1096
rect 490 1093 493 1126
rect 506 1116 509 1153
rect 514 1143 533 1146
rect 514 1133 517 1143
rect 474 993 477 1086
rect 482 1013 485 1026
rect 474 943 493 946
rect 474 933 477 943
rect 458 853 477 856
rect 474 806 477 853
rect 482 823 485 936
rect 490 923 493 943
rect 498 933 501 1116
rect 506 1113 513 1116
rect 510 1036 513 1113
rect 522 1103 525 1136
rect 530 1123 533 1143
rect 538 1083 541 1326
rect 546 1293 549 1326
rect 546 1193 549 1206
rect 506 1033 513 1036
rect 546 1033 549 1176
rect 554 1163 557 1506
rect 562 1493 565 1513
rect 562 1196 565 1426
rect 570 1203 573 1516
rect 578 1406 581 1573
rect 586 1503 589 1546
rect 594 1513 597 1633
rect 602 1593 605 1616
rect 610 1613 613 1626
rect 626 1613 629 1646
rect 642 1613 645 1663
rect 602 1506 605 1526
rect 594 1503 605 1506
rect 586 1413 589 1486
rect 594 1463 597 1503
rect 578 1403 585 1406
rect 582 1346 585 1403
rect 594 1383 597 1406
rect 582 1343 589 1346
rect 578 1253 581 1326
rect 578 1203 581 1216
rect 562 1193 581 1196
rect 554 1086 557 1156
rect 562 1113 565 1136
rect 570 1103 573 1136
rect 554 1083 565 1086
rect 578 1083 581 1193
rect 586 1093 589 1343
rect 602 1336 605 1496
rect 594 1333 605 1336
rect 610 1333 613 1606
rect 650 1556 653 1833
rect 658 1763 661 1836
rect 666 1796 669 1806
rect 674 1803 677 1893
rect 682 1796 685 1816
rect 666 1793 685 1796
rect 690 1783 693 1806
rect 666 1733 669 1746
rect 658 1596 661 1606
rect 666 1603 669 1616
rect 674 1596 677 1616
rect 658 1593 677 1596
rect 618 1506 621 1556
rect 650 1553 661 1556
rect 626 1543 645 1546
rect 626 1523 629 1543
rect 634 1513 637 1536
rect 642 1533 645 1543
rect 618 1503 625 1506
rect 622 1426 625 1503
rect 642 1436 645 1526
rect 658 1466 661 1553
rect 682 1533 685 1606
rect 690 1526 693 1776
rect 698 1696 701 1876
rect 706 1803 709 1893
rect 706 1713 709 1726
rect 698 1693 705 1696
rect 702 1616 705 1693
rect 618 1423 625 1426
rect 634 1433 645 1436
rect 650 1463 661 1466
rect 618 1393 621 1423
rect 594 1316 597 1333
rect 594 1313 605 1316
rect 602 1246 605 1313
rect 594 1243 605 1246
rect 594 1153 597 1243
rect 602 1213 605 1226
rect 618 1213 621 1326
rect 626 1303 629 1406
rect 634 1336 637 1433
rect 650 1413 653 1463
rect 674 1413 677 1526
rect 682 1523 693 1526
rect 698 1613 705 1616
rect 682 1493 685 1523
rect 650 1393 653 1406
rect 642 1343 645 1356
rect 634 1333 645 1336
rect 642 1313 645 1333
rect 642 1213 645 1226
rect 650 1206 653 1356
rect 594 1133 597 1146
rect 506 956 509 1033
rect 562 1026 565 1083
rect 602 1073 605 1206
rect 618 1193 621 1206
rect 642 1203 653 1206
rect 610 1066 613 1136
rect 618 1113 621 1126
rect 586 1063 613 1066
rect 514 993 517 1016
rect 522 1013 525 1026
rect 562 1023 573 1026
rect 506 953 517 956
rect 514 936 517 953
rect 530 946 533 1016
rect 538 996 541 1006
rect 546 1003 549 1016
rect 554 996 557 1016
rect 538 993 557 996
rect 510 933 517 936
rect 522 943 533 946
rect 510 866 513 933
rect 522 923 525 943
rect 530 923 533 936
rect 538 923 541 956
rect 554 933 557 956
rect 562 936 565 1006
rect 570 943 573 1023
rect 562 933 573 936
rect 510 863 517 866
rect 498 813 501 826
rect 474 803 485 806
rect 410 743 429 746
rect 410 733 413 743
rect 418 703 421 736
rect 426 723 429 743
rect 402 693 421 696
rect 418 646 421 693
rect 418 643 425 646
rect 362 573 373 576
rect 394 573 397 606
rect 422 596 425 643
rect 434 633 437 736
rect 458 716 461 736
rect 474 733 477 796
rect 482 733 485 803
rect 450 713 461 716
rect 450 666 453 713
rect 466 673 469 726
rect 450 663 461 666
rect 458 646 461 663
rect 458 643 465 646
rect 442 613 445 626
rect 418 593 425 596
rect 418 576 421 593
rect 462 576 465 643
rect 474 613 477 726
rect 482 646 485 726
rect 490 723 493 736
rect 498 696 501 746
rect 506 703 509 736
rect 514 713 517 863
rect 522 796 525 916
rect 530 806 533 816
rect 538 813 541 826
rect 546 806 549 816
rect 530 803 549 806
rect 522 793 533 796
rect 522 733 525 786
rect 530 716 533 793
rect 538 723 541 736
rect 546 733 549 803
rect 554 743 557 926
rect 562 913 565 926
rect 578 923 581 1006
rect 586 933 589 1063
rect 602 1023 621 1026
rect 594 933 597 1016
rect 562 796 565 806
rect 570 803 573 816
rect 578 796 581 816
rect 562 793 581 796
rect 586 793 589 806
rect 570 733 573 756
rect 546 723 565 726
rect 546 716 549 723
rect 530 713 549 716
rect 562 703 565 723
rect 498 693 509 696
rect 482 643 493 646
rect 482 613 485 626
rect 490 606 493 643
rect 482 603 493 606
rect 498 593 501 606
rect 402 573 421 576
rect 458 573 465 576
rect 322 446 325 526
rect 338 513 341 526
rect 322 443 333 446
rect 322 413 325 426
rect 330 406 333 443
rect 306 403 317 406
rect 322 403 333 406
rect 270 353 277 356
rect 234 313 253 316
rect 210 196 213 206
rect 218 203 221 216
rect 226 196 229 216
rect 210 193 229 196
rect 194 183 205 186
rect 234 183 237 306
rect 258 303 261 336
rect 266 286 269 336
rect 274 303 277 353
rect 282 333 285 376
rect 258 283 269 286
rect 250 213 253 226
rect 154 133 157 146
rect 178 133 181 146
rect 202 143 205 183
rect 226 113 229 126
rect 258 123 261 283
rect 266 133 269 216
rect 274 203 277 216
rect 282 213 285 316
rect 290 306 293 336
rect 298 333 301 396
rect 314 356 317 403
rect 338 393 341 406
rect 310 353 317 356
rect 346 356 349 416
rect 346 353 357 356
rect 310 306 313 353
rect 330 333 333 346
rect 354 323 357 353
rect 362 343 365 573
rect 402 556 405 573
rect 394 553 405 556
rect 394 506 397 553
rect 410 513 413 526
rect 442 523 445 556
rect 450 513 453 526
rect 458 523 461 573
rect 474 543 493 546
rect 474 533 477 543
rect 474 513 477 526
rect 394 503 405 506
rect 402 306 405 503
rect 410 413 413 426
rect 442 413 445 436
rect 450 413 453 426
rect 458 396 461 416
rect 466 413 469 446
rect 482 426 485 536
rect 490 523 493 543
rect 498 533 501 556
rect 506 466 509 693
rect 514 603 517 616
rect 522 573 525 606
rect 530 566 533 626
rect 538 603 541 616
rect 530 563 541 566
rect 514 516 517 536
rect 538 523 541 563
rect 546 553 549 606
rect 514 513 525 516
rect 498 463 509 466
rect 474 423 485 426
rect 418 333 421 356
rect 410 316 413 326
rect 426 316 429 336
rect 434 323 437 396
rect 450 393 461 396
rect 466 396 469 406
rect 474 403 477 423
rect 482 396 485 416
rect 490 403 493 436
rect 466 393 485 396
rect 450 333 453 393
rect 466 333 469 366
rect 498 353 501 463
rect 522 456 525 513
rect 546 483 549 536
rect 554 523 557 606
rect 514 453 525 456
rect 514 433 517 453
rect 410 313 437 316
rect 290 303 301 306
rect 310 303 317 306
rect 402 303 413 306
rect 298 206 301 303
rect 314 213 317 303
rect 290 203 301 206
rect 266 113 269 126
rect 290 53 293 203
rect 346 193 349 206
rect 354 136 357 216
rect 362 203 365 216
rect 378 213 381 256
rect 410 213 413 303
rect 426 213 429 236
rect 370 176 373 206
rect 418 203 429 206
rect 434 203 437 313
rect 450 253 453 326
rect 506 323 509 416
rect 530 393 533 406
rect 538 403 541 426
rect 546 403 549 416
rect 554 413 557 466
rect 562 366 565 696
rect 570 613 573 726
rect 578 713 581 766
rect 594 756 597 856
rect 602 803 605 1023
rect 618 1013 621 1023
rect 626 1006 629 1166
rect 634 1126 637 1176
rect 642 1133 645 1203
rect 658 1173 661 1376
rect 666 1336 669 1396
rect 674 1353 677 1406
rect 682 1373 685 1426
rect 666 1333 673 1336
rect 670 1266 673 1333
rect 682 1296 685 1356
rect 690 1333 693 1506
rect 682 1293 693 1296
rect 666 1263 673 1266
rect 634 1123 645 1126
rect 634 1013 637 1046
rect 610 993 613 1006
rect 626 1003 637 1006
rect 586 753 597 756
rect 586 723 589 753
rect 594 733 597 746
rect 602 693 605 736
rect 610 733 613 946
rect 618 913 621 926
rect 634 893 637 1003
rect 642 993 645 1036
rect 650 1013 653 1136
rect 666 1133 669 1263
rect 682 1166 685 1226
rect 690 1216 693 1293
rect 698 1223 701 1613
rect 706 1583 709 1596
rect 706 1463 709 1526
rect 714 1393 717 2026
rect 722 1993 725 2006
rect 722 1943 725 1966
rect 730 1956 733 2103
rect 738 1976 741 2016
rect 746 2003 749 2096
rect 754 1993 757 2026
rect 762 1976 765 2143
rect 738 1973 749 1976
rect 730 1953 737 1956
rect 722 1773 725 1936
rect 734 1876 737 1953
rect 730 1873 737 1876
rect 722 1523 725 1686
rect 722 1416 725 1516
rect 730 1423 733 1873
rect 746 1856 749 1973
rect 742 1853 749 1856
rect 758 1973 765 1976
rect 758 1856 761 1973
rect 770 1943 773 2006
rect 758 1853 765 1856
rect 742 1766 745 1853
rect 754 1813 757 1836
rect 738 1763 745 1766
rect 738 1706 741 1763
rect 746 1723 749 1746
rect 754 1713 757 1726
rect 738 1703 753 1706
rect 738 1483 741 1656
rect 750 1636 753 1703
rect 750 1633 757 1636
rect 746 1533 749 1616
rect 754 1603 757 1633
rect 754 1523 757 1546
rect 762 1516 765 1853
rect 770 1683 773 1916
rect 778 1766 781 2173
rect 794 2166 797 2296
rect 802 2263 805 2313
rect 818 2303 821 2326
rect 826 2323 829 2386
rect 818 2246 821 2296
rect 810 2243 821 2246
rect 794 2163 801 2166
rect 798 2086 801 2163
rect 810 2146 813 2243
rect 826 2226 829 2316
rect 834 2293 837 2566
rect 822 2223 829 2226
rect 822 2166 825 2223
rect 834 2193 837 2216
rect 842 2186 845 2596
rect 850 2483 853 2536
rect 858 2516 861 2726
rect 866 2613 869 2666
rect 866 2593 869 2606
rect 866 2533 869 2576
rect 874 2563 877 2676
rect 858 2513 865 2516
rect 862 2436 865 2513
rect 874 2503 877 2546
rect 858 2433 865 2436
rect 850 2293 853 2336
rect 850 2203 853 2286
rect 858 2243 861 2433
rect 866 2413 877 2416
rect 882 2413 885 2753
rect 890 2706 893 2966
rect 922 2946 925 2973
rect 942 2946 945 3033
rect 906 2933 909 2946
rect 922 2943 933 2946
rect 898 2723 901 2806
rect 890 2703 897 2706
rect 894 2636 897 2703
rect 890 2633 897 2636
rect 890 2506 893 2633
rect 898 2603 901 2616
rect 898 2523 901 2546
rect 890 2503 897 2506
rect 894 2436 897 2503
rect 890 2433 897 2436
rect 866 2373 869 2413
rect 882 2393 885 2406
rect 866 2333 869 2356
rect 866 2293 869 2326
rect 858 2233 869 2236
rect 858 2213 861 2233
rect 822 2163 829 2166
rect 810 2143 821 2146
rect 794 2083 801 2086
rect 786 2013 789 2046
rect 794 2003 797 2083
rect 802 2013 805 2026
rect 802 1936 805 2006
rect 794 1933 805 1936
rect 786 1803 789 1926
rect 794 1813 797 1836
rect 802 1813 805 1826
rect 794 1783 797 1806
rect 778 1763 789 1766
rect 786 1676 789 1763
rect 802 1713 805 1736
rect 778 1673 789 1676
rect 778 1626 781 1673
rect 778 1623 789 1626
rect 770 1533 773 1616
rect 786 1566 789 1623
rect 802 1616 805 1686
rect 810 1626 813 2126
rect 818 2116 821 2143
rect 826 2133 829 2163
rect 818 2113 825 2116
rect 822 1966 825 2113
rect 818 1963 825 1966
rect 834 1963 837 2186
rect 842 2183 853 2186
rect 818 1886 821 1963
rect 850 1956 853 2183
rect 866 2133 869 2196
rect 874 2183 877 2326
rect 882 2253 885 2386
rect 890 2316 893 2433
rect 898 2383 901 2416
rect 898 2333 901 2356
rect 890 2313 897 2316
rect 874 2133 877 2146
rect 866 2003 869 2126
rect 874 1983 877 2016
rect 882 1976 885 2246
rect 894 2236 897 2313
rect 890 2233 897 2236
rect 890 2113 893 2233
rect 898 2123 901 2216
rect 906 2123 909 2886
rect 930 2876 933 2943
rect 938 2943 945 2946
rect 938 2903 941 2943
rect 922 2873 933 2876
rect 914 2783 917 2796
rect 922 2673 925 2873
rect 938 2806 941 2866
rect 946 2833 949 2926
rect 954 2913 957 3016
rect 962 2996 965 3203
rect 978 3163 981 3196
rect 986 3013 989 3206
rect 994 3103 997 3226
rect 1002 3193 1005 3216
rect 1002 3113 1005 3126
rect 962 2993 973 2996
rect 986 2993 989 3006
rect 1002 2993 1005 3066
rect 962 2963 965 2993
rect 970 2883 973 2986
rect 842 1953 853 1956
rect 866 1973 885 1976
rect 826 1893 829 1946
rect 834 1933 837 1946
rect 842 1916 845 1953
rect 838 1913 845 1916
rect 818 1883 829 1886
rect 818 1803 821 1816
rect 818 1733 821 1756
rect 818 1643 821 1726
rect 826 1696 829 1883
rect 838 1826 841 1913
rect 838 1823 845 1826
rect 834 1733 837 1806
rect 834 1713 837 1726
rect 826 1693 833 1696
rect 830 1626 833 1693
rect 810 1623 821 1626
rect 802 1613 813 1616
rect 802 1603 813 1606
rect 778 1563 789 1566
rect 754 1493 757 1516
rect 762 1513 769 1516
rect 722 1413 733 1416
rect 738 1413 741 1466
rect 706 1323 709 1376
rect 738 1366 741 1406
rect 722 1363 741 1366
rect 722 1353 725 1363
rect 714 1333 717 1346
rect 714 1293 717 1326
rect 722 1276 725 1336
rect 718 1273 725 1276
rect 718 1216 721 1273
rect 690 1213 701 1216
rect 682 1163 697 1166
rect 650 993 653 1006
rect 666 1003 669 1126
rect 682 1036 685 1086
rect 694 1046 697 1163
rect 706 1123 709 1216
rect 718 1213 725 1216
rect 722 1196 725 1213
rect 730 1203 733 1326
rect 722 1193 733 1196
rect 694 1043 701 1046
rect 678 1033 685 1036
rect 678 966 681 1033
rect 690 1013 693 1026
rect 674 963 681 966
rect 698 966 701 1043
rect 706 1033 709 1086
rect 698 963 705 966
rect 658 913 661 926
rect 674 886 677 963
rect 674 883 693 886
rect 674 813 677 826
rect 626 793 629 806
rect 610 656 613 726
rect 618 676 621 746
rect 618 673 629 676
rect 578 593 581 606
rect 586 603 589 656
rect 602 653 613 656
rect 570 413 573 426
rect 578 403 581 536
rect 594 533 597 606
rect 602 603 605 653
rect 618 613 621 626
rect 626 613 629 673
rect 634 666 637 726
rect 658 666 661 796
rect 690 766 693 883
rect 702 836 705 963
rect 714 916 717 1156
rect 730 1086 733 1193
rect 722 1083 733 1086
rect 722 1003 725 1083
rect 730 1046 733 1066
rect 738 1053 741 1356
rect 746 1333 749 1416
rect 754 1353 757 1466
rect 766 1426 769 1513
rect 762 1423 769 1426
rect 762 1336 765 1423
rect 770 1373 773 1406
rect 778 1353 781 1563
rect 786 1533 789 1546
rect 786 1513 789 1526
rect 794 1463 797 1526
rect 794 1403 797 1426
rect 802 1403 805 1596
rect 818 1546 821 1623
rect 826 1623 833 1626
rect 826 1603 829 1623
rect 810 1543 821 1546
rect 786 1383 789 1396
rect 746 1313 749 1326
rect 754 1276 757 1336
rect 762 1333 773 1336
rect 750 1273 757 1276
rect 750 1146 753 1273
rect 770 1266 773 1333
rect 786 1323 789 1356
rect 794 1313 797 1376
rect 746 1143 753 1146
rect 762 1263 773 1266
rect 746 1123 749 1143
rect 762 1136 765 1263
rect 778 1193 781 1206
rect 802 1196 805 1396
rect 810 1373 813 1543
rect 818 1513 821 1536
rect 834 1526 837 1536
rect 842 1533 845 1823
rect 850 1803 853 1926
rect 858 1853 861 1936
rect 866 1933 869 1973
rect 890 1946 893 2016
rect 898 2013 901 2116
rect 906 2006 909 2116
rect 902 2003 909 2006
rect 902 1946 905 2003
rect 850 1733 853 1746
rect 850 1703 853 1726
rect 826 1503 829 1526
rect 834 1523 845 1526
rect 834 1443 837 1516
rect 842 1503 845 1523
rect 794 1193 805 1196
rect 794 1136 797 1193
rect 762 1133 769 1136
rect 730 1043 741 1046
rect 730 1003 733 1026
rect 738 1013 741 1043
rect 754 1023 757 1126
rect 766 1046 769 1133
rect 790 1133 797 1136
rect 790 1056 793 1133
rect 790 1053 797 1056
rect 762 1043 769 1046
rect 746 983 749 1006
rect 754 993 757 1016
rect 762 983 765 1043
rect 770 1003 773 1026
rect 770 993 781 996
rect 722 943 725 966
rect 762 943 765 956
rect 722 923 725 936
rect 786 926 789 1036
rect 794 933 797 1053
rect 802 1013 805 1126
rect 778 923 789 926
rect 714 913 725 916
rect 686 763 693 766
rect 698 833 705 836
rect 686 696 689 763
rect 674 676 677 696
rect 686 693 693 696
rect 698 693 701 833
rect 706 793 709 816
rect 714 813 717 826
rect 706 723 709 736
rect 674 673 681 676
rect 634 663 641 666
rect 658 663 669 666
rect 638 606 641 663
rect 658 613 661 626
rect 634 603 641 606
rect 602 526 605 546
rect 594 523 605 526
rect 610 543 629 546
rect 610 523 613 543
rect 618 523 621 536
rect 626 533 629 543
rect 634 526 637 603
rect 666 583 669 663
rect 678 576 681 673
rect 690 653 693 693
rect 674 573 681 576
rect 626 523 637 526
rect 594 513 597 523
rect 594 413 597 446
rect 626 443 629 523
rect 650 513 653 526
rect 658 523 669 526
rect 674 516 677 573
rect 706 553 709 606
rect 722 586 725 913
rect 778 836 781 923
rect 794 883 797 926
rect 738 813 741 836
rect 778 833 789 836
rect 754 796 757 806
rect 762 803 765 816
rect 770 796 773 816
rect 754 793 773 796
rect 778 793 781 806
rect 786 756 789 833
rect 802 813 805 1006
rect 810 933 813 1316
rect 818 1153 821 1436
rect 826 1333 829 1416
rect 842 1346 845 1466
rect 850 1433 853 1616
rect 858 1533 861 1766
rect 866 1753 869 1926
rect 874 1923 877 1946
rect 882 1943 893 1946
rect 898 1943 905 1946
rect 866 1533 869 1746
rect 874 1603 877 1896
rect 882 1763 885 1943
rect 890 1923 893 1936
rect 890 1743 893 1916
rect 898 1893 901 1943
rect 906 1873 909 1926
rect 914 1913 917 2606
rect 922 2563 925 2646
rect 922 2513 925 2536
rect 922 2376 925 2416
rect 930 2396 933 2806
rect 938 2803 949 2806
rect 938 2613 941 2796
rect 946 2763 949 2803
rect 946 2743 949 2756
rect 946 2613 949 2666
rect 954 2613 957 2876
rect 962 2813 965 2846
rect 938 2533 941 2546
rect 946 2513 949 2606
rect 930 2393 941 2396
rect 922 2373 933 2376
rect 922 2343 925 2366
rect 922 2003 925 2336
rect 930 2333 933 2373
rect 938 2326 941 2393
rect 934 2323 941 2326
rect 934 2226 937 2323
rect 930 2223 937 2226
rect 930 1996 933 2223
rect 938 2163 941 2206
rect 946 2203 949 2446
rect 954 2333 957 2526
rect 962 2403 965 2746
rect 970 2736 973 2816
rect 978 2743 981 2966
rect 970 2733 977 2736
rect 974 2676 977 2733
rect 974 2673 981 2676
rect 970 2603 973 2656
rect 970 2403 973 2596
rect 978 2543 981 2673
rect 986 2603 989 2986
rect 1010 2973 1013 3206
rect 1026 3203 1029 3216
rect 1034 3213 1037 3326
rect 1042 3196 1045 3373
rect 1026 3193 1045 3196
rect 1026 3116 1029 3193
rect 1034 3126 1037 3136
rect 1034 3123 1045 3126
rect 1026 3113 1037 3116
rect 1018 3013 1021 3056
rect 1034 3036 1037 3113
rect 1034 3033 1045 3036
rect 1018 2963 1021 3006
rect 1026 3003 1029 3016
rect 994 2913 997 2926
rect 994 2596 997 2906
rect 1010 2846 1013 2946
rect 1034 2923 1037 3016
rect 1002 2843 1013 2846
rect 1002 2803 1005 2843
rect 1002 2603 1005 2756
rect 1010 2746 1013 2816
rect 1018 2813 1021 2836
rect 1026 2753 1029 2826
rect 1034 2813 1037 2876
rect 1010 2743 1021 2746
rect 1010 2643 1013 2736
rect 1018 2673 1021 2743
rect 1026 2723 1029 2746
rect 1034 2723 1037 2736
rect 1026 2626 1029 2646
rect 1010 2623 1029 2626
rect 1010 2613 1021 2616
rect 1034 2613 1037 2706
rect 994 2593 1005 2596
rect 986 2536 989 2586
rect 978 2533 989 2536
rect 986 2523 997 2526
rect 978 2413 981 2476
rect 962 2306 965 2366
rect 970 2313 981 2316
rect 962 2303 973 2306
rect 954 2196 957 2216
rect 962 2203 965 2246
rect 970 2213 973 2303
rect 970 2196 973 2206
rect 954 2193 973 2196
rect 978 2193 981 2296
rect 962 2156 965 2176
rect 962 2153 969 2156
rect 938 2116 941 2136
rect 938 2113 945 2116
rect 926 1993 933 1996
rect 926 1906 929 1993
rect 942 1986 945 2113
rect 922 1903 929 1906
rect 938 1983 945 1986
rect 898 1803 901 1826
rect 882 1673 885 1736
rect 898 1733 901 1756
rect 906 1723 909 1856
rect 882 1613 885 1636
rect 906 1613 909 1626
rect 882 1533 885 1606
rect 858 1513 861 1526
rect 858 1363 861 1486
rect 874 1463 877 1526
rect 834 1333 837 1346
rect 842 1343 853 1346
rect 826 1283 829 1326
rect 850 1246 853 1343
rect 882 1316 885 1506
rect 890 1333 893 1606
rect 906 1526 909 1576
rect 914 1536 917 1806
rect 922 1803 925 1903
rect 930 1813 933 1836
rect 938 1803 941 1983
rect 954 1933 957 2126
rect 966 2026 969 2153
rect 978 2123 981 2146
rect 986 2116 989 2516
rect 994 2493 997 2523
rect 994 2203 997 2416
rect 1002 2403 1005 2593
rect 1010 2573 1013 2613
rect 1018 2543 1021 2606
rect 1042 2583 1045 3033
rect 1050 2736 1053 3416
rect 1058 3183 1061 3423
rect 1066 3413 1069 3426
rect 1078 3366 1081 3433
rect 1090 3413 1093 3436
rect 1090 3383 1093 3396
rect 1078 3363 1085 3366
rect 1082 3286 1085 3363
rect 1098 3336 1101 3406
rect 1074 3283 1085 3286
rect 1094 3333 1101 3336
rect 1114 3333 1117 3406
rect 1094 3286 1097 3333
rect 1094 3283 1101 3286
rect 1066 3203 1069 3226
rect 1058 3113 1061 3126
rect 1058 2853 1061 3076
rect 1066 3003 1069 3156
rect 1074 2823 1077 3283
rect 1098 3263 1101 3283
rect 1082 3163 1085 3256
rect 1090 3216 1093 3226
rect 1090 3213 1101 3216
rect 1090 3196 1093 3206
rect 1106 3203 1109 3326
rect 1114 3283 1117 3326
rect 1122 3226 1125 3536
rect 1130 3523 1133 3543
rect 1138 3533 1141 3556
rect 1146 3496 1149 3613
rect 1154 3536 1157 3616
rect 1178 3593 1181 3723
rect 1186 3703 1189 3736
rect 1194 3613 1197 3816
rect 1202 3813 1205 3826
rect 1202 3783 1205 3806
rect 1210 3803 1213 3833
rect 1202 3706 1205 3766
rect 1210 3723 1213 3736
rect 1218 3733 1221 3816
rect 1234 3813 1237 3926
rect 1250 3873 1253 3936
rect 1226 3793 1229 3806
rect 1226 3716 1229 3746
rect 1222 3713 1229 3716
rect 1202 3703 1213 3706
rect 1210 3636 1213 3703
rect 1206 3633 1213 3636
rect 1222 3636 1225 3713
rect 1222 3633 1229 3636
rect 1186 3573 1189 3606
rect 1154 3533 1165 3536
rect 1178 3533 1181 3566
rect 1186 3533 1189 3556
rect 1138 3493 1149 3496
rect 1138 3436 1141 3493
rect 1154 3463 1157 3526
rect 1162 3523 1165 3533
rect 1170 3523 1181 3526
rect 1186 3513 1189 3526
rect 1194 3483 1197 3596
rect 1206 3556 1209 3633
rect 1218 3603 1221 3616
rect 1226 3613 1229 3633
rect 1202 3553 1209 3556
rect 1138 3433 1149 3436
rect 1130 3393 1133 3416
rect 1146 3413 1149 3433
rect 1130 3323 1133 3346
rect 1138 3306 1141 3406
rect 1154 3326 1157 3416
rect 1170 3333 1173 3416
rect 1202 3346 1205 3553
rect 1210 3423 1213 3536
rect 1218 3533 1221 3576
rect 1234 3553 1237 3806
rect 1242 3793 1245 3816
rect 1258 3813 1261 3936
rect 1266 3913 1269 3936
rect 1274 3933 1277 3946
rect 1282 3883 1285 3946
rect 1290 3843 1293 3936
rect 1298 3933 1301 4016
rect 1330 4013 1333 4026
rect 1378 3993 1381 4006
rect 1394 3976 1397 4016
rect 1306 3943 1317 3946
rect 1298 3903 1301 3926
rect 1306 3836 1309 3943
rect 1322 3923 1325 3976
rect 1394 3973 1405 3976
rect 1330 3853 1333 3936
rect 1338 3933 1341 3966
rect 1338 3896 1341 3926
rect 1338 3893 1349 3896
rect 1346 3836 1349 3893
rect 1362 3883 1365 3936
rect 1306 3833 1321 3836
rect 1274 3773 1277 3806
rect 1242 3723 1245 3736
rect 1250 3713 1253 3736
rect 1258 3613 1261 3726
rect 1266 3703 1269 3726
rect 1274 3663 1277 3736
rect 1290 3733 1293 3746
rect 1298 3733 1301 3816
rect 1282 3713 1285 3726
rect 1306 3693 1309 3826
rect 1318 3776 1321 3833
rect 1342 3833 1349 3836
rect 1342 3776 1345 3833
rect 1354 3793 1357 3816
rect 1370 3803 1373 3926
rect 1378 3916 1381 3936
rect 1386 3933 1389 3946
rect 1402 3923 1405 3973
rect 1410 3943 1429 3946
rect 1410 3923 1413 3943
rect 1378 3913 1389 3916
rect 1386 3806 1389 3913
rect 1418 3863 1421 3936
rect 1426 3933 1429 3943
rect 1426 3913 1429 3926
rect 1450 3923 1453 4016
rect 1546 4013 1549 4026
rect 1458 3916 1461 3996
rect 1474 3993 1477 4006
rect 1498 3993 1501 4006
rect 1578 3986 1581 4016
rect 1586 4013 1589 4026
rect 1658 4013 1661 4026
rect 1578 3983 1589 3986
rect 1466 3923 1469 3936
rect 1450 3913 1461 3916
rect 1506 3913 1509 3936
rect 1402 3813 1405 3826
rect 1378 3803 1389 3806
rect 1378 3783 1381 3803
rect 1410 3783 1413 3816
rect 1442 3813 1445 3826
rect 1318 3773 1325 3776
rect 1306 3566 1309 3636
rect 1322 3613 1325 3773
rect 1338 3773 1345 3776
rect 1330 3616 1333 3726
rect 1338 3723 1341 3773
rect 1370 3743 1389 3746
rect 1370 3723 1373 3743
rect 1378 3723 1381 3736
rect 1386 3733 1389 3743
rect 1330 3613 1341 3616
rect 1330 3606 1333 3613
rect 1322 3603 1333 3606
rect 1330 3576 1333 3603
rect 1346 3586 1349 3646
rect 1378 3616 1381 3626
rect 1386 3616 1389 3726
rect 1402 3713 1405 3726
rect 1410 3723 1421 3726
rect 1442 3713 1445 3726
rect 1450 3696 1453 3913
rect 1458 3806 1461 3846
rect 1466 3823 1469 3886
rect 1514 3883 1517 3926
rect 1522 3903 1525 3936
rect 1538 3933 1541 3946
rect 1546 3933 1557 3936
rect 1530 3906 1533 3926
rect 1530 3903 1541 3906
rect 1530 3873 1533 3903
rect 1506 3813 1509 3836
rect 1458 3803 1465 3806
rect 1446 3693 1453 3696
rect 1362 3596 1365 3616
rect 1370 3603 1373 3616
rect 1378 3613 1389 3616
rect 1394 3613 1397 3626
rect 1402 3613 1413 3616
rect 1434 3613 1437 3626
rect 1378 3596 1381 3606
rect 1362 3593 1381 3596
rect 1346 3583 1357 3586
rect 1302 3563 1309 3566
rect 1218 3513 1221 3526
rect 1226 3503 1229 3536
rect 1234 3523 1237 3536
rect 1242 3523 1245 3536
rect 1250 3446 1253 3456
rect 1258 3446 1261 3536
rect 1282 3523 1285 3536
rect 1250 3443 1261 3446
rect 1186 3343 1205 3346
rect 1134 3303 1141 3306
rect 1146 3323 1157 3326
rect 1134 3226 1137 3303
rect 1114 3223 1125 3226
rect 1130 3223 1137 3226
rect 1114 3196 1117 3223
rect 1090 3193 1117 3196
rect 1082 3113 1085 3136
rect 1090 3133 1093 3193
rect 1106 3133 1117 3136
rect 1090 3083 1093 3126
rect 1106 3113 1109 3126
rect 1082 2983 1085 3046
rect 1090 3013 1101 3016
rect 1090 2963 1093 3006
rect 1058 2813 1077 2816
rect 1058 2803 1061 2813
rect 1066 2796 1069 2806
rect 1082 2803 1085 2916
rect 1090 2813 1093 2886
rect 1090 2796 1093 2806
rect 1066 2793 1093 2796
rect 1050 2733 1061 2736
rect 1050 2713 1053 2726
rect 1058 2706 1061 2733
rect 1054 2703 1061 2706
rect 1066 2703 1069 2736
rect 1074 2733 1077 2786
rect 1098 2776 1101 3006
rect 1106 2923 1109 3006
rect 1114 2933 1117 3036
rect 1122 2993 1125 3216
rect 1130 3043 1133 3223
rect 1146 3216 1149 3323
rect 1138 3213 1149 3216
rect 1154 3213 1157 3246
rect 1170 3206 1173 3256
rect 1186 3243 1189 3343
rect 1194 3323 1197 3336
rect 1186 3213 1189 3236
rect 1154 3203 1165 3206
rect 1170 3203 1189 3206
rect 1138 3166 1141 3186
rect 1138 3163 1145 3166
rect 1142 3026 1145 3163
rect 1138 3023 1145 3026
rect 1138 3003 1141 3023
rect 1154 3006 1157 3176
rect 1178 3133 1181 3146
rect 1170 3056 1173 3126
rect 1186 3056 1189 3203
rect 1162 3053 1173 3056
rect 1178 3053 1189 3056
rect 1162 3013 1165 3053
rect 1154 3003 1165 3006
rect 1170 3003 1173 3026
rect 1178 3013 1181 3053
rect 1122 2916 1125 2966
rect 1118 2913 1125 2916
rect 1106 2813 1109 2866
rect 1118 2846 1121 2913
rect 1114 2843 1121 2846
rect 1094 2773 1101 2776
rect 1094 2726 1097 2773
rect 1106 2733 1109 2806
rect 1114 2803 1117 2843
rect 1130 2826 1133 2926
rect 1138 2913 1141 2936
rect 1146 2883 1149 2996
rect 1162 2863 1165 3003
rect 1122 2813 1125 2826
rect 1130 2823 1149 2826
rect 1130 2813 1141 2816
rect 1154 2813 1157 2836
rect 1130 2753 1133 2813
rect 1138 2793 1141 2806
rect 1054 2636 1057 2703
rect 1050 2633 1057 2636
rect 1050 2593 1053 2633
rect 1058 2586 1061 2616
rect 1074 2603 1077 2726
rect 1082 2653 1085 2726
rect 1094 2723 1101 2726
rect 1138 2723 1141 2766
rect 1162 2746 1165 2856
rect 1170 2803 1173 2826
rect 1146 2743 1165 2746
rect 1058 2583 1069 2586
rect 1026 2536 1029 2566
rect 994 2133 997 2196
rect 1002 2123 1005 2306
rect 962 2023 969 2026
rect 978 2113 989 2116
rect 962 1933 965 2023
rect 970 1943 973 2006
rect 978 2003 981 2113
rect 986 2013 989 2076
rect 1010 2003 1013 2536
rect 1018 2533 1029 2536
rect 1018 2133 1021 2533
rect 1026 2416 1029 2526
rect 1034 2486 1037 2526
rect 1042 2523 1045 2576
rect 1050 2513 1053 2526
rect 1058 2503 1061 2536
rect 1066 2533 1069 2583
rect 1090 2533 1093 2576
rect 1076 2523 1086 2527
rect 1090 2486 1093 2526
rect 1034 2483 1045 2486
rect 1042 2426 1045 2483
rect 1082 2483 1093 2486
rect 1042 2423 1053 2426
rect 1026 2413 1037 2416
rect 1026 2316 1029 2406
rect 1034 2386 1037 2413
rect 1034 2383 1045 2386
rect 1034 2333 1037 2376
rect 1026 2313 1033 2316
rect 1030 2246 1033 2313
rect 1026 2243 1033 2246
rect 1018 2003 1021 2016
rect 994 1936 997 1966
rect 986 1933 997 1936
rect 946 1786 949 1816
rect 938 1783 949 1786
rect 922 1573 925 1706
rect 922 1543 925 1566
rect 930 1543 933 1606
rect 938 1593 941 1783
rect 954 1726 957 1926
rect 970 1883 973 1926
rect 986 1866 989 1933
rect 1010 1926 1013 1946
rect 1026 1933 1029 2243
rect 1034 2213 1037 2226
rect 1034 2133 1037 2196
rect 1042 2116 1045 2383
rect 1050 2253 1053 2423
rect 1058 2363 1061 2416
rect 1066 2403 1069 2416
rect 1058 2323 1061 2346
rect 1066 2256 1069 2376
rect 1074 2363 1077 2476
rect 1082 2443 1085 2483
rect 1090 2413 1093 2476
rect 1090 2333 1093 2346
rect 1062 2253 1069 2256
rect 1050 2133 1053 2246
rect 1062 2176 1065 2253
rect 1082 2213 1085 2226
rect 1062 2173 1069 2176
rect 1090 2173 1093 2326
rect 1098 2296 1101 2723
rect 1106 2616 1109 2656
rect 1106 2613 1117 2616
rect 1106 2563 1109 2606
rect 1106 2473 1109 2536
rect 1114 2513 1117 2613
rect 1122 2603 1125 2616
rect 1138 2593 1141 2656
rect 1146 2536 1149 2743
rect 1154 2653 1157 2726
rect 1162 2613 1165 2736
rect 1170 2733 1173 2756
rect 1178 2716 1181 2886
rect 1174 2713 1181 2716
rect 1174 2636 1177 2713
rect 1174 2633 1181 2636
rect 1154 2603 1165 2606
rect 1170 2603 1173 2616
rect 1154 2593 1157 2603
rect 1138 2523 1141 2536
rect 1146 2533 1165 2536
rect 1146 2523 1157 2526
rect 1114 2466 1117 2506
rect 1106 2463 1117 2466
rect 1106 2413 1109 2463
rect 1114 2403 1117 2446
rect 1122 2373 1125 2416
rect 1106 2313 1109 2336
rect 1098 2293 1105 2296
rect 1102 2226 1105 2293
rect 1098 2223 1105 2226
rect 1098 2193 1101 2223
rect 1106 2186 1109 2206
rect 1130 2203 1133 2426
rect 1138 2403 1141 2416
rect 1146 2263 1149 2496
rect 1154 2413 1157 2523
rect 1162 2476 1165 2533
rect 1162 2473 1169 2476
rect 1166 2406 1169 2473
rect 1162 2403 1169 2406
rect 1162 2323 1165 2403
rect 1178 2316 1181 2633
rect 1186 2333 1189 3046
rect 1194 2943 1197 3266
rect 1202 3116 1205 3336
rect 1210 3333 1213 3356
rect 1210 3253 1213 3326
rect 1218 3323 1221 3416
rect 1226 3333 1229 3346
rect 1250 3316 1253 3443
rect 1266 3403 1269 3416
rect 1274 3413 1277 3486
rect 1282 3393 1285 3406
rect 1242 3313 1253 3316
rect 1242 3246 1245 3313
rect 1234 3243 1245 3246
rect 1234 3173 1237 3243
rect 1242 3213 1245 3226
rect 1210 3133 1213 3146
rect 1226 3133 1229 3156
rect 1266 3153 1269 3346
rect 1282 3213 1285 3226
rect 1290 3166 1293 3556
rect 1302 3456 1305 3563
rect 1322 3553 1325 3576
rect 1330 3573 1349 3576
rect 1338 3506 1341 3566
rect 1298 3453 1305 3456
rect 1330 3503 1341 3506
rect 1298 3343 1301 3453
rect 1306 3426 1309 3446
rect 1330 3436 1333 3503
rect 1346 3483 1349 3573
rect 1354 3563 1357 3583
rect 1354 3533 1357 3556
rect 1362 3543 1381 3546
rect 1362 3523 1365 3543
rect 1370 3503 1373 3536
rect 1378 3533 1381 3543
rect 1330 3433 1341 3436
rect 1306 3423 1317 3426
rect 1314 3376 1317 3423
rect 1330 3403 1333 3416
rect 1338 3413 1341 3433
rect 1306 3373 1317 3376
rect 1306 3323 1309 3373
rect 1314 3313 1317 3326
rect 1306 3186 1309 3306
rect 1330 3303 1333 3376
rect 1338 3326 1341 3396
rect 1346 3373 1349 3446
rect 1362 3333 1365 3416
rect 1370 3403 1373 3496
rect 1378 3376 1381 3486
rect 1386 3443 1389 3613
rect 1446 3596 1449 3693
rect 1462 3686 1465 3803
rect 1458 3683 1465 3686
rect 1446 3593 1453 3596
rect 1450 3573 1453 3593
rect 1394 3523 1397 3536
rect 1402 3503 1405 3526
rect 1418 3503 1421 3556
rect 1458 3546 1461 3683
rect 1490 3636 1493 3806
rect 1514 3783 1517 3806
rect 1522 3793 1525 3816
rect 1538 3813 1541 3836
rect 1546 3826 1549 3926
rect 1562 3893 1565 3936
rect 1578 3933 1581 3956
rect 1586 3933 1589 3983
rect 1570 3903 1573 3926
rect 1586 3833 1589 3926
rect 1602 3923 1605 4006
rect 1546 3823 1581 3826
rect 1506 3656 1509 3726
rect 1482 3633 1493 3636
rect 1498 3653 1509 3656
rect 1482 3603 1485 3633
rect 1450 3543 1461 3546
rect 1434 3523 1437 3536
rect 1450 3496 1453 3543
rect 1450 3493 1461 3496
rect 1442 3413 1445 3426
rect 1394 3393 1397 3406
rect 1378 3373 1405 3376
rect 1370 3333 1373 3356
rect 1338 3323 1349 3326
rect 1354 3313 1357 3326
rect 1362 3303 1365 3326
rect 1378 3256 1381 3336
rect 1386 3333 1397 3336
rect 1362 3253 1381 3256
rect 1314 3196 1317 3206
rect 1322 3203 1325 3236
rect 1330 3196 1333 3216
rect 1314 3193 1333 3196
rect 1306 3183 1325 3186
rect 1290 3163 1297 3166
rect 1202 3113 1209 3116
rect 1206 2966 1209 3113
rect 1218 2986 1221 3106
rect 1226 2993 1229 3006
rect 1234 3003 1237 3026
rect 1242 2996 1245 3046
rect 1250 3013 1253 3126
rect 1294 3086 1297 3163
rect 1314 3133 1317 3146
rect 1322 3126 1325 3183
rect 1338 3163 1341 3206
rect 1290 3083 1297 3086
rect 1290 3043 1293 3083
rect 1306 3066 1309 3126
rect 1298 3063 1309 3066
rect 1314 3123 1325 3126
rect 1234 2993 1245 2996
rect 1218 2983 1229 2986
rect 1202 2963 1209 2966
rect 1194 2833 1197 2926
rect 1202 2826 1205 2963
rect 1210 2833 1213 2946
rect 1226 2883 1229 2983
rect 1234 2906 1237 2993
rect 1250 2983 1253 3006
rect 1242 2913 1245 2926
rect 1234 2903 1245 2906
rect 1250 2903 1253 2936
rect 1194 2813 1197 2826
rect 1202 2823 1217 2826
rect 1202 2733 1205 2816
rect 1214 2776 1217 2823
rect 1234 2813 1237 2826
rect 1242 2793 1245 2903
rect 1214 2773 1221 2776
rect 1154 2296 1157 2316
rect 1154 2293 1161 2296
rect 1158 2226 1161 2293
rect 1146 2213 1149 2226
rect 1154 2223 1161 2226
rect 1106 2183 1113 2186
rect 1038 2113 1045 2116
rect 1038 1956 1041 2113
rect 1038 1953 1045 1956
rect 986 1863 997 1866
rect 970 1803 973 1846
rect 970 1733 973 1776
rect 986 1733 989 1796
rect 994 1733 997 1863
rect 954 1723 973 1726
rect 978 1723 989 1726
rect 954 1713 965 1716
rect 970 1706 973 1723
rect 954 1703 973 1706
rect 946 1603 949 1626
rect 954 1586 957 1703
rect 962 1676 965 1696
rect 962 1673 969 1676
rect 950 1583 957 1586
rect 914 1533 925 1536
rect 898 1413 901 1526
rect 906 1523 917 1526
rect 906 1413 909 1426
rect 922 1383 925 1533
rect 930 1356 933 1526
rect 938 1413 941 1536
rect 950 1486 953 1583
rect 966 1566 969 1673
rect 978 1593 981 1666
rect 994 1626 997 1726
rect 1002 1693 1005 1926
rect 1010 1923 1017 1926
rect 1014 1836 1017 1923
rect 1034 1843 1037 1936
rect 1010 1833 1017 1836
rect 994 1623 1005 1626
rect 994 1573 997 1616
rect 962 1563 969 1566
rect 962 1533 965 1563
rect 950 1483 957 1486
rect 954 1463 957 1483
rect 946 1413 949 1426
rect 954 1403 957 1416
rect 962 1393 965 1526
rect 954 1366 957 1386
rect 954 1363 961 1366
rect 922 1353 933 1356
rect 874 1303 877 1316
rect 882 1313 889 1316
rect 842 1243 853 1246
rect 826 1213 829 1226
rect 842 1203 845 1243
rect 850 1213 861 1216
rect 866 1213 869 1226
rect 858 1156 861 1196
rect 834 1153 861 1156
rect 874 1153 877 1286
rect 886 1216 889 1313
rect 882 1213 889 1216
rect 834 1133 837 1153
rect 858 1133 861 1153
rect 834 1026 837 1126
rect 830 1023 837 1026
rect 818 926 821 1006
rect 830 966 833 1023
rect 842 973 845 1016
rect 850 1006 853 1106
rect 858 1013 861 1126
rect 874 1013 877 1026
rect 850 1003 861 1006
rect 830 963 837 966
rect 810 923 821 926
rect 770 753 789 756
rect 730 723 741 726
rect 746 723 749 736
rect 730 613 733 686
rect 746 603 749 616
rect 754 596 757 616
rect 762 603 765 636
rect 770 613 773 753
rect 786 743 805 746
rect 786 733 789 743
rect 794 723 797 736
rect 802 723 805 743
rect 770 596 773 606
rect 754 593 773 596
rect 714 583 725 586
rect 658 513 677 516
rect 690 513 693 526
rect 602 413 605 426
rect 610 413 613 436
rect 594 403 613 406
rect 642 403 645 416
rect 538 363 565 366
rect 538 346 541 363
rect 534 343 541 346
rect 442 213 445 226
rect 338 133 357 136
rect 362 173 373 176
rect 362 126 365 173
rect 434 133 437 146
rect 346 113 349 126
rect 354 123 365 126
rect 386 113 389 126
rect 458 123 461 206
rect 466 196 469 216
rect 474 203 477 216
rect 490 213 493 286
rect 482 196 485 206
rect 466 193 485 196
rect 498 123 501 216
rect 506 213 509 246
rect 506 193 509 206
rect 514 113 517 306
rect 534 296 537 343
rect 546 333 557 336
rect 546 306 549 333
rect 562 326 565 356
rect 554 323 565 326
rect 570 323 573 396
rect 578 333 581 346
rect 594 333 597 356
rect 546 303 557 306
rect 534 293 541 296
rect 522 203 525 256
rect 530 193 533 236
rect 538 213 541 293
rect 554 226 557 303
rect 586 283 589 326
rect 602 313 605 336
rect 610 323 613 403
rect 658 383 661 513
rect 618 333 621 346
rect 642 333 645 366
rect 546 223 557 226
rect 546 203 549 223
rect 578 203 581 226
rect 538 133 541 146
rect 562 133 565 146
rect 586 123 589 216
rect 594 163 597 306
rect 626 303 629 326
rect 666 323 669 426
rect 690 403 693 416
rect 706 393 709 486
rect 714 403 717 583
rect 738 496 741 556
rect 738 493 745 496
rect 730 423 733 486
rect 742 436 745 493
rect 762 486 765 586
rect 786 523 789 616
rect 794 573 797 596
rect 810 543 813 923
rect 818 733 821 876
rect 834 826 837 963
rect 850 923 853 946
rect 858 906 861 1003
rect 866 933 869 1006
rect 874 923 877 996
rect 850 903 861 906
rect 850 853 853 903
rect 826 823 837 826
rect 826 806 829 823
rect 834 813 845 816
rect 850 813 853 826
rect 826 803 837 806
rect 826 723 829 736
rect 834 716 837 803
rect 842 723 845 813
rect 850 753 853 796
rect 834 713 845 716
rect 818 603 821 706
rect 826 603 829 636
rect 834 613 837 626
rect 842 613 845 713
rect 834 603 845 606
rect 842 523 845 603
rect 850 516 853 746
rect 858 613 861 896
rect 866 803 869 826
rect 866 773 869 796
rect 866 713 869 756
rect 874 733 877 886
rect 882 743 885 1213
rect 890 1183 893 1196
rect 890 1103 893 1156
rect 898 1133 901 1336
rect 906 1213 909 1326
rect 914 1213 917 1336
rect 922 1333 925 1353
rect 890 923 893 1036
rect 898 1013 901 1126
rect 906 1086 909 1206
rect 922 1203 925 1326
rect 930 1303 933 1336
rect 930 1203 933 1216
rect 938 1196 941 1346
rect 926 1193 941 1196
rect 946 1193 949 1356
rect 958 1256 961 1363
rect 970 1323 973 1506
rect 978 1483 981 1536
rect 978 1403 981 1436
rect 986 1386 989 1466
rect 982 1383 989 1386
rect 982 1306 985 1383
rect 994 1323 997 1486
rect 1002 1316 1005 1623
rect 1010 1586 1013 1833
rect 1042 1826 1045 1953
rect 1038 1823 1045 1826
rect 1018 1793 1021 1816
rect 1018 1596 1021 1736
rect 1038 1726 1041 1823
rect 1026 1706 1029 1726
rect 1038 1723 1045 1726
rect 1026 1703 1033 1706
rect 1030 1626 1033 1703
rect 1026 1623 1033 1626
rect 1026 1603 1029 1623
rect 1018 1593 1029 1596
rect 1010 1583 1021 1586
rect 1010 1523 1013 1576
rect 1018 1503 1021 1583
rect 1010 1343 1013 1466
rect 1026 1446 1029 1593
rect 1042 1483 1045 1723
rect 1050 1716 1053 2126
rect 1066 2063 1069 2173
rect 1098 2133 1101 2146
rect 1110 2126 1113 2183
rect 1106 2123 1113 2126
rect 1058 1923 1061 1946
rect 1066 1933 1069 1996
rect 1058 1813 1061 1846
rect 1066 1823 1069 1926
rect 1066 1803 1069 1816
rect 1066 1733 1069 1796
rect 1074 1716 1077 2016
rect 1082 1923 1085 2036
rect 1082 1793 1085 1916
rect 1090 1843 1093 1946
rect 1098 1826 1101 2016
rect 1094 1823 1101 1826
rect 1094 1736 1097 1823
rect 1090 1733 1097 1736
rect 1106 1736 1109 2123
rect 1114 1963 1117 2006
rect 1122 2003 1125 2116
rect 1138 2026 1141 2186
rect 1154 2133 1157 2223
rect 1162 2126 1165 2206
rect 1154 2123 1165 2126
rect 1154 2106 1157 2123
rect 1170 2116 1173 2316
rect 1178 2313 1185 2316
rect 1182 2146 1185 2313
rect 1178 2143 1185 2146
rect 1178 2123 1181 2143
rect 1150 2103 1157 2106
rect 1162 2113 1173 2116
rect 1150 2046 1153 2103
rect 1150 2043 1157 2046
rect 1138 2023 1145 2026
rect 1114 1913 1117 1946
rect 1114 1753 1117 1826
rect 1106 1733 1113 1736
rect 1050 1713 1061 1716
rect 1058 1636 1061 1713
rect 1054 1633 1061 1636
rect 1070 1713 1077 1716
rect 1070 1636 1073 1713
rect 1082 1703 1085 1726
rect 1082 1643 1085 1666
rect 1070 1633 1077 1636
rect 1054 1566 1057 1633
rect 1066 1593 1069 1616
rect 1050 1563 1057 1566
rect 1050 1463 1053 1563
rect 1074 1546 1077 1633
rect 1090 1613 1093 1733
rect 1058 1523 1061 1546
rect 1074 1543 1081 1546
rect 1066 1496 1069 1536
rect 1058 1493 1069 1496
rect 1078 1466 1081 1543
rect 1074 1463 1081 1466
rect 1026 1443 1069 1446
rect 1018 1333 1021 1426
rect 1042 1423 1045 1436
rect 1026 1413 1037 1416
rect 1026 1356 1029 1413
rect 1034 1393 1037 1406
rect 1042 1403 1045 1416
rect 1026 1353 1037 1356
rect 1026 1333 1029 1346
rect 1034 1333 1037 1353
rect 954 1253 961 1256
rect 978 1303 985 1306
rect 994 1303 997 1316
rect 1002 1313 1013 1316
rect 906 1083 917 1086
rect 898 836 901 1006
rect 906 1003 909 1026
rect 906 933 909 996
rect 914 916 917 1083
rect 926 1026 929 1193
rect 910 913 917 916
rect 922 1023 929 1026
rect 922 913 925 1023
rect 930 993 933 1006
rect 938 983 941 1126
rect 946 976 949 1126
rect 954 1003 957 1253
rect 978 1236 981 1303
rect 966 1233 981 1236
rect 966 1176 969 1233
rect 978 1193 981 1216
rect 962 1173 969 1176
rect 962 1086 965 1173
rect 962 1083 973 1086
rect 930 973 949 976
rect 910 856 913 913
rect 910 853 917 856
rect 898 833 905 836
rect 890 813 893 826
rect 890 783 893 796
rect 902 776 905 833
rect 914 803 917 853
rect 922 803 925 886
rect 930 803 933 973
rect 962 966 965 1026
rect 970 986 973 1083
rect 978 1023 981 1186
rect 978 1003 981 1016
rect 970 983 977 986
rect 946 963 965 966
rect 946 926 949 963
rect 954 933 957 946
rect 938 923 949 926
rect 898 773 905 776
rect 874 673 877 726
rect 882 693 885 736
rect 890 646 893 726
rect 898 703 901 773
rect 866 633 877 636
rect 866 603 869 626
rect 874 613 877 633
rect 874 593 877 606
rect 858 533 861 576
rect 850 513 857 516
rect 762 483 773 486
rect 738 433 745 436
rect 706 366 709 386
rect 738 383 741 433
rect 754 413 757 456
rect 754 393 757 406
rect 706 363 713 366
rect 602 203 605 216
rect 610 213 613 226
rect 626 213 629 236
rect 634 213 637 246
rect 642 123 645 206
rect 658 183 661 206
rect 666 173 669 216
rect 674 203 677 316
rect 710 286 713 363
rect 738 333 741 346
rect 722 313 725 326
rect 762 323 765 416
rect 770 343 773 483
rect 778 413 781 466
rect 778 396 781 406
rect 786 403 789 416
rect 794 396 797 416
rect 818 413 821 446
rect 778 393 797 396
rect 802 326 805 406
rect 818 393 821 406
rect 826 353 829 416
rect 834 413 837 506
rect 842 363 845 466
rect 854 436 857 513
rect 866 463 869 546
rect 882 526 885 646
rect 890 643 901 646
rect 906 643 909 736
rect 914 716 917 736
rect 930 723 933 736
rect 914 713 921 716
rect 890 553 893 616
rect 898 603 901 643
rect 918 636 921 713
rect 938 693 941 916
rect 946 873 949 923
rect 946 733 949 816
rect 954 733 957 916
rect 962 793 965 946
rect 974 916 977 983
rect 986 933 989 1226
rect 994 1183 997 1286
rect 1010 1226 1013 1313
rect 1026 1303 1029 1316
rect 1002 1223 1013 1226
rect 994 1013 997 1126
rect 970 913 977 916
rect 970 893 973 913
rect 994 906 997 926
rect 986 903 997 906
rect 962 716 965 786
rect 970 733 973 876
rect 986 826 989 903
rect 986 823 997 826
rect 994 803 997 823
rect 1002 783 1005 1223
rect 1010 1193 1013 1206
rect 1026 1133 1029 1296
rect 1010 1006 1013 1026
rect 1010 1003 1021 1006
rect 1010 823 1013 936
rect 1010 803 1013 816
rect 1018 776 1021 1003
rect 1026 926 1029 1016
rect 1034 1013 1037 1036
rect 1034 933 1037 1006
rect 1042 996 1045 1326
rect 1050 1283 1053 1406
rect 1058 1323 1061 1416
rect 1066 1413 1069 1443
rect 1066 1333 1069 1406
rect 1074 1386 1077 1463
rect 1082 1403 1085 1446
rect 1074 1383 1081 1386
rect 1078 1326 1081 1383
rect 1074 1323 1081 1326
rect 1066 1213 1069 1226
rect 1074 1223 1077 1323
rect 1090 1313 1093 1516
rect 1098 1256 1101 1726
rect 1110 1666 1113 1733
rect 1106 1663 1113 1666
rect 1106 1643 1109 1663
rect 1122 1633 1125 1996
rect 1130 1616 1133 2016
rect 1142 1966 1145 2023
rect 1138 1963 1145 1966
rect 1138 1896 1141 1963
rect 1154 1923 1157 2043
rect 1162 2023 1165 2113
rect 1170 2076 1173 2096
rect 1170 2073 1181 2076
rect 1178 2016 1181 2073
rect 1194 2026 1197 2726
rect 1202 2573 1205 2676
rect 1210 2603 1213 2646
rect 1218 2573 1221 2773
rect 1250 2753 1253 2836
rect 1258 2746 1261 3036
rect 1274 3003 1277 3016
rect 1290 3013 1293 3026
rect 1298 2993 1301 3063
rect 1306 3003 1309 3036
rect 1314 3013 1317 3123
rect 1330 3113 1333 3126
rect 1338 3083 1341 3136
rect 1346 3133 1349 3246
rect 1362 3233 1365 3253
rect 1386 3246 1389 3326
rect 1370 3243 1389 3246
rect 1370 3203 1373 3243
rect 1378 3213 1381 3226
rect 1386 3213 1389 3236
rect 1346 3016 1349 3126
rect 1354 3113 1357 3136
rect 1378 3113 1381 3126
rect 1386 3123 1389 3146
rect 1370 3016 1373 3026
rect 1266 2843 1269 2936
rect 1274 2873 1277 2946
rect 1282 2933 1285 2956
rect 1322 2936 1325 3016
rect 1282 2823 1285 2926
rect 1290 2913 1293 2936
rect 1298 2933 1309 2936
rect 1314 2933 1325 2936
rect 1330 2933 1333 3016
rect 1338 3013 1349 3016
rect 1354 2996 1357 3016
rect 1362 3003 1365 3016
rect 1370 3013 1381 3016
rect 1386 3013 1389 3026
rect 1370 2996 1373 3006
rect 1354 2993 1373 2996
rect 1378 2986 1381 3013
rect 1362 2983 1381 2986
rect 1298 2883 1301 2926
rect 1314 2913 1317 2933
rect 1322 2903 1325 2926
rect 1234 2743 1261 2746
rect 1234 2656 1237 2743
rect 1242 2663 1245 2736
rect 1250 2676 1253 2726
rect 1250 2673 1261 2676
rect 1250 2656 1253 2673
rect 1226 2653 1237 2656
rect 1242 2653 1253 2656
rect 1226 2613 1229 2653
rect 1242 2613 1245 2653
rect 1202 2524 1205 2536
rect 1202 2486 1205 2516
rect 1202 2483 1209 2486
rect 1206 2336 1209 2483
rect 1218 2393 1221 2456
rect 1226 2423 1229 2596
rect 1234 2553 1237 2606
rect 1242 2496 1245 2526
rect 1238 2493 1245 2496
rect 1238 2416 1241 2493
rect 1226 2413 1241 2416
rect 1202 2333 1209 2336
rect 1202 2266 1205 2333
rect 1210 2283 1213 2316
rect 1202 2263 1209 2266
rect 1206 2146 1209 2263
rect 1202 2143 1209 2146
rect 1202 2093 1205 2143
rect 1218 2126 1221 2326
rect 1226 2183 1229 2413
rect 1234 2386 1237 2406
rect 1234 2383 1241 2386
rect 1238 2246 1241 2383
rect 1234 2243 1241 2246
rect 1210 2123 1221 2126
rect 1170 2013 1181 2016
rect 1190 2023 1197 2026
rect 1170 1943 1173 2013
rect 1190 1966 1193 2023
rect 1190 1963 1197 1966
rect 1186 1923 1189 1946
rect 1138 1893 1145 1896
rect 1142 1756 1145 1893
rect 1138 1753 1145 1756
rect 1138 1733 1141 1753
rect 1138 1623 1141 1726
rect 1154 1693 1157 1896
rect 1106 1603 1109 1616
rect 1106 1353 1109 1526
rect 1114 1416 1117 1616
rect 1122 1613 1133 1616
rect 1122 1523 1125 1613
rect 1130 1543 1133 1606
rect 1138 1526 1141 1616
rect 1134 1523 1141 1526
rect 1122 1503 1125 1516
rect 1122 1423 1125 1466
rect 1134 1436 1137 1523
rect 1134 1433 1141 1436
rect 1146 1433 1149 1646
rect 1162 1623 1165 1826
rect 1170 1696 1173 1876
rect 1186 1823 1189 1916
rect 1194 1893 1197 1963
rect 1202 1873 1205 2016
rect 1210 2013 1213 2123
rect 1186 1803 1189 1816
rect 1202 1813 1205 1846
rect 1178 1713 1181 1736
rect 1194 1733 1197 1806
rect 1210 1783 1213 1806
rect 1170 1693 1181 1696
rect 1178 1636 1181 1693
rect 1178 1633 1189 1636
rect 1154 1613 1165 1616
rect 1154 1523 1157 1613
rect 1162 1593 1165 1606
rect 1162 1503 1165 1536
rect 1170 1533 1173 1626
rect 1178 1603 1181 1616
rect 1186 1523 1189 1633
rect 1114 1413 1133 1416
rect 1130 1356 1133 1413
rect 1122 1353 1133 1356
rect 1122 1326 1125 1353
rect 1138 1346 1141 1433
rect 1146 1403 1149 1416
rect 1162 1383 1165 1406
rect 1186 1396 1189 1436
rect 1178 1393 1189 1396
rect 1178 1376 1181 1393
rect 1170 1373 1181 1376
rect 1106 1323 1125 1326
rect 1082 1253 1101 1256
rect 1074 1193 1077 1206
rect 1082 1186 1085 1253
rect 1090 1213 1093 1246
rect 1106 1223 1109 1316
rect 1122 1306 1125 1323
rect 1118 1303 1125 1306
rect 1118 1236 1121 1303
rect 1118 1233 1125 1236
rect 1098 1203 1101 1216
rect 1122 1213 1125 1233
rect 1130 1223 1133 1346
rect 1138 1343 1149 1346
rect 1138 1283 1141 1336
rect 1074 1183 1085 1186
rect 1050 1143 1061 1146
rect 1074 1133 1077 1183
rect 1082 1123 1085 1146
rect 1058 1013 1061 1026
rect 1074 1013 1077 1086
rect 1098 1036 1101 1196
rect 1090 1033 1101 1036
rect 1050 1003 1061 1006
rect 1042 993 1053 996
rect 1026 923 1037 926
rect 1002 773 1021 776
rect 954 713 965 716
rect 954 646 957 713
rect 970 703 973 716
rect 978 713 981 726
rect 994 723 997 746
rect 1002 716 1005 773
rect 1034 766 1037 923
rect 1050 836 1053 993
rect 1066 973 1069 1006
rect 1066 923 1069 936
rect 1026 763 1037 766
rect 1046 833 1053 836
rect 1010 733 1013 756
rect 1018 726 1021 736
rect 1010 723 1021 726
rect 1002 713 1013 716
rect 954 643 961 646
rect 914 633 921 636
rect 906 613 909 626
rect 914 613 917 633
rect 890 543 917 546
rect 890 533 893 543
rect 914 536 917 543
rect 874 513 877 526
rect 882 523 893 526
rect 854 433 861 436
rect 850 393 853 416
rect 858 386 861 433
rect 866 413 869 446
rect 890 443 893 523
rect 898 513 901 536
rect 914 533 925 536
rect 874 413 877 436
rect 866 393 869 406
rect 858 383 877 386
rect 802 323 821 326
rect 706 283 713 286
rect 682 193 685 206
rect 666 133 669 146
rect 690 123 693 216
rect 698 193 701 206
rect 706 203 709 283
rect 714 203 717 216
rect 722 213 725 306
rect 834 296 837 346
rect 858 323 861 356
rect 826 293 837 296
rect 730 203 733 216
rect 738 193 741 216
rect 762 213 765 236
rect 770 213 773 246
rect 786 223 789 286
rect 826 236 829 293
rect 858 276 861 306
rect 850 273 861 276
rect 826 233 837 236
rect 746 123 749 206
rect 778 203 789 206
rect 770 133 773 146
rect 794 123 797 216
rect 802 133 805 216
rect 810 196 813 206
rect 818 203 821 216
rect 826 196 829 216
rect 810 193 829 196
rect 834 143 837 233
rect 842 213 845 236
rect 850 213 853 273
rect 874 266 877 383
rect 906 366 909 446
rect 914 433 917 533
rect 930 526 933 636
rect 946 613 949 626
rect 958 586 961 643
rect 958 583 965 586
rect 946 533 949 556
rect 954 543 957 566
rect 866 263 877 266
rect 902 363 909 366
rect 850 123 853 206
rect 866 193 869 263
rect 902 256 905 363
rect 914 323 917 416
rect 922 413 925 526
rect 930 523 941 526
rect 902 253 909 256
rect 906 233 909 253
rect 874 203 877 226
rect 882 213 901 216
rect 882 203 885 213
rect 882 183 885 196
rect 890 193 893 206
rect 874 133 877 146
rect 906 123 909 216
rect 914 213 917 276
rect 922 253 925 346
rect 930 333 933 516
rect 938 453 941 523
rect 954 353 957 526
rect 962 513 965 583
rect 970 533 973 696
rect 970 503 973 516
rect 970 413 973 446
rect 970 366 973 406
rect 962 363 973 366
rect 938 323 941 346
rect 922 196 925 206
rect 930 203 933 246
rect 938 196 941 216
rect 946 203 949 336
rect 954 303 957 326
rect 962 243 965 363
rect 978 356 981 596
rect 986 503 989 566
rect 994 523 997 696
rect 1026 623 1029 763
rect 1034 733 1037 756
rect 1046 746 1049 833
rect 1046 743 1053 746
rect 1034 703 1037 726
rect 1010 603 1013 616
rect 1042 586 1045 726
rect 1050 593 1053 743
rect 1058 693 1061 826
rect 1074 816 1077 966
rect 1090 946 1093 1033
rect 1106 1003 1109 1026
rect 1114 996 1117 1086
rect 1122 1013 1125 1126
rect 1130 1083 1133 1196
rect 1110 993 1117 996
rect 1090 943 1101 946
rect 1090 906 1093 926
rect 1086 903 1093 906
rect 1086 826 1089 903
rect 1086 823 1093 826
rect 1098 823 1101 943
rect 1110 836 1113 993
rect 1130 986 1133 1026
rect 1122 983 1133 986
rect 1122 923 1125 983
rect 1130 923 1133 936
rect 1106 833 1113 836
rect 1066 813 1077 816
rect 1066 633 1069 813
rect 1074 803 1085 806
rect 1090 803 1093 823
rect 1098 773 1101 816
rect 1106 756 1109 833
rect 1102 753 1109 756
rect 1074 733 1077 746
rect 1082 723 1085 736
rect 1066 606 1069 626
rect 1090 613 1093 736
rect 1058 603 1069 606
rect 1082 603 1093 606
rect 1042 583 1053 586
rect 1002 523 1005 536
rect 1010 506 1013 536
rect 1026 533 1037 536
rect 1042 533 1045 566
rect 1050 526 1053 583
rect 1002 503 1013 506
rect 1002 446 1005 503
rect 1018 463 1021 526
rect 1034 513 1037 526
rect 1042 523 1053 526
rect 1058 523 1061 603
rect 1102 596 1105 753
rect 1114 673 1117 816
rect 1122 733 1125 776
rect 1138 773 1141 1216
rect 1146 1203 1149 1343
rect 1154 1166 1157 1366
rect 1170 1226 1173 1373
rect 1194 1293 1197 1696
rect 1202 1563 1205 1746
rect 1210 1613 1213 1756
rect 1218 1716 1221 2096
rect 1226 2003 1229 2126
rect 1234 2106 1237 2243
rect 1250 2213 1253 2576
rect 1258 2496 1261 2586
rect 1266 2533 1269 2796
rect 1274 2706 1277 2756
rect 1282 2723 1285 2816
rect 1298 2813 1301 2866
rect 1298 2773 1301 2806
rect 1290 2733 1293 2756
rect 1298 2723 1301 2736
rect 1306 2706 1309 2876
rect 1330 2836 1333 2926
rect 1338 2863 1341 2946
rect 1346 2923 1349 2936
rect 1354 2933 1357 2956
rect 1314 2833 1333 2836
rect 1314 2773 1317 2833
rect 1362 2816 1365 2983
rect 1370 2933 1381 2936
rect 1378 2913 1381 2926
rect 1386 2923 1389 2956
rect 1394 2916 1397 3326
rect 1402 3243 1405 3373
rect 1418 3263 1421 3396
rect 1458 3376 1461 3493
rect 1446 3373 1461 3376
rect 1446 3296 1449 3373
rect 1466 3336 1469 3446
rect 1474 3393 1477 3486
rect 1482 3443 1485 3576
rect 1498 3553 1501 3653
rect 1514 3576 1517 3696
rect 1522 3683 1525 3756
rect 1530 3676 1533 3806
rect 1538 3793 1541 3806
rect 1546 3693 1549 3823
rect 1570 3723 1573 3816
rect 1578 3813 1581 3823
rect 1602 3813 1605 3906
rect 1618 3853 1621 3926
rect 1626 3883 1629 3926
rect 1634 3876 1637 3936
rect 1642 3923 1645 4006
rect 1650 3933 1653 3956
rect 1666 3953 1669 4016
rect 1698 4013 1701 4026
rect 1746 3993 1749 4006
rect 1658 3886 1661 3926
rect 1666 3913 1669 3926
rect 1626 3873 1637 3876
rect 1650 3883 1661 3886
rect 1578 3793 1581 3806
rect 1586 3803 1597 3806
rect 1610 3803 1613 3816
rect 1618 3813 1621 3826
rect 1594 3746 1597 3786
rect 1618 3783 1621 3806
rect 1626 3803 1629 3873
rect 1650 3816 1653 3883
rect 1634 3796 1637 3816
rect 1642 3803 1645 3816
rect 1650 3813 1661 3816
rect 1682 3813 1685 3826
rect 1690 3813 1701 3816
rect 1650 3796 1653 3806
rect 1634 3793 1653 3796
rect 1658 3786 1661 3813
rect 1706 3806 1709 3956
rect 1762 3953 1765 4016
rect 1834 4013 1837 4053
rect 1858 4013 1861 4140
rect 1770 3976 1773 3996
rect 1858 3993 1861 4006
rect 1874 3976 1877 4140
rect 1770 3973 1781 3976
rect 1722 3913 1725 3926
rect 1722 3813 1725 3826
rect 1642 3783 1661 3786
rect 1698 3803 1709 3806
rect 1586 3743 1597 3746
rect 1586 3686 1589 3743
rect 1618 3733 1621 3746
rect 1642 3736 1645 3783
rect 1698 3746 1701 3803
rect 1690 3743 1701 3746
rect 1642 3733 1649 3736
rect 1634 3696 1637 3726
rect 1626 3693 1637 3696
rect 1522 3673 1533 3676
rect 1522 3603 1525 3673
rect 1530 3613 1541 3616
rect 1546 3613 1549 3686
rect 1586 3683 1613 3686
rect 1538 3593 1541 3606
rect 1554 3603 1557 3636
rect 1562 3603 1565 3626
rect 1570 3596 1573 3616
rect 1578 3613 1589 3616
rect 1562 3593 1573 3596
rect 1514 3573 1525 3576
rect 1490 3476 1493 3506
rect 1498 3483 1501 3536
rect 1490 3473 1501 3476
rect 1482 3413 1485 3426
rect 1442 3293 1449 3296
rect 1458 3333 1469 3336
rect 1442 3246 1445 3293
rect 1458 3256 1461 3333
rect 1466 3313 1469 3326
rect 1490 3283 1493 3466
rect 1498 3413 1501 3473
rect 1506 3463 1509 3526
rect 1514 3473 1517 3536
rect 1522 3513 1525 3573
rect 1498 3396 1501 3406
rect 1506 3403 1509 3416
rect 1514 3396 1517 3416
rect 1498 3393 1517 3396
rect 1522 3393 1525 3406
rect 1530 3376 1533 3556
rect 1546 3533 1549 3556
rect 1554 3523 1557 3536
rect 1562 3523 1565 3593
rect 1578 3583 1581 3606
rect 1586 3566 1589 3613
rect 1594 3603 1597 3616
rect 1602 3613 1605 3666
rect 1610 3586 1613 3683
rect 1618 3596 1621 3616
rect 1626 3603 1629 3693
rect 1646 3686 1649 3733
rect 1674 3686 1677 3726
rect 1690 3696 1693 3743
rect 1690 3693 1701 3696
rect 1642 3683 1649 3686
rect 1658 3683 1677 3686
rect 1634 3596 1637 3606
rect 1618 3593 1637 3596
rect 1610 3583 1621 3586
rect 1578 3563 1589 3566
rect 1570 3533 1573 3546
rect 1506 3373 1533 3376
rect 1458 3253 1469 3256
rect 1434 3243 1445 3246
rect 1418 3213 1421 3226
rect 1434 3196 1437 3243
rect 1434 3193 1445 3196
rect 1418 3113 1421 3126
rect 1434 3103 1437 3166
rect 1402 3013 1413 3016
rect 1418 2936 1421 3066
rect 1434 3013 1437 3026
rect 1386 2913 1397 2916
rect 1386 2896 1389 2913
rect 1322 2803 1325 2816
rect 1322 2766 1325 2796
rect 1314 2763 1325 2766
rect 1330 2763 1333 2816
rect 1346 2813 1365 2816
rect 1378 2893 1389 2896
rect 1314 2746 1317 2763
rect 1338 2753 1341 2806
rect 1346 2796 1349 2813
rect 1378 2806 1381 2893
rect 1402 2886 1405 2936
rect 1418 2933 1433 2936
rect 1418 2913 1421 2926
rect 1394 2883 1405 2886
rect 1394 2813 1397 2883
rect 1378 2803 1389 2806
rect 1346 2793 1365 2796
rect 1314 2743 1341 2746
rect 1338 2736 1341 2743
rect 1274 2703 1281 2706
rect 1278 2546 1281 2703
rect 1302 2703 1309 2706
rect 1290 2613 1293 2656
rect 1302 2616 1305 2703
rect 1314 2653 1317 2736
rect 1302 2613 1309 2616
rect 1322 2613 1325 2726
rect 1330 2723 1333 2736
rect 1338 2733 1357 2736
rect 1362 2733 1365 2793
rect 1338 2723 1349 2726
rect 1370 2723 1373 2776
rect 1274 2543 1281 2546
rect 1274 2513 1277 2543
rect 1306 2533 1309 2613
rect 1330 2606 1333 2706
rect 1330 2603 1341 2606
rect 1258 2493 1269 2496
rect 1258 2343 1261 2426
rect 1266 2413 1269 2493
rect 1282 2423 1285 2526
rect 1282 2406 1285 2416
rect 1266 2403 1285 2406
rect 1290 2403 1293 2496
rect 1306 2493 1309 2526
rect 1314 2476 1317 2576
rect 1310 2473 1317 2476
rect 1298 2403 1301 2466
rect 1266 2283 1269 2336
rect 1290 2296 1293 2346
rect 1298 2313 1301 2326
rect 1290 2293 1297 2296
rect 1250 2193 1253 2206
rect 1274 2196 1277 2216
rect 1266 2193 1277 2196
rect 1242 2123 1245 2136
rect 1234 2103 1241 2106
rect 1238 1996 1241 2103
rect 1250 2096 1253 2186
rect 1266 2133 1269 2193
rect 1282 2186 1285 2286
rect 1274 2183 1285 2186
rect 1258 2113 1261 2126
rect 1274 2123 1277 2183
rect 1294 2176 1297 2293
rect 1310 2266 1313 2473
rect 1310 2263 1317 2266
rect 1290 2173 1297 2176
rect 1250 2093 1261 2096
rect 1290 2093 1293 2173
rect 1258 2036 1261 2093
rect 1234 1993 1241 1996
rect 1250 2033 1261 2036
rect 1234 1926 1237 1993
rect 1234 1923 1241 1926
rect 1226 1803 1229 1916
rect 1238 1826 1241 1923
rect 1234 1823 1241 1826
rect 1234 1803 1237 1823
rect 1226 1726 1229 1796
rect 1234 1733 1237 1756
rect 1242 1733 1245 1806
rect 1226 1723 1237 1726
rect 1218 1713 1229 1716
rect 1234 1713 1237 1723
rect 1218 1456 1221 1626
rect 1202 1453 1221 1456
rect 1202 1363 1205 1453
rect 1210 1393 1213 1416
rect 1146 1163 1157 1166
rect 1162 1223 1173 1226
rect 1162 1166 1165 1223
rect 1186 1213 1189 1266
rect 1170 1183 1173 1206
rect 1162 1163 1169 1166
rect 1146 1076 1149 1163
rect 1166 1086 1169 1163
rect 1178 1133 1181 1206
rect 1194 1203 1197 1216
rect 1202 1213 1205 1226
rect 1186 1133 1189 1146
rect 1162 1083 1169 1086
rect 1146 1073 1153 1076
rect 1150 936 1153 1073
rect 1162 986 1165 1083
rect 1178 1036 1181 1126
rect 1170 1033 1181 1036
rect 1170 1003 1173 1033
rect 1186 1006 1189 1116
rect 1178 1003 1189 1006
rect 1162 983 1173 986
rect 1146 933 1153 936
rect 1146 913 1149 933
rect 1170 916 1173 983
rect 1194 963 1197 1126
rect 1202 1123 1205 1206
rect 1210 1203 1213 1326
rect 1218 1193 1221 1366
rect 1226 1243 1229 1713
rect 1242 1693 1245 1716
rect 1234 1286 1237 1626
rect 1242 1413 1245 1536
rect 1250 1363 1253 2033
rect 1290 2016 1293 2026
rect 1274 2013 1293 2016
rect 1306 2013 1309 2116
rect 1314 2083 1317 2263
rect 1314 2013 1317 2026
rect 1322 2013 1325 2536
rect 1330 2516 1333 2603
rect 1338 2533 1341 2556
rect 1330 2513 1337 2516
rect 1334 2446 1337 2513
rect 1330 2443 1337 2446
rect 1330 2413 1333 2443
rect 1274 2003 1277 2013
rect 1258 1923 1261 1966
rect 1266 1913 1269 1986
rect 1282 1933 1285 2006
rect 1298 2003 1309 2006
rect 1306 1933 1309 1946
rect 1258 1813 1261 1846
rect 1258 1743 1261 1806
rect 1258 1713 1261 1726
rect 1266 1693 1269 1736
rect 1274 1656 1277 1926
rect 1282 1923 1301 1926
rect 1314 1843 1317 1966
rect 1330 1933 1333 2406
rect 1338 2203 1341 2426
rect 1346 2386 1349 2706
rect 1378 2636 1381 2756
rect 1386 2703 1389 2803
rect 1394 2713 1397 2736
rect 1370 2633 1381 2636
rect 1370 2553 1373 2633
rect 1354 2456 1357 2536
rect 1362 2493 1365 2546
rect 1386 2526 1389 2616
rect 1402 2583 1405 2736
rect 1410 2733 1413 2766
rect 1418 2676 1421 2846
rect 1430 2836 1433 2933
rect 1442 2873 1445 3193
rect 1466 3163 1469 3253
rect 1482 3203 1485 3256
rect 1450 2976 1453 3046
rect 1458 2983 1461 3086
rect 1466 3043 1469 3156
rect 1450 2973 1469 2976
rect 1466 2836 1469 2973
rect 1482 2946 1485 3106
rect 1490 3063 1493 3266
rect 1498 3206 1501 3326
rect 1506 3306 1509 3373
rect 1538 3336 1541 3416
rect 1530 3333 1541 3336
rect 1530 3313 1533 3326
rect 1506 3303 1517 3306
rect 1514 3236 1517 3303
rect 1506 3233 1517 3236
rect 1506 3216 1509 3233
rect 1506 3213 1525 3216
rect 1530 3213 1533 3286
rect 1546 3263 1549 3426
rect 1554 3353 1557 3406
rect 1570 3403 1573 3436
rect 1554 3343 1573 3346
rect 1554 3333 1557 3343
rect 1562 3303 1565 3336
rect 1570 3323 1573 3343
rect 1498 3203 1517 3206
rect 1514 3013 1517 3126
rect 1522 3083 1525 3213
rect 1538 3203 1541 3216
rect 1546 3213 1549 3236
rect 1578 3233 1581 3563
rect 1594 3523 1597 3566
rect 1610 3533 1613 3546
rect 1618 3526 1621 3583
rect 1602 3523 1621 3526
rect 1626 3523 1629 3536
rect 1634 3533 1637 3546
rect 1594 3413 1597 3426
rect 1602 3406 1605 3523
rect 1642 3516 1645 3683
rect 1658 3613 1661 3683
rect 1698 3646 1701 3693
rect 1694 3643 1701 3646
rect 1650 3523 1653 3546
rect 1658 3533 1661 3606
rect 1674 3566 1677 3616
rect 1682 3613 1685 3626
rect 1694 3576 1697 3643
rect 1722 3596 1725 3746
rect 1738 3723 1741 3796
rect 1746 3786 1749 3946
rect 1762 3913 1765 3926
rect 1778 3906 1781 3973
rect 1802 3943 1821 3946
rect 1802 3933 1805 3943
rect 1770 3903 1781 3906
rect 1746 3783 1753 3786
rect 1750 3716 1753 3783
rect 1770 3743 1773 3903
rect 1786 3793 1789 3806
rect 1746 3713 1753 3716
rect 1746 3643 1749 3713
rect 1778 3653 1781 3756
rect 1794 3736 1797 3926
rect 1810 3923 1813 3936
rect 1818 3923 1821 3943
rect 1826 3886 1829 3936
rect 1834 3903 1837 3966
rect 1850 3946 1853 3976
rect 1870 3973 1877 3976
rect 1882 3973 1885 4016
rect 1850 3943 1861 3946
rect 1818 3883 1829 3886
rect 1810 3763 1813 3816
rect 1818 3783 1821 3883
rect 1826 3813 1829 3836
rect 1834 3813 1837 3826
rect 1842 3803 1845 3936
rect 1858 3846 1861 3943
rect 1850 3843 1861 3846
rect 1786 3733 1797 3736
rect 1738 3603 1741 3616
rect 1762 3603 1765 3646
rect 1778 3603 1781 3626
rect 1722 3593 1733 3596
rect 1694 3573 1701 3576
rect 1674 3563 1685 3566
rect 1682 3523 1685 3563
rect 1642 3513 1653 3516
rect 1610 3413 1613 3496
rect 1586 3393 1589 3406
rect 1594 3403 1613 3406
rect 1586 3323 1589 3336
rect 1594 3323 1597 3356
rect 1602 3333 1605 3403
rect 1618 3383 1621 3416
rect 1634 3413 1637 3426
rect 1650 3413 1653 3513
rect 1698 3426 1701 3573
rect 1730 3503 1733 3593
rect 1746 3523 1749 3536
rect 1754 3523 1757 3576
rect 1786 3573 1789 3733
rect 1794 3713 1797 3726
rect 1794 3566 1797 3656
rect 1810 3636 1813 3666
rect 1818 3643 1821 3736
rect 1834 3733 1837 3766
rect 1850 3753 1853 3843
rect 1870 3826 1873 3973
rect 1858 3823 1873 3826
rect 1858 3736 1861 3823
rect 1866 3796 1869 3816
rect 1874 3803 1877 3816
rect 1882 3813 1885 3886
rect 1882 3796 1885 3806
rect 1866 3793 1885 3796
rect 1850 3733 1861 3736
rect 1834 3713 1837 3726
rect 1850 3706 1853 3733
rect 1834 3703 1853 3706
rect 1810 3633 1821 3636
rect 1802 3613 1805 3626
rect 1818 3613 1821 3633
rect 1786 3563 1797 3566
rect 1778 3533 1781 3546
rect 1770 3513 1773 3526
rect 1650 3393 1653 3406
rect 1658 3403 1661 3426
rect 1682 3413 1685 3426
rect 1698 3423 1709 3426
rect 1690 3413 1701 3416
rect 1698 3393 1701 3413
rect 1706 3386 1709 3423
rect 1722 3413 1725 3426
rect 1746 3406 1749 3426
rect 1690 3383 1709 3386
rect 1738 3403 1749 3406
rect 1666 3346 1669 3366
rect 1666 3343 1673 3346
rect 1554 3113 1557 3216
rect 1562 3203 1565 3216
rect 1594 3213 1597 3246
rect 1570 3203 1581 3206
rect 1586 3193 1589 3206
rect 1610 3196 1613 3216
rect 1602 3193 1613 3196
rect 1602 3183 1605 3193
rect 1610 3183 1621 3186
rect 1578 3133 1589 3136
rect 1522 3006 1525 3076
rect 1530 3013 1533 3036
rect 1498 3003 1509 3006
rect 1522 3003 1533 3006
rect 1482 2943 1493 2946
rect 1482 2903 1485 2936
rect 1490 2843 1493 2943
rect 1498 2873 1501 2986
rect 1506 2933 1509 2996
rect 1506 2903 1509 2926
rect 1514 2846 1517 2976
rect 1522 2923 1525 2936
rect 1530 2883 1533 3003
rect 1538 2983 1541 3006
rect 1546 3003 1549 3016
rect 1562 3013 1565 3026
rect 1554 2976 1557 3006
rect 1570 3003 1573 3126
rect 1578 3113 1581 3126
rect 1538 2973 1557 2976
rect 1538 2933 1541 2973
rect 1546 2933 1549 2946
rect 1506 2843 1517 2846
rect 1430 2833 1437 2836
rect 1426 2723 1429 2816
rect 1434 2776 1437 2833
rect 1458 2833 1469 2836
rect 1434 2773 1445 2776
rect 1434 2693 1437 2766
rect 1410 2673 1421 2676
rect 1442 2676 1445 2773
rect 1458 2753 1461 2833
rect 1450 2683 1453 2736
rect 1466 2703 1469 2736
rect 1490 2723 1493 2816
rect 1498 2793 1501 2816
rect 1442 2673 1469 2676
rect 1410 2556 1413 2673
rect 1418 2593 1421 2666
rect 1434 2616 1437 2646
rect 1426 2613 1453 2616
rect 1442 2593 1445 2606
rect 1370 2523 1389 2526
rect 1394 2553 1413 2556
rect 1354 2453 1365 2456
rect 1354 2403 1357 2416
rect 1346 2383 1353 2386
rect 1350 2306 1353 2383
rect 1362 2343 1365 2453
rect 1370 2353 1373 2523
rect 1394 2516 1397 2553
rect 1418 2546 1421 2566
rect 1402 2533 1405 2546
rect 1418 2543 1425 2546
rect 1386 2513 1397 2516
rect 1386 2436 1389 2513
rect 1410 2506 1413 2526
rect 1378 2433 1389 2436
rect 1402 2503 1413 2506
rect 1378 2403 1381 2433
rect 1346 2303 1353 2306
rect 1346 2196 1349 2303
rect 1354 2213 1357 2286
rect 1362 2213 1365 2336
rect 1386 2326 1389 2416
rect 1402 2403 1405 2503
rect 1410 2413 1413 2496
rect 1422 2426 1425 2543
rect 1434 2463 1437 2586
rect 1466 2573 1469 2673
rect 1474 2613 1477 2646
rect 1482 2596 1485 2686
rect 1490 2603 1493 2706
rect 1498 2613 1501 2786
rect 1506 2776 1509 2843
rect 1538 2826 1541 2926
rect 1546 2903 1549 2926
rect 1514 2823 1541 2826
rect 1514 2813 1517 2823
rect 1514 2796 1517 2806
rect 1522 2803 1525 2816
rect 1530 2796 1533 2816
rect 1546 2813 1549 2846
rect 1554 2813 1557 2956
rect 1562 2893 1565 2936
rect 1570 2933 1573 2996
rect 1578 2933 1581 3016
rect 1586 3013 1589 3066
rect 1594 3053 1597 3136
rect 1618 3133 1621 3156
rect 1602 3073 1605 3126
rect 1618 3093 1621 3126
rect 1602 3053 1613 3056
rect 1586 2936 1589 3006
rect 1594 3003 1597 3046
rect 1602 3033 1605 3053
rect 1626 3043 1629 3336
rect 1634 3213 1653 3216
rect 1642 3183 1645 3206
rect 1650 3203 1653 3213
rect 1634 3123 1637 3146
rect 1642 3133 1645 3156
rect 1650 3133 1653 3146
rect 1658 3126 1661 3266
rect 1670 3246 1673 3343
rect 1682 3313 1685 3326
rect 1690 3296 1693 3383
rect 1738 3346 1741 3403
rect 1770 3366 1773 3506
rect 1786 3423 1789 3563
rect 1810 3536 1813 3606
rect 1826 3603 1829 3616
rect 1794 3513 1797 3536
rect 1802 3533 1813 3536
rect 1754 3363 1773 3366
rect 1738 3343 1749 3346
rect 1714 3303 1717 3336
rect 1730 3313 1733 3326
rect 1690 3293 1701 3296
rect 1746 3293 1749 3343
rect 1754 3316 1757 3363
rect 1762 3323 1765 3336
rect 1770 3333 1773 3356
rect 1786 3343 1789 3416
rect 1802 3406 1805 3533
rect 1810 3513 1813 3526
rect 1818 3523 1829 3526
rect 1794 3403 1805 3406
rect 1754 3313 1765 3316
rect 1770 3313 1773 3326
rect 1778 3323 1789 3326
rect 1698 3256 1701 3293
rect 1666 3243 1673 3246
rect 1694 3253 1701 3256
rect 1666 3196 1669 3243
rect 1674 3213 1677 3226
rect 1666 3193 1673 3196
rect 1650 3123 1661 3126
rect 1650 3033 1653 3123
rect 1670 3116 1673 3193
rect 1682 3183 1685 3216
rect 1694 3176 1697 3253
rect 1714 3213 1717 3226
rect 1738 3196 1741 3236
rect 1738 3193 1749 3196
rect 1694 3173 1701 3176
rect 1666 3113 1673 3116
rect 1682 3113 1685 3126
rect 1690 3123 1693 3156
rect 1666 3056 1669 3113
rect 1698 3106 1701 3173
rect 1746 3146 1749 3193
rect 1762 3176 1765 3313
rect 1778 3193 1781 3286
rect 1762 3173 1773 3176
rect 1738 3143 1749 3146
rect 1722 3113 1725 3126
rect 1658 3053 1669 3056
rect 1682 3103 1701 3106
rect 1618 3016 1621 3026
rect 1602 2996 1605 3016
rect 1610 3003 1613 3016
rect 1618 3013 1629 3016
rect 1634 3013 1637 3026
rect 1642 3013 1653 3016
rect 1618 2996 1621 3006
rect 1602 2993 1621 2996
rect 1602 2943 1621 2946
rect 1586 2933 1597 2936
rect 1562 2813 1565 2856
rect 1570 2836 1573 2926
rect 1578 2893 1581 2926
rect 1586 2913 1589 2926
rect 1594 2916 1597 2933
rect 1602 2923 1605 2943
rect 1594 2913 1605 2916
rect 1570 2833 1581 2836
rect 1578 2813 1581 2833
rect 1514 2793 1533 2796
rect 1506 2773 1513 2776
rect 1510 2706 1513 2773
rect 1538 2726 1541 2806
rect 1562 2803 1573 2806
rect 1586 2803 1589 2826
rect 1594 2813 1597 2866
rect 1506 2703 1513 2706
rect 1530 2723 1549 2726
rect 1554 2723 1557 2756
rect 1570 2723 1573 2776
rect 1506 2683 1509 2703
rect 1506 2613 1509 2676
rect 1514 2603 1517 2636
rect 1522 2613 1525 2646
rect 1530 2603 1533 2723
rect 1578 2706 1581 2736
rect 1586 2723 1589 2796
rect 1574 2703 1581 2706
rect 1574 2636 1577 2703
rect 1594 2686 1597 2806
rect 1602 2753 1605 2913
rect 1610 2823 1613 2936
rect 1618 2933 1621 2943
rect 1610 2766 1613 2816
rect 1626 2813 1629 3013
rect 1634 2913 1637 2926
rect 1642 2923 1653 2926
rect 1658 2866 1661 3053
rect 1674 3013 1677 3026
rect 1674 2913 1677 2926
rect 1682 2896 1685 3103
rect 1738 3096 1741 3143
rect 1690 3076 1693 3096
rect 1738 3093 1749 3096
rect 1690 3073 1697 3076
rect 1694 2896 1697 3073
rect 1650 2863 1661 2866
rect 1678 2893 1685 2896
rect 1690 2893 1697 2896
rect 1634 2816 1637 2836
rect 1634 2813 1645 2816
rect 1650 2813 1653 2863
rect 1658 2813 1661 2856
rect 1618 2793 1621 2806
rect 1610 2763 1629 2766
rect 1626 2753 1629 2763
rect 1634 2736 1637 2813
rect 1626 2733 1637 2736
rect 1574 2633 1581 2636
rect 1482 2593 1493 2596
rect 1442 2523 1445 2536
rect 1450 2513 1453 2526
rect 1418 2423 1425 2426
rect 1418 2333 1421 2423
rect 1426 2373 1429 2406
rect 1442 2386 1445 2406
rect 1442 2383 1449 2386
rect 1370 2306 1373 2326
rect 1378 2323 1389 2326
rect 1370 2303 1377 2306
rect 1374 2226 1377 2303
rect 1426 2246 1429 2346
rect 1434 2333 1437 2356
rect 1446 2316 1449 2383
rect 1458 2323 1461 2346
rect 1466 2323 1469 2566
rect 1474 2533 1485 2536
rect 1490 2533 1493 2593
rect 1546 2526 1549 2606
rect 1474 2413 1477 2456
rect 1506 2383 1509 2466
rect 1506 2356 1509 2376
rect 1498 2353 1509 2356
rect 1442 2313 1449 2316
rect 1442 2293 1445 2313
rect 1482 2276 1485 2326
rect 1498 2296 1501 2353
rect 1514 2343 1517 2526
rect 1546 2523 1557 2526
rect 1522 2366 1525 2456
rect 1530 2413 1533 2426
rect 1554 2403 1557 2523
rect 1562 2513 1565 2526
rect 1570 2523 1573 2616
rect 1578 2613 1581 2633
rect 1578 2463 1581 2526
rect 1586 2523 1589 2686
rect 1594 2683 1613 2686
rect 1610 2666 1613 2683
rect 1626 2676 1629 2733
rect 1634 2713 1637 2726
rect 1642 2686 1645 2796
rect 1650 2743 1653 2806
rect 1666 2783 1669 2836
rect 1678 2826 1681 2893
rect 1678 2823 1685 2826
rect 1674 2766 1677 2806
rect 1682 2793 1685 2823
rect 1690 2783 1693 2893
rect 1674 2763 1693 2766
rect 1666 2703 1669 2746
rect 1682 2733 1685 2756
rect 1682 2713 1685 2726
rect 1642 2683 1649 2686
rect 1626 2673 1637 2676
rect 1610 2663 1617 2666
rect 1594 2593 1597 2616
rect 1614 2596 1617 2663
rect 1610 2593 1617 2596
rect 1610 2576 1613 2593
rect 1606 2573 1613 2576
rect 1570 2413 1573 2426
rect 1586 2403 1589 2426
rect 1594 2403 1597 2546
rect 1606 2436 1609 2573
rect 1626 2533 1629 2616
rect 1634 2613 1637 2673
rect 1646 2606 1649 2683
rect 1690 2643 1693 2763
rect 1698 2713 1701 2876
rect 1714 2766 1717 2886
rect 1710 2763 1717 2766
rect 1642 2603 1649 2606
rect 1618 2513 1621 2526
rect 1602 2433 1609 2436
rect 1522 2363 1533 2366
rect 1498 2293 1509 2296
rect 1482 2273 1497 2276
rect 1370 2223 1377 2226
rect 1418 2243 1429 2246
rect 1370 2206 1373 2223
rect 1338 2193 1349 2196
rect 1354 2203 1373 2206
rect 1338 2106 1341 2193
rect 1354 2123 1357 2203
rect 1362 2133 1365 2196
rect 1402 2193 1405 2216
rect 1362 2106 1365 2126
rect 1338 2103 1349 2106
rect 1346 2026 1349 2103
rect 1342 2023 1349 2026
rect 1358 2103 1365 2106
rect 1358 2026 1361 2103
rect 1370 2026 1373 2126
rect 1386 2036 1389 2136
rect 1410 2123 1413 2186
rect 1418 2106 1421 2243
rect 1414 2103 1421 2106
rect 1414 2036 1417 2103
rect 1426 2046 1429 2166
rect 1442 2156 1445 2206
rect 1466 2166 1469 2206
rect 1494 2186 1497 2273
rect 1494 2183 1501 2186
rect 1466 2163 1493 2166
rect 1442 2153 1453 2156
rect 1450 2106 1453 2153
rect 1466 2113 1469 2126
rect 1450 2103 1461 2106
rect 1426 2043 1433 2046
rect 1386 2033 1393 2036
rect 1414 2033 1421 2036
rect 1358 2023 1365 2026
rect 1370 2023 1381 2026
rect 1342 1956 1345 2023
rect 1338 1953 1345 1956
rect 1282 1716 1285 1756
rect 1290 1726 1293 1736
rect 1298 1733 1301 1746
rect 1314 1733 1317 1816
rect 1322 1793 1325 1926
rect 1338 1773 1341 1953
rect 1346 1866 1349 1936
rect 1354 1873 1357 2006
rect 1362 1926 1365 2023
rect 1378 1966 1381 2023
rect 1390 1986 1393 2033
rect 1410 2003 1413 2016
rect 1370 1963 1381 1966
rect 1386 1983 1393 1986
rect 1386 1963 1389 1983
rect 1370 1933 1373 1946
rect 1362 1923 1373 1926
rect 1378 1923 1381 1963
rect 1386 1933 1413 1936
rect 1370 1916 1373 1923
rect 1386 1916 1389 1926
rect 1370 1913 1389 1916
rect 1346 1863 1365 1866
rect 1330 1733 1341 1736
rect 1290 1723 1309 1726
rect 1282 1713 1297 1716
rect 1306 1713 1309 1723
rect 1274 1653 1285 1656
rect 1274 1613 1277 1646
rect 1282 1606 1285 1653
rect 1294 1636 1297 1713
rect 1294 1633 1301 1636
rect 1298 1613 1301 1633
rect 1266 1573 1269 1606
rect 1274 1603 1285 1606
rect 1258 1483 1261 1526
rect 1274 1476 1277 1603
rect 1290 1593 1293 1606
rect 1258 1473 1277 1476
rect 1258 1333 1261 1473
rect 1282 1413 1285 1486
rect 1234 1283 1253 1286
rect 1210 1113 1213 1136
rect 1218 1123 1221 1186
rect 1202 1013 1205 1066
rect 1226 1026 1229 1206
rect 1234 1203 1237 1216
rect 1242 1213 1245 1226
rect 1250 1206 1253 1283
rect 1242 1203 1253 1206
rect 1242 1033 1245 1203
rect 1258 1113 1261 1236
rect 1274 1203 1277 1406
rect 1290 1393 1293 1406
rect 1298 1233 1301 1556
rect 1306 1416 1309 1696
rect 1314 1553 1317 1676
rect 1314 1523 1317 1536
rect 1306 1413 1317 1416
rect 1322 1413 1325 1726
rect 1330 1713 1333 1726
rect 1330 1596 1333 1636
rect 1338 1603 1341 1733
rect 1346 1693 1349 1746
rect 1354 1733 1357 1816
rect 1362 1736 1365 1863
rect 1370 1813 1381 1816
rect 1378 1803 1381 1813
rect 1362 1733 1373 1736
rect 1378 1723 1381 1756
rect 1386 1733 1389 1806
rect 1394 1743 1397 1846
rect 1354 1603 1357 1616
rect 1330 1593 1341 1596
rect 1378 1593 1381 1616
rect 1394 1593 1397 1666
rect 1338 1576 1341 1593
rect 1338 1573 1345 1576
rect 1342 1486 1345 1573
rect 1338 1483 1345 1486
rect 1338 1426 1341 1483
rect 1334 1423 1341 1426
rect 1354 1426 1357 1566
rect 1402 1563 1405 1876
rect 1410 1843 1413 1933
rect 1418 1856 1421 2033
rect 1430 1976 1433 2043
rect 1458 1976 1461 2103
rect 1426 1973 1433 1976
rect 1450 1973 1461 1976
rect 1474 1973 1477 2016
rect 1426 1873 1429 1973
rect 1442 1923 1445 1946
rect 1450 1856 1453 1973
rect 1482 1966 1485 2056
rect 1490 1983 1493 2163
rect 1498 2156 1501 2183
rect 1506 2163 1509 2293
rect 1514 2213 1517 2326
rect 1522 2273 1525 2356
rect 1530 2166 1533 2363
rect 1538 2306 1541 2386
rect 1538 2303 1545 2306
rect 1526 2163 1533 2166
rect 1498 2153 1517 2156
rect 1506 2113 1509 2126
rect 1514 2106 1517 2153
rect 1498 2103 1517 2106
rect 1498 1976 1501 2103
rect 1526 2056 1529 2163
rect 1542 2156 1545 2303
rect 1554 2196 1557 2346
rect 1562 2343 1581 2346
rect 1562 2333 1565 2343
rect 1570 2203 1573 2336
rect 1578 2323 1581 2343
rect 1586 2226 1589 2336
rect 1602 2323 1605 2433
rect 1618 2413 1621 2426
rect 1626 2403 1629 2456
rect 1634 2413 1637 2526
rect 1642 2383 1645 2603
rect 1658 2593 1661 2606
rect 1650 2566 1653 2586
rect 1674 2583 1677 2606
rect 1650 2563 1661 2566
rect 1658 2436 1661 2563
rect 1650 2433 1661 2436
rect 1634 2333 1637 2346
rect 1650 2343 1653 2433
rect 1578 2223 1589 2226
rect 1554 2193 1573 2196
rect 1538 2153 1545 2156
rect 1526 2053 1533 2056
rect 1538 2053 1541 2153
rect 1554 2133 1557 2166
rect 1530 2033 1533 2053
rect 1498 1973 1509 1976
rect 1458 1893 1461 1966
rect 1466 1963 1485 1966
rect 1466 1876 1469 1963
rect 1490 1923 1493 1936
rect 1418 1853 1429 1856
rect 1410 1803 1413 1816
rect 1410 1693 1413 1796
rect 1426 1766 1429 1853
rect 1418 1763 1429 1766
rect 1442 1853 1453 1856
rect 1462 1873 1469 1876
rect 1418 1656 1421 1763
rect 1426 1706 1429 1736
rect 1442 1733 1445 1853
rect 1462 1766 1465 1873
rect 1462 1763 1469 1766
rect 1466 1743 1469 1763
rect 1466 1723 1469 1736
rect 1426 1703 1437 1706
rect 1418 1653 1425 1656
rect 1422 1576 1425 1653
rect 1434 1613 1437 1703
rect 1418 1573 1425 1576
rect 1370 1503 1373 1526
rect 1378 1483 1381 1536
rect 1402 1533 1413 1536
rect 1402 1503 1405 1526
rect 1418 1486 1421 1573
rect 1410 1483 1421 1486
rect 1354 1423 1361 1426
rect 1306 1373 1309 1406
rect 1314 1383 1317 1413
rect 1334 1356 1337 1423
rect 1334 1353 1341 1356
rect 1314 1313 1317 1336
rect 1322 1333 1333 1336
rect 1282 1213 1301 1216
rect 1314 1213 1317 1226
rect 1330 1223 1333 1326
rect 1338 1316 1341 1353
rect 1346 1323 1349 1416
rect 1338 1313 1345 1316
rect 1282 1183 1285 1213
rect 1226 1023 1245 1026
rect 1218 963 1221 1006
rect 1162 913 1173 916
rect 1194 913 1197 936
rect 1162 883 1165 913
rect 1202 906 1205 936
rect 1210 923 1213 936
rect 1218 933 1229 936
rect 1234 933 1237 1016
rect 1242 1006 1245 1023
rect 1242 1003 1249 1006
rect 1246 946 1249 1003
rect 1242 943 1249 946
rect 1194 903 1205 906
rect 1154 813 1157 826
rect 1178 756 1181 896
rect 1170 753 1181 756
rect 1130 723 1133 746
rect 1138 723 1141 736
rect 1146 723 1149 736
rect 1154 666 1157 736
rect 1146 663 1157 666
rect 1102 593 1109 596
rect 1106 576 1109 593
rect 1106 573 1117 576
rect 1042 503 1045 523
rect 1066 513 1069 536
rect 1074 526 1077 536
rect 1074 523 1085 526
rect 1090 523 1093 536
rect 1002 443 1013 446
rect 986 363 989 406
rect 994 403 997 416
rect 1010 413 1013 443
rect 1010 393 1013 406
rect 1034 403 1037 416
rect 978 353 989 356
rect 970 333 973 346
rect 978 323 981 346
rect 986 333 989 353
rect 994 323 997 336
rect 970 296 973 316
rect 970 293 981 296
rect 978 236 981 293
rect 994 256 997 296
rect 1002 263 1005 356
rect 1010 266 1013 336
rect 1018 323 1021 366
rect 1034 333 1037 346
rect 1034 286 1037 326
rect 1026 283 1037 286
rect 1010 263 1021 266
rect 994 253 1013 256
rect 954 213 957 236
rect 970 233 981 236
rect 970 213 973 233
rect 922 193 941 196
rect 954 123 957 206
rect 994 193 997 206
rect 978 133 981 146
rect 1002 123 1005 216
rect 1010 213 1013 253
rect 1018 203 1021 263
rect 1026 233 1029 283
rect 1042 236 1045 336
rect 1050 326 1053 466
rect 1074 456 1077 516
rect 1082 483 1085 523
rect 1098 473 1101 536
rect 1106 523 1109 536
rect 1106 503 1109 516
rect 1114 496 1117 573
rect 1106 493 1117 496
rect 1074 453 1081 456
rect 1078 386 1081 453
rect 1074 383 1081 386
rect 1074 363 1077 383
rect 1058 333 1069 336
rect 1074 333 1077 346
rect 1090 343 1093 416
rect 1106 403 1109 493
rect 1122 443 1125 636
rect 1146 613 1149 663
rect 1130 503 1133 536
rect 1138 523 1141 596
rect 1170 576 1173 753
rect 1186 746 1189 776
rect 1178 743 1189 746
rect 1194 736 1197 903
rect 1226 886 1229 926
rect 1234 913 1237 926
rect 1242 896 1245 943
rect 1218 883 1229 886
rect 1238 893 1245 896
rect 1202 743 1205 816
rect 1210 803 1213 826
rect 1218 736 1221 883
rect 1226 803 1229 856
rect 1238 826 1241 893
rect 1238 823 1245 826
rect 1234 783 1237 806
rect 1242 776 1245 823
rect 1250 813 1253 926
rect 1258 813 1261 1006
rect 1266 1003 1269 1056
rect 1274 976 1277 1016
rect 1266 973 1277 976
rect 1266 853 1269 973
rect 1282 966 1285 1166
rect 1290 1116 1293 1136
rect 1306 1123 1309 1206
rect 1322 1163 1325 1206
rect 1330 1203 1333 1216
rect 1342 1166 1345 1313
rect 1358 1306 1361 1423
rect 1370 1413 1373 1426
rect 1378 1393 1381 1406
rect 1386 1403 1389 1416
rect 1410 1376 1413 1483
rect 1426 1413 1429 1526
rect 1434 1513 1437 1536
rect 1450 1503 1453 1606
rect 1426 1383 1429 1406
rect 1410 1373 1421 1376
rect 1354 1303 1361 1306
rect 1342 1163 1349 1166
rect 1330 1133 1333 1156
rect 1290 1113 1297 1116
rect 1294 966 1297 1113
rect 1274 963 1285 966
rect 1290 963 1297 966
rect 1274 886 1277 963
rect 1290 943 1293 963
rect 1290 923 1293 936
rect 1274 883 1285 886
rect 1178 723 1181 736
rect 1186 733 1197 736
rect 1186 723 1189 733
rect 1194 613 1197 726
rect 1202 706 1205 736
rect 1210 733 1221 736
rect 1226 773 1245 776
rect 1226 733 1229 773
rect 1258 746 1261 806
rect 1266 793 1269 816
rect 1274 813 1277 826
rect 1282 803 1285 883
rect 1298 803 1301 816
rect 1306 776 1309 1116
rect 1346 1076 1349 1163
rect 1338 1073 1349 1076
rect 1314 1013 1317 1066
rect 1338 1006 1341 1073
rect 1354 1053 1357 1303
rect 1370 1276 1373 1336
rect 1386 1333 1389 1366
rect 1410 1323 1413 1336
rect 1370 1273 1381 1276
rect 1378 1226 1381 1273
rect 1370 1223 1381 1226
rect 1370 1203 1373 1223
rect 1402 1213 1405 1286
rect 1402 1166 1405 1206
rect 1398 1163 1405 1166
rect 1370 1133 1373 1156
rect 1398 1116 1401 1163
rect 1410 1123 1413 1206
rect 1398 1113 1405 1116
rect 1338 1003 1349 1006
rect 1338 893 1341 986
rect 1346 973 1349 1003
rect 1354 906 1357 1016
rect 1370 983 1373 1006
rect 1394 996 1397 1016
rect 1386 993 1397 996
rect 1378 923 1381 966
rect 1386 933 1389 993
rect 1354 903 1365 906
rect 1314 786 1317 806
rect 1314 783 1325 786
rect 1306 773 1313 776
rect 1210 723 1213 733
rect 1202 703 1213 706
rect 1210 636 1213 703
rect 1242 686 1245 746
rect 1258 743 1269 746
rect 1266 723 1269 743
rect 1310 716 1313 773
rect 1322 723 1325 783
rect 1330 723 1333 806
rect 1310 713 1317 716
rect 1242 683 1253 686
rect 1202 633 1213 636
rect 1202 606 1205 633
rect 1186 593 1189 606
rect 1194 603 1205 606
rect 1210 603 1213 616
rect 1170 573 1181 576
rect 1178 486 1181 573
rect 1194 523 1197 603
rect 1250 586 1253 683
rect 1314 656 1317 713
rect 1338 706 1341 806
rect 1346 773 1349 846
rect 1362 836 1365 903
rect 1354 833 1365 836
rect 1354 803 1357 833
rect 1362 803 1365 816
rect 1334 703 1341 706
rect 1314 653 1325 656
rect 1298 603 1301 616
rect 1242 583 1253 586
rect 1218 533 1221 546
rect 1162 483 1181 486
rect 1162 466 1165 483
rect 1158 463 1165 466
rect 1098 373 1101 396
rect 1114 333 1117 416
rect 1158 406 1161 463
rect 1130 383 1133 406
rect 1158 403 1165 406
rect 1050 323 1069 326
rect 1058 263 1061 306
rect 1074 303 1077 316
rect 1106 283 1109 326
rect 1114 313 1117 326
rect 1034 233 1045 236
rect 1026 193 1029 216
rect 1034 206 1037 233
rect 1050 223 1053 236
rect 1034 203 1045 206
rect 1050 203 1053 216
rect 1066 213 1069 226
rect 1090 213 1093 236
rect 1098 213 1101 226
rect 1114 213 1117 236
rect 1122 213 1125 366
rect 1130 313 1133 346
rect 1146 333 1157 336
rect 1138 233 1141 326
rect 1146 303 1149 326
rect 1154 293 1157 316
rect 1162 286 1165 403
rect 1154 283 1165 286
rect 1170 283 1173 446
rect 1178 403 1181 416
rect 1226 413 1229 506
rect 1242 403 1245 583
rect 1322 576 1325 653
rect 1334 626 1337 703
rect 1334 623 1341 626
rect 1338 606 1341 623
rect 1346 616 1349 756
rect 1370 723 1373 806
rect 1346 613 1365 616
rect 1338 603 1357 606
rect 1362 603 1373 606
rect 1306 573 1325 576
rect 1306 556 1309 573
rect 1354 566 1357 603
rect 1378 586 1381 816
rect 1386 696 1389 856
rect 1394 813 1397 926
rect 1402 906 1405 1113
rect 1418 1056 1421 1373
rect 1434 1356 1437 1376
rect 1442 1363 1445 1406
rect 1466 1393 1469 1416
rect 1474 1366 1477 1876
rect 1506 1816 1509 1973
rect 1514 1953 1517 2006
rect 1530 1983 1533 2006
rect 1554 1996 1557 2126
rect 1562 2013 1565 2126
rect 1550 1993 1557 1996
rect 1530 1916 1533 1966
rect 1490 1813 1509 1816
rect 1522 1913 1533 1916
rect 1482 1783 1485 1806
rect 1466 1363 1477 1366
rect 1430 1353 1437 1356
rect 1430 1286 1433 1353
rect 1466 1316 1469 1363
rect 1482 1323 1485 1776
rect 1490 1713 1493 1746
rect 1506 1676 1509 1806
rect 1522 1796 1525 1913
rect 1538 1896 1541 1946
rect 1534 1893 1541 1896
rect 1534 1826 1537 1893
rect 1550 1886 1553 1993
rect 1562 1943 1565 2006
rect 1570 1953 1573 2193
rect 1578 2113 1581 2223
rect 1594 2216 1597 2256
rect 1586 2213 1597 2216
rect 1586 2123 1589 2213
rect 1594 2193 1597 2206
rect 1602 2163 1605 2216
rect 1610 2183 1613 2206
rect 1618 2156 1621 2326
rect 1594 2153 1621 2156
rect 1594 2123 1597 2153
rect 1602 2143 1621 2146
rect 1602 2133 1605 2143
rect 1594 2066 1597 2086
rect 1594 2063 1601 2066
rect 1578 2003 1581 2036
rect 1546 1883 1553 1886
rect 1534 1823 1541 1826
rect 1538 1803 1541 1823
rect 1490 1673 1509 1676
rect 1514 1793 1525 1796
rect 1466 1313 1485 1316
rect 1430 1283 1437 1286
rect 1426 1213 1429 1226
rect 1414 1053 1421 1056
rect 1414 986 1417 1053
rect 1414 983 1421 986
rect 1410 923 1413 966
rect 1402 903 1409 906
rect 1406 846 1409 903
rect 1402 843 1409 846
rect 1418 843 1421 983
rect 1434 976 1437 1283
rect 1442 1193 1445 1216
rect 1450 1206 1453 1226
rect 1458 1213 1461 1256
rect 1450 1203 1461 1206
rect 1442 1136 1445 1156
rect 1442 1133 1449 1136
rect 1446 1036 1449 1133
rect 1426 973 1437 976
rect 1442 1033 1449 1036
rect 1426 933 1429 973
rect 1434 853 1437 956
rect 1442 893 1445 1033
rect 1458 1016 1461 1203
rect 1466 1123 1469 1246
rect 1474 1203 1477 1236
rect 1482 1196 1485 1313
rect 1490 1306 1493 1673
rect 1514 1653 1517 1793
rect 1522 1723 1525 1786
rect 1498 1613 1501 1646
rect 1522 1636 1525 1716
rect 1530 1643 1533 1726
rect 1538 1663 1541 1786
rect 1546 1746 1549 1883
rect 1554 1753 1557 1806
rect 1562 1773 1565 1936
rect 1578 1803 1581 1986
rect 1598 1976 1601 2063
rect 1610 1983 1613 2136
rect 1618 2123 1621 2143
rect 1626 2133 1629 2206
rect 1618 2003 1621 2116
rect 1634 2083 1637 2326
rect 1658 2253 1661 2406
rect 1666 2323 1669 2416
rect 1674 2396 1677 2536
rect 1690 2513 1693 2526
rect 1698 2523 1701 2616
rect 1710 2566 1713 2763
rect 1722 2743 1725 3036
rect 1738 3013 1741 3026
rect 1738 2923 1741 3006
rect 1746 2976 1749 3093
rect 1762 3026 1765 3066
rect 1770 3033 1773 3173
rect 1786 3096 1789 3296
rect 1794 3193 1797 3403
rect 1810 3396 1813 3466
rect 1834 3413 1837 3703
rect 1842 3603 1845 3626
rect 1850 3446 1853 3616
rect 1858 3613 1861 3726
rect 1858 3593 1861 3606
rect 1866 3603 1869 3786
rect 1874 3613 1877 3746
rect 1874 3596 1877 3606
rect 1866 3593 1877 3596
rect 1858 3513 1861 3526
rect 1866 3463 1869 3593
rect 1882 3586 1885 3646
rect 1890 3623 1893 4016
rect 1898 3796 1901 4140
rect 1914 4056 1917 4140
rect 1914 4053 1921 4056
rect 1918 3996 1921 4053
rect 1914 3993 1921 3996
rect 1914 3973 1917 3993
rect 1930 3966 1933 4140
rect 1946 4056 1949 4140
rect 1938 4053 1949 4056
rect 1938 4013 1941 4053
rect 1970 4033 1973 4140
rect 1986 4036 1989 4140
rect 2002 4053 2005 4140
rect 2018 4043 2021 4140
rect 1978 4033 1989 4036
rect 1914 3963 1933 3966
rect 1906 3813 1909 3926
rect 1898 3793 1905 3796
rect 1902 3726 1905 3793
rect 1898 3723 1905 3726
rect 1914 3723 1917 3963
rect 1938 3933 1941 3946
rect 1954 3876 1957 3976
rect 1962 3956 1965 4006
rect 1978 3966 1981 4033
rect 2018 4013 2021 4036
rect 2026 4006 2029 4056
rect 1994 3993 1997 4006
rect 2018 4003 2029 4006
rect 1978 3963 1997 3966
rect 1962 3953 1973 3956
rect 1946 3873 1957 3876
rect 1922 3743 1925 3846
rect 1946 3776 1949 3873
rect 1970 3856 1973 3953
rect 1962 3853 1973 3856
rect 1962 3796 1965 3853
rect 1994 3846 1997 3963
rect 2002 3926 2005 3946
rect 2002 3923 2009 3926
rect 2018 3923 2021 4003
rect 2006 3846 2009 3923
rect 1986 3843 1997 3846
rect 2002 3843 2009 3846
rect 1962 3793 1973 3796
rect 1946 3773 1957 3776
rect 1898 3643 1901 3723
rect 1890 3596 1893 3616
rect 1898 3603 1901 3636
rect 1906 3596 1909 3606
rect 1890 3593 1909 3596
rect 1846 3443 1853 3446
rect 1802 3393 1813 3396
rect 1846 3396 1849 3443
rect 1846 3393 1853 3396
rect 1874 3393 1877 3586
rect 1882 3583 1901 3586
rect 1898 3533 1901 3583
rect 1914 3573 1917 3616
rect 1914 3533 1917 3556
rect 1890 3403 1893 3416
rect 1802 3333 1805 3393
rect 1810 3316 1813 3336
rect 1806 3313 1813 3316
rect 1806 3236 1809 3313
rect 1802 3233 1809 3236
rect 1802 3213 1805 3233
rect 1802 3203 1813 3206
rect 1818 3186 1821 3316
rect 1810 3183 1821 3186
rect 1782 3093 1789 3096
rect 1782 3036 1785 3093
rect 1794 3076 1797 3136
rect 1810 3096 1813 3183
rect 1810 3093 1821 3096
rect 1794 3073 1805 3076
rect 1782 3033 1789 3036
rect 1762 3023 1773 3026
rect 1754 2996 1757 3016
rect 1762 3003 1765 3016
rect 1770 3013 1773 3023
rect 1770 2996 1773 3006
rect 1754 2993 1773 2996
rect 1746 2973 1753 2976
rect 1750 2896 1753 2973
rect 1778 2923 1781 3016
rect 1746 2893 1753 2896
rect 1746 2873 1749 2893
rect 1730 2736 1733 2856
rect 1738 2813 1741 2826
rect 1722 2733 1733 2736
rect 1710 2563 1717 2566
rect 1706 2533 1709 2546
rect 1714 2533 1717 2563
rect 1722 2543 1725 2733
rect 1730 2713 1733 2726
rect 1706 2473 1709 2526
rect 1682 2413 1685 2466
rect 1714 2423 1717 2456
rect 1690 2413 1717 2416
rect 1690 2403 1693 2413
rect 1674 2393 1681 2396
rect 1678 2316 1681 2393
rect 1698 2323 1701 2386
rect 1706 2366 1709 2406
rect 1722 2373 1725 2536
rect 1730 2413 1733 2576
rect 1738 2473 1741 2796
rect 1738 2413 1741 2466
rect 1706 2363 1717 2366
rect 1674 2313 1681 2316
rect 1642 2033 1645 2216
rect 1650 2206 1653 2216
rect 1658 2213 1661 2246
rect 1674 2236 1677 2313
rect 1714 2306 1717 2363
rect 1730 2356 1733 2406
rect 1746 2383 1749 2736
rect 1754 2723 1757 2736
rect 1754 2633 1757 2716
rect 1762 2663 1765 2816
rect 1778 2813 1781 2826
rect 1786 2806 1789 3033
rect 1794 3013 1797 3026
rect 1802 3003 1805 3073
rect 1818 3023 1821 3093
rect 1810 2996 1813 3016
rect 1818 3003 1821 3016
rect 1826 3013 1829 3346
rect 1834 3223 1837 3326
rect 1842 3133 1845 3326
rect 1826 2996 1829 3006
rect 1810 2993 1829 2996
rect 1794 2863 1797 2986
rect 1794 2813 1797 2826
rect 1778 2803 1789 2806
rect 1770 2656 1773 2786
rect 1778 2713 1781 2803
rect 1794 2796 1797 2806
rect 1802 2803 1805 2836
rect 1810 2796 1813 2816
rect 1818 2813 1821 2946
rect 1834 2933 1837 3016
rect 1842 3013 1845 3126
rect 1834 2903 1837 2926
rect 1842 2906 1845 2936
rect 1850 2933 1853 3393
rect 1898 3323 1901 3526
rect 1922 3523 1925 3646
rect 1930 3503 1933 3626
rect 1938 3583 1941 3746
rect 1954 3736 1957 3773
rect 1970 3743 1973 3793
rect 1954 3733 1969 3736
rect 1954 3646 1957 3726
rect 1966 3686 1969 3733
rect 1966 3683 1973 3686
rect 1954 3643 1965 3646
rect 1946 3613 1949 3626
rect 1954 3613 1957 3636
rect 1962 3606 1965 3643
rect 1946 3603 1965 3606
rect 1938 3436 1941 3576
rect 1946 3493 1949 3603
rect 1962 3533 1965 3596
rect 1970 3546 1973 3683
rect 1986 3633 1989 3843
rect 1986 3613 1989 3626
rect 1970 3543 1989 3546
rect 1954 3513 1957 3526
rect 1962 3523 1973 3526
rect 1962 3446 1965 3523
rect 1978 3513 1981 3536
rect 1962 3443 1969 3446
rect 1922 3433 1941 3436
rect 1922 3356 1925 3433
rect 1938 3393 1941 3406
rect 1966 3396 1969 3443
rect 1978 3413 1981 3506
rect 1986 3406 1989 3543
rect 1994 3483 1997 3836
rect 2002 3723 2005 3843
rect 2010 3813 2013 3826
rect 2034 3823 2037 4140
rect 2050 4056 2053 4140
rect 2042 4053 2053 4056
rect 2042 3833 2045 4053
rect 2066 4026 2069 4140
rect 2062 4023 2069 4026
rect 2062 3966 2065 4023
rect 2062 3963 2069 3966
rect 2074 3963 2077 4016
rect 2066 3943 2069 3963
rect 2082 3943 2085 4140
rect 2098 4013 2101 4140
rect 2114 4056 2117 4140
rect 2114 4053 2125 4056
rect 2122 4013 2125 4053
rect 2162 4026 2165 4046
rect 2682 4026 2685 4140
rect 2738 4126 2741 4140
rect 2730 4123 2741 4126
rect 2730 4046 2733 4123
rect 2754 4056 2757 4140
rect 2754 4053 2765 4056
rect 2730 4043 2741 4046
rect 2162 4023 2169 4026
rect 2682 4023 2693 4026
rect 2098 3993 2101 4006
rect 2138 3956 2141 4016
rect 2166 3976 2169 4023
rect 2162 3973 2169 3976
rect 2138 3953 2149 3956
rect 2034 3733 2037 3806
rect 2050 3753 2053 3926
rect 2066 3773 2069 3936
rect 2114 3913 2117 3926
rect 2090 3773 2093 3806
rect 2058 3686 2061 3736
rect 2106 3723 2109 3746
rect 2058 3683 2069 3686
rect 2002 3616 2005 3636
rect 2002 3613 2009 3616
rect 2006 3546 2009 3613
rect 2002 3543 2009 3546
rect 2002 3503 2005 3543
rect 2010 3513 2013 3526
rect 2018 3523 2021 3556
rect 2034 3506 2037 3616
rect 2066 3573 2069 3683
rect 2122 3656 2125 3826
rect 2098 3653 2125 3656
rect 2098 3586 2101 3653
rect 2114 3593 2117 3616
rect 2098 3583 2109 3586
rect 2066 3536 2069 3556
rect 2062 3533 2069 3536
rect 2050 3513 2053 3526
rect 2026 3503 2037 3506
rect 2026 3446 2029 3503
rect 2026 3443 2037 3446
rect 1962 3393 1969 3396
rect 1978 3403 1989 3406
rect 1922 3353 1941 3356
rect 1922 3333 1925 3346
rect 1858 3043 1861 3276
rect 1874 3213 1877 3226
rect 1898 3186 1901 3226
rect 1898 3183 1909 3186
rect 1858 3013 1861 3026
rect 1858 2993 1861 3006
rect 1866 2983 1869 3136
rect 1890 3026 1893 3146
rect 1882 3023 1893 3026
rect 1874 2976 1877 3016
rect 1866 2973 1877 2976
rect 1858 2933 1861 2956
rect 1850 2923 1861 2926
rect 1842 2903 1849 2906
rect 1826 2813 1829 2896
rect 1794 2793 1813 2796
rect 1818 2776 1821 2806
rect 1834 2793 1837 2866
rect 1846 2836 1849 2903
rect 1858 2863 1861 2916
rect 1842 2833 1849 2836
rect 1842 2803 1845 2833
rect 1850 2813 1861 2816
rect 1866 2813 1869 2973
rect 1882 2943 1885 3023
rect 1890 2996 1893 3016
rect 1898 3003 1901 3016
rect 1906 3013 1909 3183
rect 1922 3143 1925 3306
rect 1938 3213 1941 3353
rect 1946 3223 1949 3376
rect 1946 3203 1949 3216
rect 1954 3213 1957 3326
rect 1962 3233 1965 3393
rect 1978 3346 1981 3403
rect 1978 3343 1985 3346
rect 1970 3213 1973 3336
rect 1982 3236 1985 3343
rect 2002 3336 2005 3426
rect 2034 3423 2037 3443
rect 2018 3373 2021 3416
rect 1994 3333 2005 3336
rect 1994 3256 1997 3333
rect 2002 3266 2005 3326
rect 2018 3276 2021 3346
rect 2034 3343 2037 3416
rect 2042 3323 2045 3486
rect 2050 3316 2053 3506
rect 2062 3466 2065 3533
rect 2062 3463 2069 3466
rect 2066 3366 2069 3463
rect 2074 3413 2077 3566
rect 2106 3553 2109 3583
rect 2098 3533 2101 3546
rect 2122 3523 2125 3576
rect 2130 3563 2133 3946
rect 2146 3866 2149 3953
rect 2138 3863 2149 3866
rect 2138 3823 2141 3863
rect 2138 3793 2141 3816
rect 2138 3736 2141 3756
rect 2138 3733 2149 3736
rect 2146 3686 2149 3733
rect 2138 3683 2149 3686
rect 2138 3553 2141 3683
rect 2146 3496 2149 3666
rect 2138 3493 2149 3496
rect 2042 3313 2053 3316
rect 2062 3363 2069 3366
rect 2018 3273 2029 3276
rect 2002 3263 2021 3266
rect 1994 3253 2005 3256
rect 1978 3233 1985 3236
rect 1914 3106 1917 3126
rect 1954 3123 1957 3206
rect 1962 3176 1965 3206
rect 1978 3203 1981 3233
rect 1986 3213 1997 3216
rect 1962 3173 1969 3176
rect 1966 3116 1969 3173
rect 2002 3156 2005 3253
rect 2018 3213 2021 3263
rect 2018 3163 2021 3206
rect 2002 3153 2013 3156
rect 1994 3133 1997 3146
rect 1962 3113 1969 3116
rect 1914 3103 1925 3106
rect 1922 3046 1925 3103
rect 1914 3043 1925 3046
rect 1906 2996 1909 3006
rect 1890 2993 1909 2996
rect 1914 2946 1917 3043
rect 1922 3013 1925 3026
rect 1938 3016 1941 3036
rect 1930 2993 1933 3016
rect 1938 3013 1945 3016
rect 1962 3013 1965 3113
rect 1978 3013 1981 3026
rect 1874 2923 1877 2936
rect 1898 2933 1901 2946
rect 1914 2943 1933 2946
rect 1882 2913 1885 2926
rect 1922 2913 1925 2926
rect 1930 2903 1933 2943
rect 1942 2936 1945 3013
rect 1938 2933 1945 2936
rect 1858 2796 1861 2806
rect 1874 2803 1877 2816
rect 1842 2793 1861 2796
rect 1802 2773 1821 2776
rect 1786 2676 1789 2726
rect 1794 2706 1797 2766
rect 1802 2723 1805 2773
rect 1810 2713 1813 2726
rect 1826 2723 1829 2756
rect 1834 2706 1837 2786
rect 1794 2703 1801 2706
rect 1762 2653 1773 2656
rect 1778 2673 1789 2676
rect 1778 2653 1781 2673
rect 1762 2573 1765 2653
rect 1798 2636 1801 2703
rect 1770 2536 1773 2616
rect 1778 2613 1781 2626
rect 1754 2523 1757 2536
rect 1770 2533 1781 2536
rect 1754 2403 1757 2496
rect 1762 2413 1765 2516
rect 1770 2463 1773 2526
rect 1778 2493 1781 2533
rect 1786 2516 1789 2636
rect 1794 2633 1801 2636
rect 1826 2703 1837 2706
rect 1826 2636 1829 2703
rect 1842 2643 1845 2793
rect 1882 2716 1885 2866
rect 1938 2833 1941 2933
rect 1978 2923 1981 2956
rect 2010 2953 2013 3153
rect 2026 3086 2029 3273
rect 2034 3173 2037 3236
rect 2042 3196 2045 3313
rect 2062 3286 2065 3363
rect 2114 3353 2117 3406
rect 2090 3333 2109 3336
rect 2062 3283 2069 3286
rect 2066 3213 2069 3283
rect 2082 3213 2085 3246
rect 2090 3213 2093 3333
rect 2098 3283 2101 3326
rect 2106 3323 2109 3333
rect 2114 3246 2117 3346
rect 2130 3333 2133 3416
rect 2138 3413 2141 3493
rect 2154 3403 2157 3606
rect 2162 3476 2165 3973
rect 2178 3846 2181 4016
rect 2186 3863 2189 4016
rect 2194 3963 2197 4006
rect 2202 4003 2205 4016
rect 2234 3976 2237 4016
rect 2218 3973 2237 3976
rect 2194 3893 2197 3926
rect 2210 3866 2213 3936
rect 2218 3933 2221 3973
rect 2234 3926 2237 3966
rect 2242 3933 2245 4006
rect 2282 3966 2285 4006
rect 2314 3993 2317 4006
rect 2274 3963 2285 3966
rect 2202 3863 2213 3866
rect 2226 3923 2237 3926
rect 2178 3843 2189 3846
rect 2186 3766 2189 3843
rect 2178 3763 2189 3766
rect 2202 3766 2205 3863
rect 2226 3856 2229 3923
rect 2250 3903 2253 3926
rect 2218 3853 2229 3856
rect 2218 3783 2221 3853
rect 2202 3763 2213 3766
rect 2178 3746 2181 3763
rect 2174 3743 2181 3746
rect 2174 3656 2177 3743
rect 2174 3653 2181 3656
rect 2178 3633 2181 3653
rect 2170 3563 2173 3616
rect 2178 3566 2181 3626
rect 2186 3583 2189 3736
rect 2202 3733 2205 3746
rect 2210 3726 2213 3763
rect 2226 3743 2229 3816
rect 2234 3793 2237 3806
rect 2194 3703 2197 3726
rect 2202 3723 2213 3726
rect 2194 3573 2197 3616
rect 2202 3613 2205 3723
rect 2210 3613 2213 3716
rect 2218 3616 2221 3736
rect 2242 3733 2245 3836
rect 2250 3793 2253 3866
rect 2258 3813 2261 3926
rect 2266 3813 2269 3896
rect 2258 3783 2261 3806
rect 2274 3733 2277 3963
rect 2314 3923 2317 3946
rect 2290 3803 2293 3916
rect 2226 3723 2253 3726
rect 2226 3663 2229 3723
rect 2298 3656 2301 3846
rect 2306 3793 2309 3806
rect 2314 3803 2317 3816
rect 2294 3653 2301 3656
rect 2218 3613 2229 3616
rect 2202 3593 2205 3606
rect 2178 3563 2197 3566
rect 2170 3523 2173 3546
rect 2186 3476 2189 3556
rect 2162 3473 2173 3476
rect 2170 3396 2173 3473
rect 2162 3393 2173 3396
rect 2182 3473 2189 3476
rect 2162 3343 2165 3393
rect 2182 3356 2185 3473
rect 2194 3366 2197 3563
rect 2202 3403 2205 3526
rect 2210 3413 2213 3566
rect 2218 3553 2221 3613
rect 2226 3533 2229 3606
rect 2218 3413 2221 3526
rect 2234 3416 2237 3636
rect 2250 3593 2253 3606
rect 2242 3533 2245 3546
rect 2258 3533 2261 3546
rect 2250 3493 2253 3526
rect 2234 3413 2245 3416
rect 2194 3363 2201 3366
rect 2182 3353 2189 3356
rect 2162 3276 2165 3336
rect 2106 3243 2117 3246
rect 2158 3273 2165 3276
rect 2042 3193 2053 3196
rect 2050 3123 2053 3193
rect 2066 3183 2069 3206
rect 2026 3083 2037 3086
rect 1890 2723 1893 2816
rect 1898 2733 1901 2816
rect 1922 2753 1925 2816
rect 1930 2763 1933 2806
rect 1882 2713 1893 2716
rect 1826 2633 1837 2636
rect 1858 2633 1861 2646
rect 1794 2613 1797 2633
rect 1802 2613 1813 2616
rect 1826 2606 1829 2616
rect 1802 2603 1829 2606
rect 1834 2603 1837 2633
rect 1826 2583 1829 2603
rect 1842 2566 1845 2626
rect 1866 2613 1869 2636
rect 1874 2623 1877 2656
rect 1882 2623 1885 2706
rect 1890 2606 1893 2713
rect 1922 2693 1925 2736
rect 1938 2723 1941 2816
rect 1946 2803 1949 2916
rect 1946 2716 1949 2746
rect 1954 2736 1957 2876
rect 1994 2866 1997 2946
rect 2034 2943 2037 3083
rect 2058 3073 2061 3176
rect 2042 2926 2045 2956
rect 2018 2913 2021 2926
rect 2034 2923 2045 2926
rect 1970 2863 1997 2866
rect 2034 2866 2037 2923
rect 2058 2886 2061 3046
rect 2066 2913 2069 3166
rect 2074 3013 2077 3176
rect 2082 2983 2085 3076
rect 2090 3053 2093 3206
rect 2098 3153 2101 3216
rect 2106 3173 2109 3243
rect 2114 3193 2117 3206
rect 2106 3063 2109 3126
rect 2114 3106 2117 3186
rect 2130 3183 2133 3206
rect 2158 3196 2161 3273
rect 2154 3193 2161 3196
rect 2138 3133 2141 3156
rect 2114 3103 2125 3106
rect 2122 3046 2125 3103
rect 2154 3066 2157 3193
rect 2170 3166 2173 3286
rect 2186 3253 2189 3353
rect 2198 3316 2201 3363
rect 2234 3356 2237 3406
rect 2242 3363 2245 3413
rect 2250 3403 2253 3426
rect 2234 3353 2245 3356
rect 2210 3323 2213 3346
rect 2242 3323 2245 3353
rect 2258 3323 2261 3416
rect 2266 3403 2269 3586
rect 2274 3523 2277 3566
rect 2282 3533 2285 3616
rect 2294 3576 2297 3653
rect 2294 3573 2301 3576
rect 2298 3556 2301 3573
rect 2298 3553 2317 3556
rect 2298 3533 2301 3546
rect 2282 3413 2285 3476
rect 2290 3463 2293 3526
rect 2306 3513 2309 3536
rect 2314 3496 2317 3553
rect 2322 3503 2325 3616
rect 2330 3583 2333 3756
rect 2338 3733 2341 3996
rect 2362 3993 2365 4016
rect 2418 3983 2421 4016
rect 2354 3923 2357 3936
rect 2370 3933 2373 3946
rect 2394 3933 2397 3946
rect 2362 3833 2365 3926
rect 2378 3826 2381 3926
rect 2402 3923 2405 3936
rect 2426 3933 2429 3996
rect 2418 3843 2421 3926
rect 2434 3906 2437 3986
rect 2442 3973 2445 4006
rect 2442 3933 2445 3946
rect 2450 3923 2453 3936
rect 2474 3923 2477 3936
rect 2482 3933 2485 4016
rect 2498 3933 2501 3946
rect 2530 3933 2533 4016
rect 2586 3956 2589 4006
rect 2610 3996 2613 4016
rect 2602 3993 2613 3996
rect 2586 3953 2597 3956
rect 2546 3906 2549 3926
rect 2430 3903 2437 3906
rect 2430 3836 2433 3903
rect 2430 3833 2437 3836
rect 2362 3823 2381 3826
rect 2362 3816 2365 3823
rect 2354 3813 2365 3816
rect 2354 3793 2357 3813
rect 2362 3783 2365 3806
rect 2346 3733 2349 3746
rect 2370 3723 2373 3816
rect 2378 3753 2381 3806
rect 2378 3676 2381 3736
rect 2386 3693 2389 3816
rect 2394 3803 2397 3816
rect 2394 3733 2397 3796
rect 2402 3783 2405 3826
rect 2402 3733 2405 3746
rect 2410 3723 2413 3816
rect 2378 3673 2397 3676
rect 2330 3506 2333 3576
rect 2338 3523 2341 3606
rect 2346 3563 2349 3616
rect 2354 3553 2357 3606
rect 2362 3603 2365 3616
rect 2370 3593 2373 3606
rect 2354 3543 2373 3546
rect 2354 3536 2357 3543
rect 2346 3533 2357 3536
rect 2354 3513 2357 3526
rect 2330 3503 2337 3506
rect 2314 3493 2325 3496
rect 2194 3313 2201 3316
rect 2194 3293 2197 3313
rect 2178 3193 2181 3216
rect 2170 3163 2181 3166
rect 2170 3123 2173 3156
rect 2154 3063 2165 3066
rect 2114 3043 2125 3046
rect 2114 3026 2117 3043
rect 2098 3023 2117 3026
rect 2050 2883 2061 2886
rect 2034 2863 2045 2866
rect 1970 2805 1973 2863
rect 1954 2733 1973 2736
rect 1938 2713 1949 2716
rect 1898 2613 1901 2626
rect 1906 2623 1909 2636
rect 1922 2633 1925 2656
rect 1930 2606 1933 2626
rect 1834 2563 1845 2566
rect 1866 2603 1893 2606
rect 1922 2603 1933 2606
rect 1834 2546 1837 2563
rect 1866 2556 1869 2603
rect 1794 2543 1821 2546
rect 1794 2533 1797 2543
rect 1802 2533 1813 2536
rect 1786 2513 1797 2516
rect 1810 2513 1813 2526
rect 1770 2413 1773 2456
rect 1778 2413 1781 2476
rect 1794 2446 1797 2513
rect 1786 2443 1797 2446
rect 1818 2446 1821 2543
rect 1830 2543 1837 2546
rect 1862 2553 1869 2556
rect 1830 2486 1833 2543
rect 1850 2513 1853 2526
rect 1862 2496 1865 2553
rect 1858 2493 1865 2496
rect 1830 2483 1837 2486
rect 1818 2443 1825 2446
rect 1770 2373 1773 2406
rect 1710 2303 1717 2306
rect 1722 2353 1733 2356
rect 1710 2236 1713 2303
rect 1674 2233 1701 2236
rect 1710 2233 1717 2236
rect 1650 2203 1661 2206
rect 1594 1973 1601 1976
rect 1586 1756 1589 1816
rect 1594 1783 1597 1973
rect 1602 1923 1605 1946
rect 1626 1806 1629 2026
rect 1634 1946 1637 2006
rect 1642 1963 1645 2016
rect 1650 2003 1653 2176
rect 1658 2003 1661 2203
rect 1666 2193 1669 2206
rect 1674 2196 1677 2216
rect 1682 2203 1685 2216
rect 1690 2213 1693 2226
rect 1690 2196 1693 2206
rect 1674 2193 1693 2196
rect 1666 2166 1669 2186
rect 1698 2173 1701 2233
rect 1666 2163 1673 2166
rect 1670 2056 1673 2163
rect 1698 2083 1701 2166
rect 1706 2123 1709 2216
rect 1714 2213 1717 2233
rect 1714 2193 1717 2206
rect 1722 2186 1725 2353
rect 1738 2333 1741 2346
rect 1778 2336 1781 2406
rect 1770 2333 1781 2336
rect 1714 2183 1725 2186
rect 1714 2106 1717 2183
rect 1738 2163 1741 2326
rect 1770 2243 1773 2333
rect 1778 2313 1781 2326
rect 1738 2133 1741 2146
rect 1710 2103 1717 2106
rect 1666 2053 1673 2056
rect 1634 1943 1645 1946
rect 1634 1903 1637 1936
rect 1618 1803 1629 1806
rect 1586 1753 1597 1756
rect 1546 1743 1557 1746
rect 1546 1643 1549 1736
rect 1522 1633 1541 1636
rect 1522 1613 1533 1616
rect 1498 1523 1501 1536
rect 1514 1483 1517 1576
rect 1498 1313 1501 1326
rect 1490 1303 1497 1306
rect 1494 1236 1497 1303
rect 1506 1246 1509 1386
rect 1522 1336 1525 1606
rect 1530 1523 1533 1576
rect 1538 1553 1541 1633
rect 1538 1523 1541 1536
rect 1546 1523 1549 1636
rect 1554 1623 1557 1743
rect 1570 1743 1589 1746
rect 1562 1633 1565 1736
rect 1570 1723 1573 1743
rect 1578 1713 1581 1736
rect 1586 1733 1589 1743
rect 1554 1533 1557 1616
rect 1562 1573 1565 1606
rect 1538 1436 1541 1456
rect 1562 1453 1565 1556
rect 1534 1433 1541 1436
rect 1534 1356 1537 1433
rect 1546 1413 1549 1426
rect 1554 1396 1557 1446
rect 1562 1403 1565 1436
rect 1554 1393 1565 1396
rect 1534 1353 1541 1356
rect 1538 1336 1541 1353
rect 1518 1333 1525 1336
rect 1530 1333 1541 1336
rect 1518 1266 1521 1333
rect 1518 1263 1525 1266
rect 1506 1243 1513 1246
rect 1494 1233 1501 1236
rect 1474 1193 1485 1196
rect 1450 933 1453 1016
rect 1458 1013 1469 1016
rect 1474 1013 1477 1193
rect 1490 1173 1493 1216
rect 1458 983 1461 1006
rect 1466 976 1469 1013
rect 1458 973 1469 976
rect 1458 953 1461 973
rect 1466 946 1469 966
rect 1490 963 1493 1156
rect 1498 1093 1501 1233
rect 1510 1156 1513 1243
rect 1522 1213 1525 1263
rect 1530 1193 1533 1333
rect 1506 1153 1513 1156
rect 1506 1013 1509 1153
rect 1514 1116 1517 1136
rect 1530 1133 1533 1166
rect 1514 1113 1525 1116
rect 1498 1003 1509 1006
rect 1458 943 1469 946
rect 1402 803 1405 843
rect 1418 776 1421 806
rect 1434 776 1437 796
rect 1418 773 1437 776
rect 1450 773 1453 866
rect 1410 733 1413 746
rect 1386 693 1397 696
rect 1394 613 1397 693
rect 1434 656 1437 773
rect 1458 743 1461 943
rect 1466 813 1469 826
rect 1482 733 1485 936
rect 1514 923 1517 1016
rect 1522 1003 1525 1113
rect 1538 1073 1541 1326
rect 1546 1323 1549 1376
rect 1546 1026 1549 1296
rect 1554 1033 1557 1336
rect 1562 1316 1565 1393
rect 1570 1333 1573 1666
rect 1578 1603 1581 1616
rect 1586 1613 1589 1726
rect 1594 1713 1597 1753
rect 1602 1723 1605 1776
rect 1618 1766 1621 1803
rect 1614 1763 1621 1766
rect 1614 1706 1617 1763
rect 1610 1703 1617 1706
rect 1610 1636 1613 1703
rect 1626 1656 1629 1796
rect 1634 1723 1637 1816
rect 1642 1756 1645 1943
rect 1650 1923 1653 1946
rect 1658 1903 1661 1996
rect 1666 1933 1669 2053
rect 1710 2036 1713 2103
rect 1674 1993 1677 2036
rect 1710 2033 1717 2036
rect 1690 2016 1693 2026
rect 1682 2013 1693 2016
rect 1642 1753 1653 1756
rect 1642 1713 1645 1736
rect 1626 1653 1645 1656
rect 1610 1633 1621 1636
rect 1578 1553 1581 1596
rect 1586 1433 1589 1526
rect 1578 1413 1581 1426
rect 1594 1403 1597 1606
rect 1602 1523 1605 1616
rect 1618 1546 1621 1633
rect 1626 1613 1629 1646
rect 1634 1603 1637 1636
rect 1610 1543 1621 1546
rect 1610 1473 1613 1543
rect 1618 1503 1621 1536
rect 1634 1533 1637 1576
rect 1634 1463 1637 1526
rect 1634 1436 1637 1456
rect 1630 1433 1637 1436
rect 1618 1413 1621 1426
rect 1562 1313 1573 1316
rect 1586 1313 1589 1326
rect 1570 1246 1573 1313
rect 1562 1243 1573 1246
rect 1562 1133 1565 1243
rect 1578 1203 1581 1216
rect 1602 1213 1605 1336
rect 1630 1316 1633 1433
rect 1630 1313 1637 1316
rect 1634 1293 1637 1313
rect 1642 1263 1645 1653
rect 1650 1593 1653 1753
rect 1658 1546 1661 1726
rect 1666 1603 1669 1876
rect 1674 1863 1677 1936
rect 1682 1923 1685 2013
rect 1682 1786 1685 1906
rect 1690 1793 1693 1936
rect 1698 1933 1701 2006
rect 1706 1923 1709 2016
rect 1714 2003 1717 2033
rect 1722 1943 1725 2096
rect 1730 1936 1733 2086
rect 1714 1906 1717 1936
rect 1710 1903 1717 1906
rect 1722 1933 1733 1936
rect 1674 1783 1685 1786
rect 1698 1783 1701 1856
rect 1710 1836 1713 1903
rect 1710 1833 1717 1836
rect 1674 1766 1677 1783
rect 1674 1763 1685 1766
rect 1682 1676 1685 1763
rect 1706 1733 1709 1816
rect 1714 1743 1717 1833
rect 1674 1673 1685 1676
rect 1674 1586 1677 1673
rect 1650 1543 1661 1546
rect 1670 1583 1677 1586
rect 1650 1523 1653 1543
rect 1670 1516 1673 1583
rect 1666 1513 1673 1516
rect 1666 1453 1669 1513
rect 1666 1366 1669 1416
rect 1674 1413 1677 1506
rect 1682 1443 1685 1656
rect 1698 1643 1709 1646
rect 1698 1603 1701 1643
rect 1714 1626 1717 1716
rect 1722 1653 1725 1933
rect 1730 1726 1733 1926
rect 1738 1853 1741 2116
rect 1754 2106 1757 2216
rect 1762 2213 1773 2216
rect 1778 2213 1781 2226
rect 1770 2186 1773 2206
rect 1750 2103 1757 2106
rect 1762 2183 1773 2186
rect 1778 2183 1781 2206
rect 1750 2026 1753 2103
rect 1762 2066 1765 2183
rect 1770 2113 1773 2176
rect 1786 2173 1789 2443
rect 1794 2413 1797 2426
rect 1810 2403 1813 2436
rect 1822 2396 1825 2443
rect 1818 2393 1825 2396
rect 1818 2336 1821 2393
rect 1802 2333 1821 2336
rect 1802 2276 1805 2333
rect 1818 2293 1821 2326
rect 1826 2313 1829 2326
rect 1798 2273 1805 2276
rect 1798 2186 1801 2273
rect 1798 2183 1805 2186
rect 1794 2093 1797 2166
rect 1802 2086 1805 2183
rect 1810 2096 1813 2276
rect 1818 2123 1821 2216
rect 1834 2163 1837 2483
rect 1858 2436 1861 2493
rect 1858 2433 1869 2436
rect 1866 2413 1869 2433
rect 1842 2273 1845 2346
rect 1850 2323 1853 2406
rect 1866 2326 1869 2406
rect 1874 2393 1877 2546
rect 1898 2533 1901 2576
rect 1922 2546 1925 2603
rect 1938 2566 1941 2706
rect 1946 2643 1949 2706
rect 1946 2613 1949 2626
rect 1954 2613 1957 2726
rect 1962 2616 1965 2716
rect 1970 2713 1973 2733
rect 1962 2613 1973 2616
rect 1938 2563 1949 2566
rect 1922 2543 1933 2546
rect 1914 2476 1917 2526
rect 1914 2473 1921 2476
rect 1882 2373 1885 2416
rect 1898 2413 1901 2426
rect 1906 2416 1909 2466
rect 1918 2426 1921 2473
rect 1930 2456 1933 2543
rect 1946 2473 1949 2563
rect 1954 2463 1957 2596
rect 1930 2453 1949 2456
rect 1918 2423 1925 2426
rect 1906 2413 1917 2416
rect 1890 2403 1909 2406
rect 1914 2386 1917 2413
rect 1922 2403 1925 2423
rect 1930 2403 1933 2426
rect 1906 2383 1917 2386
rect 1874 2343 1893 2346
rect 1874 2333 1877 2343
rect 1882 2326 1885 2336
rect 1866 2323 1885 2326
rect 1890 2323 1893 2343
rect 1866 2296 1869 2316
rect 1842 2183 1845 2216
rect 1850 2193 1853 2206
rect 1842 2113 1845 2146
rect 1858 2133 1861 2296
rect 1866 2293 1877 2296
rect 1898 2293 1901 2336
rect 1906 2333 1909 2383
rect 1914 2316 1917 2376
rect 1910 2313 1917 2316
rect 1874 2236 1877 2293
rect 1866 2233 1877 2236
rect 1910 2236 1913 2313
rect 1910 2233 1917 2236
rect 1866 2173 1869 2233
rect 1882 2176 1885 2216
rect 1898 2213 1901 2226
rect 1914 2216 1917 2233
rect 1906 2213 1917 2216
rect 1882 2173 1901 2176
rect 1858 2106 1861 2126
rect 1850 2103 1861 2106
rect 1810 2093 1829 2096
rect 1802 2083 1821 2086
rect 1762 2063 1773 2066
rect 1746 2023 1753 2026
rect 1746 1933 1749 2023
rect 1754 2003 1765 2006
rect 1770 2003 1773 2063
rect 1794 1943 1797 2036
rect 1802 1936 1805 2006
rect 1810 1973 1813 2016
rect 1818 2003 1821 2083
rect 1826 2003 1829 2093
rect 1850 2016 1853 2103
rect 1850 2013 1857 2016
rect 1866 2013 1869 2126
rect 1874 2023 1877 2136
rect 1890 2133 1893 2146
rect 1898 2133 1901 2173
rect 1906 2133 1909 2213
rect 1882 2033 1885 2126
rect 1906 2113 1909 2126
rect 1914 2123 1917 2206
rect 1898 2013 1901 2036
rect 1754 1896 1757 1936
rect 1762 1903 1765 1926
rect 1754 1893 1773 1896
rect 1746 1803 1749 1816
rect 1738 1743 1741 1756
rect 1754 1736 1757 1806
rect 1750 1733 1757 1736
rect 1730 1723 1741 1726
rect 1714 1623 1725 1626
rect 1706 1576 1709 1616
rect 1714 1593 1717 1616
rect 1690 1573 1709 1576
rect 1690 1533 1693 1573
rect 1690 1406 1693 1516
rect 1698 1506 1701 1536
rect 1722 1533 1725 1623
rect 1730 1603 1733 1616
rect 1738 1536 1741 1723
rect 1750 1656 1753 1733
rect 1750 1653 1757 1656
rect 1754 1633 1757 1653
rect 1762 1546 1765 1846
rect 1770 1813 1773 1893
rect 1778 1853 1781 1936
rect 1802 1933 1813 1936
rect 1802 1903 1805 1926
rect 1786 1773 1789 1816
rect 1778 1733 1781 1746
rect 1770 1706 1773 1726
rect 1770 1703 1777 1706
rect 1774 1626 1777 1703
rect 1786 1663 1789 1736
rect 1794 1733 1797 1846
rect 1810 1793 1813 1933
rect 1842 1876 1845 2006
rect 1854 1946 1857 2013
rect 1834 1873 1845 1876
rect 1850 1943 1857 1946
rect 1834 1736 1837 1873
rect 1850 1836 1853 1943
rect 1858 1843 1861 1926
rect 1850 1833 1861 1836
rect 1834 1733 1845 1736
rect 1850 1733 1853 1816
rect 1858 1793 1861 1833
rect 1866 1803 1869 1826
rect 1858 1733 1861 1756
rect 1794 1656 1797 1726
rect 1802 1673 1805 1726
rect 1794 1653 1801 1656
rect 1770 1623 1777 1626
rect 1770 1603 1773 1623
rect 1778 1593 1781 1606
rect 1762 1543 1773 1546
rect 1734 1533 1741 1536
rect 1706 1523 1725 1526
rect 1698 1503 1709 1506
rect 1706 1416 1709 1503
rect 1722 1423 1725 1516
rect 1706 1413 1717 1416
rect 1666 1363 1673 1366
rect 1650 1323 1653 1346
rect 1670 1306 1673 1363
rect 1682 1323 1685 1406
rect 1690 1403 1709 1406
rect 1714 1396 1717 1413
rect 1706 1393 1717 1396
rect 1722 1393 1725 1416
rect 1734 1406 1737 1533
rect 1746 1413 1749 1526
rect 1762 1516 1765 1536
rect 1758 1513 1765 1516
rect 1758 1456 1761 1513
rect 1758 1453 1765 1456
rect 1762 1436 1765 1453
rect 1770 1443 1773 1543
rect 1786 1533 1789 1626
rect 1798 1556 1801 1653
rect 1810 1573 1813 1696
rect 1798 1553 1813 1556
rect 1786 1493 1789 1516
rect 1762 1433 1773 1436
rect 1730 1403 1737 1406
rect 1666 1303 1673 1306
rect 1618 1203 1621 1216
rect 1562 1093 1565 1126
rect 1602 1076 1605 1136
rect 1594 1073 1605 1076
rect 1538 1023 1549 1026
rect 1522 906 1525 996
rect 1518 903 1525 906
rect 1490 813 1501 816
rect 1506 813 1509 826
rect 1518 806 1521 903
rect 1506 803 1521 806
rect 1506 756 1509 803
rect 1502 753 1509 756
rect 1482 703 1485 726
rect 1502 706 1505 753
rect 1514 723 1517 746
rect 1502 703 1509 706
rect 1522 703 1525 726
rect 1530 706 1533 1016
rect 1538 993 1541 1023
rect 1546 956 1549 1016
rect 1554 976 1557 1006
rect 1562 1003 1565 1016
rect 1578 1013 1581 1036
rect 1554 973 1565 976
rect 1546 953 1553 956
rect 1550 886 1553 953
rect 1562 923 1565 973
rect 1546 883 1553 886
rect 1538 723 1541 816
rect 1546 813 1549 883
rect 1546 796 1549 806
rect 1554 803 1557 816
rect 1562 796 1565 816
rect 1570 803 1573 1006
rect 1594 986 1597 1073
rect 1610 996 1613 1196
rect 1618 1013 1621 1126
rect 1610 993 1617 996
rect 1594 983 1605 986
rect 1586 886 1589 966
rect 1602 953 1605 983
rect 1586 883 1605 886
rect 1578 813 1581 836
rect 1546 793 1565 796
rect 1546 723 1549 776
rect 1554 743 1573 746
rect 1554 733 1557 743
rect 1554 706 1557 726
rect 1530 703 1541 706
rect 1506 683 1509 703
rect 1418 653 1437 656
rect 1386 603 1397 606
rect 1346 563 1357 566
rect 1370 583 1381 586
rect 1306 553 1317 556
rect 1290 523 1293 536
rect 1314 486 1317 553
rect 1346 536 1349 563
rect 1330 533 1349 536
rect 1354 533 1365 536
rect 1330 516 1333 533
rect 1306 483 1317 486
rect 1326 513 1333 516
rect 1338 523 1357 526
rect 1338 513 1341 523
rect 1306 456 1309 483
rect 1306 453 1317 456
rect 1290 393 1293 416
rect 1178 313 1181 336
rect 1186 323 1189 336
rect 1186 293 1189 316
rect 1202 303 1205 326
rect 1210 323 1213 336
rect 1226 333 1229 386
rect 1314 376 1317 453
rect 1326 406 1329 513
rect 1370 506 1373 583
rect 1362 503 1373 506
rect 1338 416 1341 476
rect 1362 436 1365 503
rect 1378 496 1381 576
rect 1402 563 1405 606
rect 1418 566 1421 653
rect 1466 613 1469 626
rect 1410 563 1421 566
rect 1410 523 1413 563
rect 1378 493 1389 496
rect 1386 436 1389 493
rect 1362 433 1373 436
rect 1338 413 1357 416
rect 1370 413 1373 433
rect 1378 433 1389 436
rect 1378 413 1381 433
rect 1326 403 1333 406
rect 1306 373 1317 376
rect 1330 386 1333 403
rect 1346 386 1349 406
rect 1362 393 1365 406
rect 1330 383 1349 386
rect 1378 383 1381 406
rect 1250 293 1253 346
rect 1042 126 1045 203
rect 1090 193 1093 206
rect 1098 203 1109 206
rect 1122 183 1125 206
rect 1042 123 1061 126
rect 1074 123 1077 166
rect 1130 163 1133 206
rect 1138 193 1141 216
rect 1130 123 1133 156
rect 1154 133 1157 283
rect 1162 203 1165 216
rect 1170 193 1173 216
rect 1170 133 1173 176
rect 1178 153 1181 206
rect 1186 193 1189 256
rect 1194 223 1221 226
rect 1194 213 1197 223
rect 1218 216 1221 223
rect 1226 216 1229 236
rect 1194 166 1197 206
rect 1202 203 1205 216
rect 1210 183 1213 216
rect 1218 213 1229 216
rect 1194 163 1205 166
rect 1186 133 1189 146
rect 1202 143 1205 163
rect 1218 123 1221 206
rect 1234 203 1237 256
rect 1242 183 1245 216
rect 1250 126 1253 206
rect 1258 203 1261 216
rect 1266 153 1269 336
rect 1274 323 1277 346
rect 1282 213 1285 236
rect 1290 213 1293 336
rect 1306 263 1309 373
rect 1330 336 1333 383
rect 1386 346 1389 406
rect 1322 333 1333 336
rect 1346 333 1349 346
rect 1362 333 1365 346
rect 1378 343 1389 346
rect 1378 336 1381 343
rect 1370 333 1381 336
rect 1314 323 1341 326
rect 1354 243 1357 326
rect 1378 313 1381 326
rect 1354 213 1357 236
rect 1386 233 1389 336
rect 1394 303 1397 416
rect 1410 413 1413 436
rect 1402 373 1405 406
rect 1410 403 1421 406
rect 1426 393 1429 416
rect 1434 403 1437 486
rect 1410 333 1413 356
rect 1394 253 1397 276
rect 1402 213 1405 316
rect 1410 213 1413 326
rect 1418 323 1421 376
rect 1450 366 1453 526
rect 1458 513 1461 526
rect 1482 383 1485 636
rect 1498 593 1501 616
rect 1506 613 1509 626
rect 1490 523 1493 536
rect 1506 526 1509 566
rect 1514 556 1517 616
rect 1522 613 1525 686
rect 1538 656 1541 703
rect 1530 653 1541 656
rect 1550 703 1557 706
rect 1530 633 1533 653
rect 1550 636 1553 703
rect 1550 633 1557 636
rect 1522 596 1525 606
rect 1530 603 1533 626
rect 1538 596 1541 616
rect 1554 613 1557 633
rect 1562 623 1565 736
rect 1570 723 1573 743
rect 1578 733 1581 746
rect 1586 733 1589 806
rect 1578 723 1589 726
rect 1522 593 1541 596
rect 1546 593 1549 606
rect 1514 553 1525 556
rect 1522 526 1525 553
rect 1530 543 1549 546
rect 1530 533 1533 543
rect 1538 526 1541 536
rect 1498 513 1501 526
rect 1506 523 1517 526
rect 1522 523 1541 526
rect 1546 523 1549 543
rect 1554 533 1557 546
rect 1562 526 1565 616
rect 1570 556 1573 656
rect 1578 583 1581 606
rect 1586 566 1589 666
rect 1594 603 1597 726
rect 1602 613 1605 883
rect 1614 876 1617 993
rect 1610 873 1617 876
rect 1610 853 1613 873
rect 1626 786 1629 1046
rect 1634 923 1637 1016
rect 1642 963 1645 1136
rect 1666 1133 1669 1303
rect 1674 1203 1677 1286
rect 1690 1246 1693 1336
rect 1682 1243 1693 1246
rect 1682 1213 1685 1243
rect 1690 1213 1701 1216
rect 1706 1213 1709 1393
rect 1730 1346 1733 1403
rect 1722 1343 1733 1346
rect 1690 1203 1701 1206
rect 1690 1146 1693 1196
rect 1722 1193 1725 1343
rect 1730 1306 1733 1336
rect 1738 1323 1741 1396
rect 1754 1393 1757 1406
rect 1762 1403 1765 1426
rect 1746 1333 1749 1346
rect 1754 1333 1765 1336
rect 1770 1326 1773 1433
rect 1794 1346 1797 1536
rect 1786 1343 1797 1346
rect 1786 1326 1789 1343
rect 1754 1323 1773 1326
rect 1782 1323 1789 1326
rect 1730 1303 1741 1306
rect 1738 1226 1741 1303
rect 1730 1223 1741 1226
rect 1730 1203 1733 1223
rect 1690 1143 1701 1146
rect 1698 1096 1701 1143
rect 1714 1123 1717 1136
rect 1754 1126 1757 1323
rect 1770 1216 1773 1316
rect 1782 1226 1785 1323
rect 1782 1223 1789 1226
rect 1762 1213 1773 1216
rect 1786 1206 1789 1223
rect 1794 1213 1797 1336
rect 1762 1133 1765 1206
rect 1778 1173 1781 1206
rect 1786 1203 1797 1206
rect 1754 1123 1765 1126
rect 1650 1003 1661 1006
rect 1666 1003 1669 1016
rect 1674 1013 1677 1036
rect 1682 1003 1685 1096
rect 1690 1093 1701 1096
rect 1690 1043 1693 1093
rect 1690 1003 1693 1016
rect 1706 1013 1709 1076
rect 1698 966 1701 1006
rect 1690 963 1701 966
rect 1650 936 1653 956
rect 1650 933 1661 936
rect 1658 886 1661 933
rect 1650 883 1661 886
rect 1622 783 1629 786
rect 1610 703 1613 736
rect 1622 726 1625 783
rect 1622 723 1629 726
rect 1634 723 1637 816
rect 1642 733 1645 806
rect 1650 773 1653 883
rect 1666 756 1669 856
rect 1674 813 1677 936
rect 1690 916 1693 963
rect 1706 923 1709 1006
rect 1714 936 1717 1036
rect 1722 1013 1733 1016
rect 1738 983 1741 1016
rect 1746 1013 1749 1096
rect 1754 1013 1757 1076
rect 1762 1013 1765 1046
rect 1770 1013 1773 1136
rect 1778 1033 1781 1126
rect 1786 1076 1789 1136
rect 1794 1123 1797 1203
rect 1802 1123 1805 1536
rect 1810 1516 1813 1553
rect 1818 1533 1821 1626
rect 1810 1513 1817 1516
rect 1814 1426 1817 1513
rect 1810 1423 1817 1426
rect 1810 1403 1813 1423
rect 1810 1126 1813 1396
rect 1826 1393 1829 1636
rect 1834 1523 1837 1716
rect 1842 1566 1845 1733
rect 1866 1723 1869 1786
rect 1866 1696 1869 1716
rect 1874 1713 1877 1976
rect 1890 1873 1893 2006
rect 1906 1933 1909 2066
rect 1914 1993 1917 2026
rect 1882 1803 1893 1806
rect 1862 1693 1869 1696
rect 1850 1603 1853 1676
rect 1862 1606 1865 1693
rect 1874 1633 1877 1706
rect 1882 1626 1885 1796
rect 1890 1653 1893 1803
rect 1898 1723 1901 1806
rect 1914 1796 1917 1986
rect 1922 1936 1925 2396
rect 1930 2343 1933 2396
rect 1930 2293 1933 2326
rect 1938 2323 1941 2446
rect 1946 2436 1949 2453
rect 1946 2433 1953 2436
rect 1950 2296 1953 2433
rect 1962 2413 1965 2526
rect 1970 2443 1973 2613
rect 1978 2553 1981 2626
rect 1986 2573 1989 2746
rect 1994 2713 1997 2726
rect 2002 2713 2005 2816
rect 2034 2766 2037 2836
rect 2030 2763 2037 2766
rect 1994 2613 1997 2656
rect 2002 2556 2005 2706
rect 2010 2613 2013 2726
rect 2018 2633 2021 2716
rect 2030 2686 2033 2763
rect 2030 2683 2037 2686
rect 2034 2663 2037 2683
rect 2026 2633 2029 2646
rect 2010 2573 2013 2606
rect 2026 2593 2029 2626
rect 2034 2613 2037 2626
rect 2002 2553 2013 2556
rect 2042 2553 2045 2863
rect 2050 2796 2053 2883
rect 2058 2813 2061 2826
rect 2074 2806 2077 2926
rect 2082 2923 2085 2976
rect 2098 2966 2101 3023
rect 2094 2963 2101 2966
rect 2094 2906 2097 2963
rect 2094 2903 2101 2906
rect 2098 2883 2101 2903
rect 2098 2813 2109 2816
rect 2074 2803 2101 2806
rect 2050 2793 2057 2796
rect 2054 2646 2057 2793
rect 2106 2783 2109 2813
rect 2114 2776 2117 3016
rect 2130 2993 2133 3006
rect 2122 2883 2125 2986
rect 2138 2923 2141 2936
rect 2162 2933 2165 3063
rect 2178 3026 2181 3163
rect 2194 3156 2197 3226
rect 2218 3213 2229 3216
rect 2242 3213 2245 3296
rect 2258 3216 2261 3236
rect 2250 3213 2261 3216
rect 2266 3206 2269 3336
rect 2282 3333 2285 3346
rect 2290 3323 2293 3416
rect 2298 3413 2309 3416
rect 2314 3413 2317 3426
rect 2322 3406 2325 3493
rect 2334 3436 2337 3503
rect 2362 3476 2365 3536
rect 2370 3533 2373 3543
rect 2378 3513 2381 3636
rect 2386 3603 2389 3616
rect 2394 3613 2397 3673
rect 2410 3626 2413 3646
rect 2418 3636 2421 3806
rect 2426 3776 2429 3816
rect 2434 3803 2437 3833
rect 2442 3786 2445 3906
rect 2538 3903 2549 3906
rect 2458 3803 2461 3856
rect 2506 3793 2509 3816
rect 2538 3786 2541 3903
rect 2442 3783 2461 3786
rect 2426 3773 2445 3776
rect 2418 3633 2429 3636
rect 2402 3623 2421 3626
rect 2394 3593 2397 3606
rect 2386 3523 2389 3586
rect 2402 3536 2405 3623
rect 2426 3616 2429 3633
rect 2418 3613 2429 3616
rect 2394 3533 2405 3536
rect 2330 3433 2337 3436
rect 2346 3473 2365 3476
rect 2330 3413 2333 3433
rect 2306 3383 2309 3406
rect 2298 3236 2301 3336
rect 2314 3333 2317 3406
rect 2322 3403 2333 3406
rect 2322 3333 2325 3356
rect 2330 3323 2333 3403
rect 2282 3233 2301 3236
rect 2234 3203 2245 3206
rect 2250 3193 2253 3206
rect 2266 3203 2277 3206
rect 2282 3203 2285 3233
rect 2338 3213 2341 3336
rect 2346 3323 2349 3473
rect 2362 3416 2365 3446
rect 2354 3413 2365 3416
rect 2378 3413 2381 3426
rect 2370 3393 2373 3406
rect 2354 3323 2357 3336
rect 2378 3316 2381 3336
rect 2370 3313 2381 3316
rect 2370 3236 2373 3313
rect 2370 3233 2381 3236
rect 2386 3233 2389 3506
rect 2394 3433 2397 3533
rect 2410 3526 2413 3536
rect 2402 3523 2413 3526
rect 2402 3493 2405 3523
rect 2394 3383 2397 3406
rect 2402 3313 2405 3486
rect 2410 3433 2413 3516
rect 2418 3413 2421 3613
rect 2426 3473 2429 3556
rect 2434 3533 2437 3736
rect 2442 3713 2445 3773
rect 2450 3733 2453 3756
rect 2458 3733 2461 3783
rect 2466 3723 2469 3736
rect 2474 3706 2477 3786
rect 2538 3783 2549 3786
rect 2442 3583 2445 3616
rect 2450 3573 2453 3606
rect 2442 3533 2453 3536
rect 2458 3533 2461 3706
rect 2470 3703 2477 3706
rect 2470 3646 2473 3703
rect 2482 3696 2485 3736
rect 2506 3733 2509 3746
rect 2514 3733 2517 3766
rect 2490 3713 2493 3726
rect 2498 3723 2509 3726
rect 2522 3703 2525 3726
rect 2482 3693 2493 3696
rect 2490 3646 2493 3693
rect 2530 3676 2533 3736
rect 2538 3693 2541 3766
rect 2546 3733 2549 3783
rect 2554 3773 2557 3946
rect 2570 3933 2589 3936
rect 2562 3913 2565 3926
rect 2586 3826 2589 3926
rect 2594 3903 2597 3953
rect 2602 3933 2605 3993
rect 2658 3946 2661 4016
rect 2666 4006 2669 4016
rect 2666 4003 2685 4006
rect 2690 4003 2693 4023
rect 2658 3943 2665 3946
rect 2610 3826 2613 3926
rect 2618 3923 2621 3936
rect 2578 3823 2589 3826
rect 2594 3823 2613 3826
rect 2554 3723 2557 3736
rect 2562 3733 2565 3816
rect 2570 3783 2573 3806
rect 2466 3643 2473 3646
rect 2482 3643 2493 3646
rect 2514 3673 2533 3676
rect 2466 3586 2469 3643
rect 2474 3616 2477 3636
rect 2482 3623 2485 3643
rect 2474 3613 2509 3616
rect 2514 3613 2517 3673
rect 2474 3593 2477 3606
rect 2466 3583 2477 3586
rect 2434 3433 2437 3526
rect 2434 3413 2437 3426
rect 2442 3413 2445 3526
rect 2450 3443 2453 3526
rect 2466 3523 2469 3536
rect 2474 3516 2477 3583
rect 2482 3523 2485 3606
rect 2490 3553 2493 3606
rect 2498 3593 2501 3606
rect 2506 3563 2517 3566
rect 2506 3533 2509 3556
rect 2514 3533 2517 3563
rect 2474 3513 2485 3516
rect 2466 3413 2469 3426
rect 2482 3406 2485 3513
rect 2490 3423 2493 3436
rect 2498 3416 2501 3426
rect 2490 3413 2501 3416
rect 2506 3413 2509 3516
rect 2514 3513 2517 3526
rect 2522 3483 2525 3646
rect 2530 3623 2533 3656
rect 2530 3583 2533 3616
rect 2538 3486 2541 3686
rect 2570 3683 2573 3776
rect 2578 3753 2581 3823
rect 2586 3793 2589 3806
rect 2594 3766 2597 3823
rect 2602 3803 2605 3816
rect 2626 3803 2629 3906
rect 2634 3863 2637 3936
rect 2662 3896 2665 3943
rect 2674 3923 2677 3946
rect 2698 3913 2701 4016
rect 2706 3996 2709 4016
rect 2722 4013 2725 4026
rect 2738 4003 2741 4043
rect 2706 3993 2717 3996
rect 2714 3926 2717 3993
rect 2762 3976 2765 4053
rect 2778 3993 2781 4016
rect 2802 4003 2805 4016
rect 2818 4003 2821 4140
rect 2754 3973 2765 3976
rect 2706 3923 2717 3926
rect 2658 3893 2665 3896
rect 2650 3773 2653 3846
rect 2594 3763 2613 3766
rect 2546 3603 2549 3636
rect 2578 3623 2581 3736
rect 2594 3733 2597 3756
rect 2602 3733 2605 3746
rect 2610 3736 2613 3763
rect 2610 3733 2621 3736
rect 2586 3713 2589 3726
rect 2594 3723 2605 3726
rect 2594 3703 2597 3723
rect 2610 3636 2613 3733
rect 2626 3716 2629 3736
rect 2634 3723 2637 3766
rect 2642 3733 2645 3756
rect 2650 3733 2653 3746
rect 2642 3723 2653 3726
rect 2622 3713 2629 3716
rect 2622 3656 2625 3713
rect 2622 3653 2629 3656
rect 2610 3633 2617 3636
rect 2570 3613 2581 3616
rect 2554 3563 2557 3606
rect 2570 3593 2573 3606
rect 2554 3543 2573 3546
rect 2554 3536 2557 3543
rect 2546 3533 2557 3536
rect 2562 3526 2565 3536
rect 2570 3533 2573 3543
rect 2586 3526 2589 3606
rect 2594 3593 2597 3606
rect 2554 3503 2557 3526
rect 2562 3523 2589 3526
rect 2602 3523 2605 3626
rect 2538 3483 2545 3486
rect 2426 3403 2437 3406
rect 2442 3393 2445 3406
rect 2466 3383 2469 3406
rect 2394 3236 2397 3256
rect 2394 3233 2401 3236
rect 2378 3213 2381 3233
rect 2298 3183 2301 3206
rect 2386 3186 2389 3216
rect 2378 3183 2389 3186
rect 2190 3153 2197 3156
rect 2190 3066 2193 3153
rect 2190 3063 2197 3066
rect 2170 3023 2181 3026
rect 2170 2953 2173 3023
rect 2178 2993 2181 3016
rect 2194 2963 2197 3063
rect 2202 2946 2205 3146
rect 2210 3013 2213 3136
rect 2234 3133 2237 3146
rect 2218 3066 2221 3126
rect 2218 3063 2237 3066
rect 2210 2983 2213 3006
rect 2218 2973 2221 3006
rect 2226 3003 2229 3016
rect 2234 3003 2237 3063
rect 2242 3013 2245 3036
rect 2258 3013 2261 3026
rect 2250 2993 2253 3006
rect 2266 2976 2269 3066
rect 2274 3013 2277 3136
rect 2282 3076 2285 3126
rect 2314 3116 2317 3126
rect 2322 3123 2325 3136
rect 2354 3133 2357 3146
rect 2370 3133 2373 3156
rect 2378 3133 2381 3183
rect 2398 3176 2401 3233
rect 2434 3226 2437 3366
rect 2474 3346 2477 3406
rect 2482 3403 2493 3406
rect 2450 3323 2453 3346
rect 2474 3343 2485 3346
rect 2482 3323 2485 3343
rect 2490 3333 2493 3366
rect 2490 3313 2493 3326
rect 2498 3323 2501 3413
rect 2506 3333 2509 3346
rect 2514 3293 2517 3466
rect 2522 3423 2525 3436
rect 2530 3413 2533 3476
rect 2542 3426 2545 3483
rect 2538 3423 2545 3426
rect 2562 3423 2565 3523
rect 2614 3506 2617 3633
rect 2626 3613 2629 3653
rect 2626 3523 2629 3536
rect 2610 3503 2617 3506
rect 2538 3406 2541 3423
rect 2522 3393 2525 3406
rect 2530 3403 2541 3406
rect 2554 3393 2557 3416
rect 2562 3356 2565 3406
rect 2578 3393 2581 3426
rect 2522 3323 2525 3356
rect 2554 3353 2573 3356
rect 2530 3333 2549 3336
rect 2546 3283 2549 3326
rect 2554 3256 2557 3353
rect 2570 3333 2581 3336
rect 2570 3326 2573 3333
rect 2562 3323 2573 3326
rect 2538 3253 2557 3256
rect 2538 3236 2541 3253
rect 2394 3173 2401 3176
rect 2426 3223 2437 3226
rect 2534 3233 2541 3236
rect 2330 3116 2333 3126
rect 2314 3113 2333 3116
rect 2282 3073 2301 3076
rect 2290 3016 2293 3036
rect 2282 3013 2293 3016
rect 2274 2993 2277 3006
rect 2282 2986 2285 3013
rect 2258 2973 2269 2976
rect 2274 2983 2285 2986
rect 2186 2933 2189 2946
rect 2202 2943 2213 2946
rect 2130 2813 2133 2826
rect 2122 2793 2125 2806
rect 2114 2773 2125 2776
rect 2066 2733 2069 2756
rect 2074 2743 2077 2766
rect 2050 2643 2057 2646
rect 2050 2593 2053 2643
rect 2058 2583 2061 2606
rect 1994 2533 1997 2546
rect 2010 2476 2013 2553
rect 1986 2366 1989 2476
rect 2002 2453 2005 2476
rect 2010 2473 2021 2476
rect 1978 2363 1989 2366
rect 2002 2366 2005 2426
rect 2010 2416 2013 2446
rect 2018 2423 2021 2473
rect 2010 2413 2021 2416
rect 2026 2373 2029 2546
rect 2050 2403 2053 2496
rect 2058 2433 2061 2576
rect 2066 2486 2069 2716
rect 2082 2643 2085 2756
rect 2090 2613 2093 2726
rect 2098 2673 2101 2716
rect 2090 2596 2093 2606
rect 2074 2593 2093 2596
rect 2074 2513 2077 2526
rect 2090 2493 2093 2556
rect 2066 2483 2085 2486
rect 2082 2436 2085 2483
rect 2078 2433 2085 2436
rect 2002 2363 2013 2366
rect 1962 2333 1965 2346
rect 1950 2293 1957 2296
rect 1954 2226 1957 2293
rect 1962 2286 1965 2326
rect 1978 2306 1981 2363
rect 1978 2303 1985 2306
rect 1962 2283 1973 2286
rect 1950 2223 1957 2226
rect 1930 2003 1933 2216
rect 1938 2193 1941 2206
rect 1950 2146 1953 2223
rect 1962 2196 1965 2216
rect 1970 2203 1973 2283
rect 1982 2246 1985 2303
rect 1982 2243 1989 2246
rect 1978 2213 1981 2226
rect 1978 2196 1981 2206
rect 1962 2193 1981 2196
rect 1986 2186 1989 2243
rect 1970 2183 1989 2186
rect 1950 2143 1957 2146
rect 1946 2113 1949 2126
rect 1946 1946 1949 2016
rect 1954 1973 1957 2143
rect 1962 2076 1965 2166
rect 1970 2096 1973 2183
rect 1994 2133 1997 2256
rect 2010 2186 2013 2363
rect 2066 2356 2069 2406
rect 2078 2376 2081 2433
rect 2078 2373 2085 2376
rect 2066 2353 2077 2356
rect 2026 2213 2029 2326
rect 2050 2253 2053 2336
rect 2066 2323 2069 2346
rect 2002 2183 2013 2186
rect 2002 2163 2005 2183
rect 2018 2123 2021 2136
rect 2042 2123 2045 2216
rect 1970 2093 1981 2096
rect 1962 2073 1969 2076
rect 1966 2006 1969 2073
rect 1962 2003 1969 2006
rect 1962 1983 1965 2003
rect 1946 1943 1957 1946
rect 1922 1933 1949 1936
rect 1938 1896 1941 1916
rect 1930 1893 1941 1896
rect 1930 1836 1933 1893
rect 1930 1833 1941 1836
rect 1922 1803 1925 1816
rect 1914 1793 1925 1796
rect 1874 1623 1901 1626
rect 1862 1603 1869 1606
rect 1842 1563 1853 1566
rect 1842 1506 1845 1556
rect 1850 1516 1853 1563
rect 1858 1533 1861 1586
rect 1866 1533 1869 1603
rect 1874 1553 1877 1623
rect 1890 1603 1893 1616
rect 1898 1613 1901 1623
rect 1898 1596 1901 1606
rect 1906 1603 1909 1756
rect 1914 1723 1917 1776
rect 1922 1706 1925 1793
rect 1930 1743 1933 1816
rect 1938 1746 1941 1833
rect 1946 1763 1949 1933
rect 1954 1856 1957 1943
rect 1978 1926 1981 2093
rect 1962 1923 1981 1926
rect 1986 1903 1989 2026
rect 1994 1923 1997 2096
rect 2002 1916 2005 1976
rect 2010 1923 2021 1926
rect 2026 1923 2029 1946
rect 2002 1913 2013 1916
rect 2018 1913 2021 1923
rect 2034 1916 2037 2026
rect 2026 1913 2037 1916
rect 1954 1853 1973 1856
rect 1962 1803 1965 1816
rect 1938 1743 1945 1746
rect 1918 1703 1925 1706
rect 1918 1636 1921 1703
rect 1918 1633 1925 1636
rect 1914 1596 1917 1616
rect 1898 1593 1917 1596
rect 1882 1536 1885 1576
rect 1922 1543 1925 1633
rect 1930 1613 1933 1726
rect 1942 1646 1945 1743
rect 1938 1643 1945 1646
rect 1938 1623 1941 1643
rect 1938 1603 1941 1616
rect 1954 1603 1957 1716
rect 1962 1673 1965 1726
rect 1970 1693 1973 1853
rect 1978 1623 1981 1896
rect 1986 1743 1989 1876
rect 2002 1733 2005 1746
rect 1978 1603 1981 1616
rect 1986 1596 1989 1716
rect 2010 1713 2013 1913
rect 2026 1793 2029 1913
rect 2042 1906 2045 2116
rect 2034 1903 2045 1906
rect 2042 1893 2045 1903
rect 2050 1876 2053 2216
rect 2058 2086 2061 2246
rect 2066 2093 2069 2316
rect 2074 2213 2077 2353
rect 2082 2313 2085 2373
rect 2058 2083 2069 2086
rect 2066 2026 2069 2083
rect 2066 2023 2077 2026
rect 2058 1993 2061 2006
rect 2058 1913 2061 1926
rect 2046 1873 2053 1876
rect 2034 1746 2037 1846
rect 2046 1756 2049 1873
rect 2058 1843 2061 1906
rect 2066 1893 2069 1906
rect 2074 1886 2077 2023
rect 2082 2013 2085 2256
rect 2090 2096 2093 2426
rect 2098 2316 2101 2646
rect 2106 2603 2109 2766
rect 2122 2696 2125 2773
rect 2138 2763 2141 2816
rect 2114 2693 2125 2696
rect 2114 2673 2117 2693
rect 2114 2606 2117 2626
rect 2122 2613 2141 2616
rect 2114 2603 2125 2606
rect 2146 2583 2149 2796
rect 2154 2736 2157 2886
rect 2210 2883 2213 2943
rect 2218 2936 2221 2956
rect 2218 2933 2225 2936
rect 2222 2846 2225 2933
rect 2234 2893 2237 2926
rect 2258 2906 2261 2973
rect 2274 2933 2277 2983
rect 2274 2913 2277 2926
rect 2258 2903 2269 2906
rect 2218 2843 2225 2846
rect 2218 2823 2221 2843
rect 2170 2743 2173 2816
rect 2218 2786 2221 2816
rect 2242 2803 2245 2886
rect 2266 2846 2269 2903
rect 2266 2843 2273 2846
rect 2270 2796 2273 2843
rect 2266 2793 2273 2796
rect 2202 2756 2205 2786
rect 2218 2783 2229 2786
rect 2202 2753 2213 2756
rect 2154 2733 2169 2736
rect 2194 2733 2197 2746
rect 2154 2643 2157 2726
rect 2166 2646 2169 2733
rect 2166 2643 2173 2646
rect 2154 2613 2157 2636
rect 2162 2603 2165 2626
rect 2114 2533 2117 2576
rect 2106 2423 2109 2526
rect 2114 2416 2117 2526
rect 2122 2506 2125 2556
rect 2130 2543 2149 2546
rect 2130 2523 2133 2543
rect 2122 2503 2129 2506
rect 2126 2426 2129 2503
rect 2138 2493 2141 2536
rect 2146 2533 2149 2543
rect 2170 2533 2173 2643
rect 2178 2613 2181 2656
rect 2186 2606 2189 2676
rect 2202 2646 2205 2666
rect 2178 2603 2189 2606
rect 2198 2643 2205 2646
rect 2146 2473 2149 2526
rect 2154 2513 2157 2526
rect 2178 2516 2181 2603
rect 2198 2596 2201 2643
rect 2210 2603 2213 2753
rect 2226 2733 2229 2783
rect 2250 2703 2253 2766
rect 2218 2613 2237 2616
rect 2198 2593 2205 2596
rect 2202 2543 2205 2593
rect 2226 2576 2229 2613
rect 2218 2573 2229 2576
rect 2170 2513 2181 2516
rect 2106 2413 2117 2416
rect 2122 2423 2129 2426
rect 2106 2383 2109 2413
rect 2122 2406 2125 2423
rect 2138 2413 2141 2446
rect 2114 2336 2117 2406
rect 2122 2403 2133 2406
rect 2106 2333 2117 2336
rect 2098 2313 2105 2316
rect 2102 2236 2105 2313
rect 2114 2253 2117 2333
rect 2122 2316 2125 2386
rect 2130 2333 2133 2376
rect 2122 2313 2133 2316
rect 2130 2266 2133 2313
rect 2122 2263 2133 2266
rect 2122 2246 2125 2263
rect 2098 2233 2105 2236
rect 2114 2243 2125 2246
rect 2098 2113 2101 2233
rect 2106 2186 2109 2216
rect 2114 2213 2117 2243
rect 2114 2196 2117 2206
rect 2122 2203 2125 2216
rect 2130 2196 2133 2216
rect 2114 2193 2133 2196
rect 2106 2183 2117 2186
rect 2090 2093 2097 2096
rect 2094 2026 2097 2093
rect 2090 2023 2097 2026
rect 2106 2023 2109 2166
rect 2114 2133 2117 2183
rect 2122 2126 2125 2176
rect 2138 2163 2141 2206
rect 2138 2133 2141 2146
rect 2114 2123 2125 2126
rect 2114 2093 2117 2123
rect 2130 2113 2133 2126
rect 2090 2003 2093 2023
rect 2122 2016 2125 2036
rect 2114 2013 2125 2016
rect 2082 1923 2085 1946
rect 2090 1916 2093 1966
rect 2114 1933 2117 1976
rect 2122 1963 2125 2006
rect 2130 2003 2133 2016
rect 2138 2003 2141 2026
rect 2146 1936 2149 2466
rect 2154 2413 2157 2496
rect 2170 2456 2173 2513
rect 2186 2493 2189 2536
rect 2218 2533 2221 2573
rect 2218 2506 2221 2526
rect 2210 2503 2221 2506
rect 2162 2453 2173 2456
rect 2154 2156 2157 2226
rect 2162 2173 2165 2453
rect 2178 2426 2181 2446
rect 2174 2423 2181 2426
rect 2174 2196 2177 2423
rect 2186 2413 2189 2476
rect 2210 2446 2213 2503
rect 2210 2443 2221 2446
rect 2218 2423 2221 2443
rect 2186 2206 2189 2406
rect 2194 2333 2221 2336
rect 2202 2313 2205 2326
rect 2202 2213 2205 2246
rect 2186 2203 2205 2206
rect 2174 2193 2181 2196
rect 2154 2153 2165 2156
rect 2154 2113 2157 2136
rect 2162 2123 2165 2153
rect 2154 1983 2157 2026
rect 2146 1933 2153 1936
rect 2082 1913 2093 1916
rect 2098 1913 2101 1926
rect 2082 1896 2085 1913
rect 2082 1893 2093 1896
rect 2066 1883 2077 1886
rect 2046 1753 2053 1756
rect 2030 1743 2037 1746
rect 1994 1603 1997 1676
rect 1978 1593 1989 1596
rect 2002 1593 2005 1636
rect 1878 1533 1885 1536
rect 1850 1513 1857 1516
rect 1834 1503 1845 1506
rect 1834 1383 1837 1503
rect 1842 1423 1845 1496
rect 1854 1416 1857 1513
rect 1866 1493 1869 1516
rect 1878 1446 1881 1533
rect 1878 1443 1885 1446
rect 1850 1413 1857 1416
rect 1874 1413 1877 1426
rect 1818 1293 1821 1336
rect 1826 1233 1829 1366
rect 1850 1343 1853 1413
rect 1866 1366 1869 1406
rect 1874 1393 1877 1406
rect 1882 1403 1885 1443
rect 1890 1423 1893 1526
rect 1898 1503 1901 1526
rect 1906 1516 1909 1536
rect 1906 1513 1913 1516
rect 1858 1363 1869 1366
rect 1834 1313 1837 1326
rect 1842 1303 1845 1326
rect 1850 1276 1853 1336
rect 1858 1313 1861 1363
rect 1874 1336 1877 1356
rect 1866 1323 1869 1336
rect 1874 1333 1885 1336
rect 1874 1303 1877 1326
rect 1882 1313 1885 1333
rect 1842 1273 1853 1276
rect 1842 1213 1845 1273
rect 1818 1143 1821 1166
rect 1810 1123 1821 1126
rect 1786 1073 1797 1076
rect 1778 1013 1789 1016
rect 1794 1006 1797 1073
rect 1714 933 1721 936
rect 1690 913 1701 916
rect 1698 896 1701 913
rect 1698 893 1705 896
rect 1682 813 1685 826
rect 1690 813 1693 866
rect 1702 836 1705 893
rect 1718 846 1721 933
rect 1718 843 1725 846
rect 1698 833 1705 836
rect 1626 703 1629 723
rect 1642 683 1645 726
rect 1610 613 1613 656
rect 1650 636 1653 756
rect 1666 753 1685 756
rect 1690 753 1693 806
rect 1698 803 1701 833
rect 1706 803 1709 816
rect 1714 803 1717 826
rect 1722 816 1725 843
rect 1730 823 1733 936
rect 1722 813 1733 816
rect 1682 746 1685 753
rect 1658 743 1677 746
rect 1682 743 1689 746
rect 1658 723 1661 743
rect 1666 723 1669 736
rect 1674 733 1677 743
rect 1642 633 1653 636
rect 1626 613 1629 626
rect 1586 563 1597 566
rect 1570 553 1581 556
rect 1554 523 1565 526
rect 1538 473 1541 523
rect 1554 506 1557 523
rect 1570 516 1573 536
rect 1578 523 1581 553
rect 1550 503 1557 506
rect 1562 513 1573 516
rect 1550 436 1553 503
rect 1498 403 1501 416
rect 1530 413 1533 436
rect 1550 433 1557 436
rect 1554 416 1557 433
rect 1538 403 1541 416
rect 1546 413 1557 416
rect 1434 363 1453 366
rect 1434 306 1437 363
rect 1546 356 1549 413
rect 1554 396 1557 406
rect 1562 403 1565 513
rect 1570 396 1573 416
rect 1554 393 1573 396
rect 1578 356 1581 476
rect 1586 453 1589 536
rect 1594 523 1597 563
rect 1602 543 1605 606
rect 1618 563 1621 606
rect 1634 593 1637 606
rect 1602 523 1613 526
rect 1586 413 1589 426
rect 1594 396 1597 516
rect 1618 473 1621 536
rect 1602 403 1605 426
rect 1610 403 1613 416
rect 1618 413 1621 436
rect 1618 396 1621 406
rect 1594 393 1621 396
rect 1538 353 1549 356
rect 1570 353 1581 356
rect 1482 313 1485 326
rect 1514 323 1517 346
rect 1522 313 1525 326
rect 1426 303 1437 306
rect 1426 236 1429 303
rect 1422 233 1429 236
rect 1274 133 1277 206
rect 1282 203 1293 206
rect 1306 186 1309 206
rect 1410 193 1413 206
rect 1422 186 1425 233
rect 1434 203 1437 216
rect 1290 183 1309 186
rect 1418 183 1425 186
rect 1250 123 1269 126
rect 1290 123 1293 183
rect 1314 123 1317 136
rect 1394 123 1397 156
rect 1418 123 1421 183
rect 1442 123 1445 216
rect 1450 103 1453 216
rect 1458 196 1461 206
rect 1466 203 1469 236
rect 1474 196 1477 216
rect 1458 193 1477 196
rect 1482 193 1485 306
rect 1530 213 1533 326
rect 1538 323 1541 353
rect 1546 343 1565 346
rect 1546 333 1549 343
rect 1554 323 1557 336
rect 1562 323 1565 343
rect 1498 123 1501 206
rect 1514 123 1517 136
rect 1538 123 1541 216
rect 1546 213 1549 316
rect 1570 236 1573 353
rect 1578 333 1581 346
rect 1602 333 1605 366
rect 1618 333 1621 393
rect 1626 326 1629 576
rect 1634 503 1637 526
rect 1642 513 1645 633
rect 1650 613 1653 626
rect 1658 533 1661 616
rect 1666 573 1669 706
rect 1666 526 1669 536
rect 1650 523 1669 526
rect 1674 506 1677 726
rect 1686 676 1689 743
rect 1698 686 1701 776
rect 1722 743 1725 806
rect 1706 703 1709 726
rect 1714 723 1725 726
rect 1730 693 1733 813
rect 1738 803 1741 936
rect 1746 903 1749 1006
rect 1754 966 1757 1006
rect 1762 983 1765 1006
rect 1786 1003 1797 1006
rect 1754 963 1765 966
rect 1754 933 1757 956
rect 1762 926 1765 963
rect 1770 953 1773 976
rect 1754 923 1765 926
rect 1754 833 1757 923
rect 1778 913 1781 936
rect 1762 813 1765 906
rect 1754 783 1757 806
rect 1770 803 1773 826
rect 1786 823 1789 976
rect 1794 863 1797 986
rect 1802 933 1805 1086
rect 1818 1066 1821 1123
rect 1810 1063 1821 1066
rect 1810 973 1813 1063
rect 1826 1013 1829 1036
rect 1802 903 1805 926
rect 1810 923 1821 926
rect 1810 853 1813 923
rect 1826 913 1829 926
rect 1786 786 1789 816
rect 1762 783 1789 786
rect 1746 703 1749 726
rect 1698 683 1709 686
rect 1686 673 1693 676
rect 1690 566 1693 673
rect 1686 563 1693 566
rect 1686 516 1689 563
rect 1698 523 1701 616
rect 1686 513 1693 516
rect 1666 503 1677 506
rect 1642 426 1645 476
rect 1666 446 1669 503
rect 1666 443 1677 446
rect 1634 413 1637 426
rect 1642 423 1661 426
rect 1642 403 1645 423
rect 1658 413 1661 423
rect 1674 406 1677 443
rect 1690 433 1693 513
rect 1706 506 1709 683
rect 1702 503 1709 506
rect 1650 403 1677 406
rect 1690 403 1693 416
rect 1578 293 1581 326
rect 1586 266 1589 326
rect 1610 323 1629 326
rect 1562 233 1573 236
rect 1578 263 1597 266
rect 1554 196 1557 206
rect 1562 203 1565 233
rect 1578 223 1581 263
rect 1570 196 1573 216
rect 1586 213 1589 256
rect 1594 213 1597 263
rect 1554 193 1573 196
rect 1578 126 1581 206
rect 1586 193 1589 206
rect 1578 123 1597 126
rect 1602 43 1605 236
rect 1610 216 1613 323
rect 1634 306 1637 356
rect 1650 336 1653 403
rect 1702 356 1705 503
rect 1714 376 1717 616
rect 1738 573 1741 606
rect 1722 533 1725 556
rect 1738 533 1741 546
rect 1762 536 1765 783
rect 1762 533 1773 536
rect 1722 513 1725 526
rect 1738 403 1741 526
rect 1762 513 1765 526
rect 1770 506 1773 533
rect 1778 523 1781 576
rect 1794 573 1797 736
rect 1802 613 1805 656
rect 1810 596 1813 826
rect 1818 813 1821 906
rect 1834 883 1837 1116
rect 1842 1113 1845 1136
rect 1826 773 1829 866
rect 1842 853 1845 1016
rect 1826 743 1845 746
rect 1826 733 1829 743
rect 1818 653 1821 726
rect 1826 683 1829 726
rect 1806 593 1813 596
rect 1806 516 1809 593
rect 1818 523 1821 546
rect 1806 513 1813 516
rect 1762 503 1773 506
rect 1762 376 1765 503
rect 1714 373 1733 376
rect 1762 373 1773 376
rect 1682 353 1705 356
rect 1626 303 1637 306
rect 1642 333 1653 336
rect 1626 236 1629 303
rect 1626 233 1637 236
rect 1610 213 1629 216
rect 1610 163 1613 213
rect 1618 173 1621 206
rect 1618 113 1621 156
rect 1626 133 1629 166
rect 1634 133 1637 233
rect 1642 213 1645 333
rect 1650 313 1653 326
rect 1634 113 1637 126
rect 1642 123 1645 206
rect 1658 163 1661 216
rect 1666 193 1669 336
rect 1682 293 1685 353
rect 1682 213 1685 236
rect 1674 113 1677 126
rect 1682 103 1685 206
rect 1690 203 1693 316
rect 1698 213 1701 346
rect 1706 313 1709 326
rect 1706 193 1709 216
rect 1714 213 1717 296
rect 1730 276 1733 373
rect 1746 333 1749 346
rect 1770 333 1773 373
rect 1746 313 1749 326
rect 1726 273 1733 276
rect 1714 183 1717 206
rect 1726 166 1729 273
rect 1738 213 1741 276
rect 1754 273 1757 296
rect 1794 293 1797 436
rect 1802 413 1805 426
rect 1722 163 1729 166
rect 1722 103 1725 163
rect 1738 123 1741 196
rect 1746 23 1749 256
rect 1762 213 1765 266
rect 1778 213 1781 256
rect 1754 173 1757 206
rect 1770 193 1773 206
rect 1786 133 1789 266
rect 1802 256 1805 326
rect 1810 263 1813 513
rect 1826 503 1829 526
rect 1834 426 1837 736
rect 1842 723 1845 743
rect 1850 706 1853 1236
rect 1890 1233 1893 1406
rect 1898 1353 1901 1486
rect 1910 1446 1913 1513
rect 1906 1443 1913 1446
rect 1906 1396 1909 1443
rect 1914 1403 1917 1426
rect 1922 1413 1925 1536
rect 1930 1533 1949 1536
rect 1954 1493 1957 1526
rect 1962 1446 1965 1546
rect 1978 1533 1981 1593
rect 1994 1473 1997 1526
rect 2002 1516 2005 1536
rect 2002 1513 2009 1516
rect 1962 1443 1969 1446
rect 1906 1393 1917 1396
rect 1906 1276 1909 1336
rect 1914 1326 1917 1393
rect 1938 1346 1941 1406
rect 1966 1396 1969 1443
rect 1962 1393 1969 1396
rect 1938 1343 1949 1346
rect 1922 1333 1941 1336
rect 1914 1323 1933 1326
rect 1938 1323 1941 1333
rect 1930 1296 1933 1316
rect 1930 1293 1937 1296
rect 1906 1273 1925 1276
rect 1922 1213 1925 1273
rect 1858 1133 1861 1196
rect 1874 1193 1877 1206
rect 1898 1193 1901 1206
rect 1898 1146 1901 1166
rect 1890 1143 1901 1146
rect 1858 1113 1861 1126
rect 1890 1046 1893 1143
rect 1922 1133 1925 1196
rect 1934 1186 1937 1293
rect 1946 1193 1949 1343
rect 1954 1303 1957 1326
rect 1962 1256 1965 1393
rect 1970 1316 1973 1336
rect 1978 1333 1981 1406
rect 1986 1393 1989 1416
rect 2006 1376 2009 1513
rect 2002 1373 2009 1376
rect 1970 1313 1981 1316
rect 1962 1253 1969 1256
rect 1966 1196 1969 1253
rect 1978 1213 1981 1313
rect 1962 1193 1969 1196
rect 1930 1183 1937 1186
rect 1930 1163 1933 1183
rect 1962 1176 1965 1193
rect 1954 1173 1965 1176
rect 1890 1043 1897 1046
rect 1858 906 1861 936
rect 1858 903 1869 906
rect 1846 703 1853 706
rect 1846 576 1849 703
rect 1846 573 1853 576
rect 1842 523 1845 556
rect 1830 423 1837 426
rect 1830 376 1833 423
rect 1842 393 1845 416
rect 1830 373 1837 376
rect 1834 343 1837 373
rect 1850 336 1853 573
rect 1858 566 1861 856
rect 1866 743 1869 903
rect 1874 813 1877 1006
rect 1894 956 1897 1043
rect 1894 953 1901 956
rect 1874 783 1877 796
rect 1866 706 1869 736
rect 1874 723 1877 776
rect 1866 703 1873 706
rect 1870 636 1873 703
rect 1882 693 1885 846
rect 1898 823 1901 953
rect 1906 923 1909 1106
rect 1954 1023 1957 1173
rect 1970 1123 1973 1136
rect 1986 1113 1989 1346
rect 1994 1133 1997 1336
rect 2002 1213 2005 1373
rect 2010 1323 2013 1336
rect 2018 1226 2021 1696
rect 2030 1686 2033 1743
rect 2042 1693 2045 1736
rect 2030 1683 2037 1686
rect 2034 1626 2037 1683
rect 2034 1623 2045 1626
rect 2026 1613 2037 1616
rect 2026 1323 2029 1596
rect 2034 1506 2037 1536
rect 2042 1523 2045 1623
rect 2034 1503 2041 1506
rect 2038 1446 2041 1503
rect 2034 1443 2041 1446
rect 2034 1373 2037 1443
rect 2050 1403 2053 1753
rect 2058 1743 2061 1816
rect 2066 1796 2069 1883
rect 2074 1803 2077 1846
rect 2090 1826 2093 1893
rect 2082 1823 2093 1826
rect 2066 1793 2077 1796
rect 2066 1733 2069 1756
rect 2074 1726 2077 1793
rect 2082 1786 2085 1823
rect 2106 1813 2109 1906
rect 2114 1853 2117 1926
rect 2138 1903 2141 1926
rect 2150 1876 2153 1933
rect 2146 1873 2153 1876
rect 2114 1813 2125 1816
rect 2090 1793 2093 1806
rect 2082 1783 2093 1786
rect 2090 1736 2093 1783
rect 2090 1733 2097 1736
rect 2058 1673 2061 1726
rect 2066 1723 2077 1726
rect 2066 1633 2069 1723
rect 2082 1713 2085 1726
rect 2074 1616 2077 1626
rect 2058 1603 2061 1616
rect 2066 1613 2077 1616
rect 2066 1533 2069 1613
rect 2082 1603 2085 1676
rect 2094 1656 2097 1733
rect 2106 1723 2109 1776
rect 2114 1753 2117 1806
rect 2122 1756 2125 1813
rect 2130 1793 2133 1816
rect 2122 1753 2133 1756
rect 2090 1653 2097 1656
rect 2090 1593 2093 1653
rect 2058 1493 2061 1516
rect 2066 1503 2069 1526
rect 2082 1396 2085 1536
rect 2090 1403 2093 1416
rect 2042 1366 2045 1386
rect 2034 1363 2045 1366
rect 2010 1223 2021 1226
rect 2002 1106 2005 1126
rect 1998 1103 2005 1106
rect 1998 1046 2001 1103
rect 2010 1083 2013 1223
rect 2034 1216 2037 1363
rect 2050 1333 2053 1346
rect 2034 1213 2041 1216
rect 2018 1106 2021 1176
rect 2026 1123 2029 1206
rect 2038 1136 2041 1213
rect 2034 1133 2041 1136
rect 2018 1103 2025 1106
rect 2022 1046 2025 1103
rect 1998 1043 2005 1046
rect 2022 1043 2029 1046
rect 1914 923 1917 1016
rect 1922 913 1925 1016
rect 1946 933 1949 1006
rect 1986 973 1989 1006
rect 2002 983 2005 1043
rect 2026 996 2029 1043
rect 2018 993 2029 996
rect 1970 943 1997 946
rect 1970 936 1973 943
rect 1954 933 1973 936
rect 1890 793 1893 806
rect 1890 733 1893 746
rect 1898 723 1901 796
rect 1906 786 1909 816
rect 1914 803 1917 816
rect 1922 803 1925 846
rect 1930 803 1933 886
rect 1938 813 1941 926
rect 1954 923 1957 933
rect 1946 806 1949 916
rect 1962 903 1965 926
rect 1978 923 1981 936
rect 1986 863 1989 936
rect 1994 933 1997 943
rect 1994 856 1997 926
rect 2002 913 2005 966
rect 1978 853 1997 856
rect 1978 833 1981 853
rect 1938 803 1949 806
rect 1906 783 1917 786
rect 1914 733 1917 783
rect 1866 633 1873 636
rect 1866 613 1869 633
rect 1858 563 1869 566
rect 1858 533 1861 546
rect 1866 433 1869 563
rect 1858 413 1861 426
rect 1874 413 1877 616
rect 1906 613 1909 626
rect 1938 623 1941 803
rect 1954 796 1957 826
rect 1946 793 1957 796
rect 1946 683 1949 793
rect 1962 756 1965 816
rect 1970 803 1973 826
rect 1986 783 1989 806
rect 2010 793 2013 926
rect 2018 776 2021 993
rect 2026 923 2029 936
rect 2034 933 2037 1133
rect 2042 1003 2045 1116
rect 2050 1093 2053 1326
rect 2058 1323 2061 1376
rect 2066 1333 2069 1396
rect 2082 1393 2093 1396
rect 2074 1213 2077 1326
rect 2082 1313 2085 1356
rect 2058 1056 2061 1206
rect 2082 1203 2085 1226
rect 2090 1213 2093 1393
rect 2098 1186 2101 1636
rect 2114 1616 2117 1746
rect 2122 1733 2125 1746
rect 2130 1743 2133 1753
rect 2130 1713 2133 1736
rect 2138 1696 2141 1856
rect 2130 1693 2141 1696
rect 2130 1636 2133 1693
rect 2106 1613 2117 1616
rect 2122 1633 2133 1636
rect 2106 1473 2109 1613
rect 2114 1533 2117 1606
rect 2114 1493 2117 1516
rect 2122 1476 2125 1633
rect 2130 1533 2133 1626
rect 2118 1473 2125 1476
rect 2118 1376 2121 1473
rect 2090 1183 2101 1186
rect 2106 1373 2121 1376
rect 2090 1126 2093 1183
rect 2106 1133 2109 1373
rect 2114 1203 2117 1346
rect 2122 1253 2125 1366
rect 2130 1243 2133 1526
rect 2138 1333 2141 1406
rect 2146 1373 2149 1873
rect 2162 1866 2165 2096
rect 2170 2003 2173 2146
rect 2178 2023 2181 2193
rect 2186 2113 2189 2126
rect 2194 2123 2197 2146
rect 2178 2003 2181 2016
rect 2194 2013 2197 2036
rect 2162 1863 2169 1866
rect 2154 1833 2157 1856
rect 2154 1773 2157 1816
rect 2166 1776 2169 1863
rect 2162 1773 2169 1776
rect 2162 1753 2165 1773
rect 2162 1726 2165 1746
rect 2178 1743 2181 1986
rect 2186 1946 2189 2006
rect 2202 2003 2205 2203
rect 2210 2003 2213 2326
rect 2218 2213 2221 2333
rect 2226 2286 2229 2546
rect 2234 2513 2237 2586
rect 2242 2573 2245 2676
rect 2266 2673 2269 2793
rect 2282 2766 2285 2966
rect 2290 2933 2293 3006
rect 2298 3003 2301 3073
rect 2306 2976 2309 3026
rect 2322 3023 2341 3026
rect 2322 3003 2325 3023
rect 2330 3003 2333 3016
rect 2338 3013 2341 3023
rect 2346 3013 2357 3016
rect 2338 3003 2349 3006
rect 2298 2973 2309 2976
rect 2298 2916 2301 2973
rect 2306 2933 2317 2936
rect 2330 2933 2333 2966
rect 2338 2933 2341 2986
rect 2354 2983 2357 3006
rect 2362 2976 2365 3126
rect 2378 3113 2381 3126
rect 2386 3103 2389 3126
rect 2370 2993 2373 3006
rect 2354 2973 2365 2976
rect 2306 2923 2317 2926
rect 2322 2916 2325 2926
rect 2346 2923 2349 2946
rect 2354 2926 2357 2973
rect 2386 2963 2389 3026
rect 2394 2973 2397 3173
rect 2410 3133 2413 3156
rect 2426 3146 2429 3223
rect 2426 3143 2437 3146
rect 2402 3023 2405 3126
rect 2410 3013 2413 3026
rect 2418 3013 2421 3126
rect 2362 2933 2365 2946
rect 2354 2923 2365 2926
rect 2370 2923 2373 2956
rect 2402 2953 2405 3006
rect 2290 2903 2293 2916
rect 2298 2913 2325 2916
rect 2330 2896 2333 2916
rect 2362 2913 2365 2923
rect 2322 2893 2333 2896
rect 2322 2836 2325 2893
rect 2322 2833 2333 2836
rect 2290 2803 2293 2816
rect 2282 2763 2293 2766
rect 2290 2746 2293 2763
rect 2290 2743 2297 2746
rect 2274 2646 2277 2696
rect 2294 2686 2297 2743
rect 2266 2643 2277 2646
rect 2290 2683 2297 2686
rect 2250 2456 2253 2616
rect 2258 2603 2261 2626
rect 2258 2523 2261 2536
rect 2242 2453 2253 2456
rect 2242 2436 2245 2453
rect 2238 2433 2245 2436
rect 2238 2376 2241 2433
rect 2258 2413 2261 2426
rect 2238 2373 2245 2376
rect 2242 2296 2245 2373
rect 2250 2313 2253 2326
rect 2242 2293 2249 2296
rect 2226 2283 2237 2286
rect 2226 2203 2229 2216
rect 2234 2133 2237 2283
rect 2246 2226 2249 2293
rect 2242 2223 2249 2226
rect 2226 2113 2229 2126
rect 2234 2016 2237 2036
rect 2242 2023 2245 2223
rect 2226 2003 2229 2016
rect 2234 2013 2245 2016
rect 2234 1983 2237 2006
rect 2242 1976 2245 2006
rect 2234 1973 2245 1976
rect 2186 1943 2205 1946
rect 2194 1836 2197 1926
rect 2210 1873 2213 1936
rect 2186 1833 2197 1836
rect 2186 1803 2189 1833
rect 2202 1826 2205 1836
rect 2194 1823 2205 1826
rect 2194 1736 2197 1823
rect 2194 1733 2205 1736
rect 2154 1713 2157 1726
rect 2162 1723 2181 1726
rect 2178 1706 2181 1723
rect 2194 1713 2197 1726
rect 2170 1703 2181 1706
rect 2170 1636 2173 1703
rect 2202 1656 2205 1733
rect 2186 1653 2205 1656
rect 2210 1656 2213 1826
rect 2218 1803 2221 1926
rect 2226 1746 2229 1926
rect 2234 1773 2237 1973
rect 2250 1933 2253 2206
rect 2258 2203 2261 2406
rect 2266 2286 2269 2643
rect 2274 2533 2277 2636
rect 2290 2626 2293 2683
rect 2282 2623 2293 2626
rect 2274 2403 2277 2526
rect 2282 2376 2285 2623
rect 2290 2443 2293 2616
rect 2298 2603 2301 2616
rect 2306 2606 2309 2826
rect 2322 2776 2325 2816
rect 2330 2813 2333 2833
rect 2338 2813 2341 2896
rect 2346 2823 2349 2906
rect 2370 2903 2373 2916
rect 2386 2913 2389 2926
rect 2394 2896 2397 2936
rect 2402 2923 2405 2946
rect 2370 2893 2397 2896
rect 2370 2813 2373 2893
rect 2410 2876 2413 2936
rect 2418 2933 2421 3006
rect 2426 2983 2429 3106
rect 2434 2956 2437 3143
rect 2442 3133 2445 3216
rect 2466 3193 2469 3206
rect 2490 3193 2493 3206
rect 2514 3166 2517 3216
rect 2498 3163 2517 3166
rect 2442 2963 2445 3126
rect 2458 3036 2461 3056
rect 2458 3033 2465 3036
rect 2462 2976 2465 3033
rect 2458 2973 2465 2976
rect 2426 2933 2429 2956
rect 2434 2953 2453 2956
rect 2402 2873 2413 2876
rect 2386 2823 2389 2836
rect 2402 2823 2405 2873
rect 2418 2866 2421 2926
rect 2410 2863 2421 2866
rect 2378 2806 2381 2816
rect 2330 2803 2349 2806
rect 2370 2803 2381 2806
rect 2322 2773 2341 2776
rect 2314 2693 2317 2736
rect 2322 2696 2325 2746
rect 2338 2733 2341 2773
rect 2330 2713 2341 2716
rect 2322 2693 2333 2696
rect 2338 2693 2341 2713
rect 2346 2703 2349 2726
rect 2330 2616 2333 2693
rect 2354 2686 2357 2776
rect 2370 2713 2373 2803
rect 2394 2733 2397 2806
rect 2402 2786 2405 2816
rect 2410 2813 2413 2863
rect 2434 2836 2437 2926
rect 2442 2923 2445 2936
rect 2450 2856 2453 2953
rect 2458 2923 2461 2973
rect 2474 2856 2477 3126
rect 2498 3123 2501 3163
rect 2522 3133 2525 3196
rect 2534 3176 2537 3233
rect 2570 3213 2573 3323
rect 2578 3313 2581 3326
rect 2586 3323 2589 3416
rect 2594 3403 2597 3416
rect 2594 3333 2597 3356
rect 2594 3313 2597 3326
rect 2602 3283 2605 3476
rect 2610 3463 2613 3503
rect 2626 3486 2629 3516
rect 2634 3496 2637 3716
rect 2642 3623 2645 3656
rect 2658 3643 2661 3893
rect 2666 3833 2677 3836
rect 2666 3783 2669 3833
rect 2706 3826 2709 3923
rect 2730 3906 2733 3926
rect 2722 3903 2733 3906
rect 2722 3836 2725 3903
rect 2738 3843 2741 3956
rect 2722 3833 2733 3836
rect 2698 3823 2709 3826
rect 2674 3793 2677 3816
rect 2666 3686 2669 3736
rect 2674 3703 2677 3726
rect 2666 3683 2673 3686
rect 2642 3563 2645 3616
rect 2642 3503 2645 3536
rect 2634 3493 2641 3496
rect 2618 3483 2629 3486
rect 2618 3446 2621 3483
rect 2610 3443 2621 3446
rect 2610 3373 2613 3443
rect 2618 3423 2621 3436
rect 2626 3413 2629 3476
rect 2638 3436 2641 3493
rect 2650 3443 2653 3596
rect 2658 3593 2661 3606
rect 2658 3473 2661 3586
rect 2670 3566 2673 3683
rect 2682 3583 2685 3776
rect 2690 3713 2693 3816
rect 2698 3726 2701 3823
rect 2706 3733 2709 3816
rect 2714 3733 2717 3816
rect 2722 3783 2725 3806
rect 2722 3736 2725 3766
rect 2730 3743 2733 3833
rect 2746 3813 2749 3826
rect 2754 3813 2757 3973
rect 2762 3933 2765 3946
rect 2778 3933 2781 3946
rect 2786 3933 2789 3966
rect 2802 3933 2805 3996
rect 2834 3993 2837 4016
rect 2850 4013 2853 4026
rect 2946 4023 2949 4140
rect 2826 3933 2829 3976
rect 2770 3823 2773 3926
rect 2786 3903 2789 3926
rect 2810 3913 2813 3926
rect 2834 3923 2837 3936
rect 2842 3933 2845 4006
rect 2882 4003 2885 4016
rect 2930 4003 2933 4016
rect 2738 3793 2741 3806
rect 2754 3773 2757 3806
rect 2722 3733 2733 3736
rect 2698 3723 2709 3726
rect 2730 3723 2733 3733
rect 2698 3616 2701 3626
rect 2690 3613 2701 3616
rect 2690 3593 2693 3606
rect 2666 3563 2673 3566
rect 2666 3533 2669 3563
rect 2706 3546 2709 3723
rect 2714 3573 2717 3606
rect 2722 3576 2725 3616
rect 2730 3613 2733 3626
rect 2738 3613 2741 3736
rect 2754 3733 2757 3746
rect 2746 3693 2749 3726
rect 2762 3626 2765 3806
rect 2770 3773 2773 3816
rect 2786 3803 2789 3866
rect 2850 3856 2853 3996
rect 2858 3916 2861 3966
rect 2866 3933 2869 3956
rect 2858 3913 2869 3916
rect 2850 3853 2857 3856
rect 2834 3813 2837 3826
rect 2854 3796 2857 3853
rect 2850 3793 2857 3796
rect 2850 3776 2853 3793
rect 2834 3773 2853 3776
rect 2786 3733 2789 3756
rect 2754 3623 2765 3626
rect 2730 3593 2733 3606
rect 2722 3573 2729 3576
rect 2674 3543 2701 3546
rect 2706 3543 2717 3546
rect 2674 3533 2677 3543
rect 2666 3523 2677 3526
rect 2682 3516 2685 3526
rect 2674 3513 2685 3516
rect 2690 3513 2693 3536
rect 2698 3533 2701 3543
rect 2706 3523 2709 3536
rect 2714 3513 2717 3543
rect 2682 3483 2685 3513
rect 2726 3486 2729 3573
rect 2738 3513 2741 3586
rect 2754 3576 2757 3623
rect 2762 3603 2765 3616
rect 2770 3593 2773 3656
rect 2794 3653 2797 3726
rect 2778 3623 2781 3646
rect 2778 3603 2781 3616
rect 2802 3613 2805 3736
rect 2810 3663 2813 3766
rect 2826 3733 2829 3746
rect 2746 3573 2757 3576
rect 2746 3496 2749 3573
rect 2754 3523 2757 3566
rect 2722 3483 2729 3486
rect 2738 3493 2749 3496
rect 2722 3463 2725 3483
rect 2738 3436 2741 3493
rect 2638 3433 2645 3436
rect 2618 3313 2621 3396
rect 2626 3353 2629 3406
rect 2634 3323 2637 3416
rect 2642 3316 2645 3433
rect 2650 3356 2653 3436
rect 2658 3363 2661 3426
rect 2666 3393 2669 3426
rect 2722 3423 2725 3436
rect 2738 3433 2749 3436
rect 2690 3396 2693 3406
rect 2698 3403 2701 3416
rect 2690 3393 2701 3396
rect 2706 3393 2709 3416
rect 2722 3396 2725 3416
rect 2746 3413 2749 3433
rect 2754 3406 2757 3516
rect 2762 3423 2765 3536
rect 2778 3513 2781 3576
rect 2786 3533 2789 3556
rect 2802 3533 2805 3606
rect 2810 3603 2813 3636
rect 2818 3596 2821 3626
rect 2810 3593 2821 3596
rect 2810 3526 2813 3593
rect 2794 3473 2797 3526
rect 2810 3523 2821 3526
rect 2826 3453 2829 3686
rect 2834 3533 2837 3773
rect 2842 3733 2845 3766
rect 2866 3756 2869 3913
rect 2850 3733 2853 3756
rect 2858 3753 2869 3756
rect 2882 3753 2885 3926
rect 2890 3883 2893 3936
rect 2906 3916 2909 3936
rect 2902 3913 2909 3916
rect 2902 3846 2905 3913
rect 2914 3856 2917 3936
rect 2922 3933 2925 3946
rect 2930 3933 2933 3966
rect 2938 3866 2941 3926
rect 2962 3923 2965 4016
rect 2978 4013 2981 4026
rect 2970 3933 2973 4006
rect 3026 4003 3029 4016
rect 3074 4003 3077 4016
rect 2986 3933 2989 3976
rect 2978 3913 2981 3926
rect 2938 3863 2945 3866
rect 2914 3853 2933 3856
rect 2902 3843 2909 3846
rect 2906 3823 2909 3843
rect 2890 3763 2893 3816
rect 2922 3776 2925 3816
rect 2898 3753 2901 3776
rect 2906 3773 2925 3776
rect 2842 3713 2845 3726
rect 2858 3696 2861 3753
rect 2850 3693 2861 3696
rect 2850 3636 2853 3693
rect 2842 3633 2853 3636
rect 2842 3583 2845 3633
rect 2850 3613 2853 3626
rect 2718 3393 2725 3396
rect 2650 3353 2661 3356
rect 2650 3333 2653 3346
rect 2634 3313 2645 3316
rect 2534 3173 2541 3176
rect 2586 3173 2589 3206
rect 2634 3203 2637 3313
rect 2658 3303 2661 3353
rect 2666 3286 2669 3336
rect 2674 3333 2677 3356
rect 2658 3283 2669 3286
rect 2658 3236 2661 3283
rect 2658 3233 2669 3236
rect 2538 3123 2541 3173
rect 2578 3123 2581 3136
rect 2482 3003 2485 3016
rect 2530 3013 2541 3016
rect 2578 3013 2581 3036
rect 2506 2986 2509 3006
rect 2586 2996 2589 3126
rect 2626 3106 2629 3176
rect 2666 3143 2669 3233
rect 2674 3223 2677 3316
rect 2690 3213 2693 3326
rect 2698 3323 2701 3393
rect 2706 3236 2709 3366
rect 2718 3336 2721 3393
rect 2718 3333 2725 3336
rect 2722 3316 2725 3333
rect 2730 3323 2733 3396
rect 2738 3383 2741 3406
rect 2746 3403 2757 3406
rect 2746 3333 2749 3403
rect 2754 3333 2757 3366
rect 2722 3313 2733 3316
rect 2698 3233 2709 3236
rect 2674 3186 2677 3206
rect 2698 3203 2701 3233
rect 2730 3213 2733 3313
rect 2754 3303 2757 3316
rect 2762 3246 2765 3416
rect 2770 3413 2773 3446
rect 2802 3343 2805 3436
rect 2770 3313 2773 3326
rect 2778 3313 2781 3336
rect 2810 3333 2813 3366
rect 2818 3323 2821 3446
rect 2842 3436 2845 3556
rect 2858 3533 2861 3616
rect 2866 3613 2869 3736
rect 2882 3726 2885 3746
rect 2898 3736 2901 3746
rect 2890 3733 2901 3736
rect 2906 3733 2909 3773
rect 2930 3766 2933 3853
rect 2942 3766 2945 3863
rect 2986 3813 2989 3826
rect 2970 3776 2973 3806
rect 2994 3803 2997 3926
rect 3002 3793 3005 3946
rect 2978 3776 2981 3786
rect 2970 3773 2981 3776
rect 2914 3763 2933 3766
rect 2938 3763 2945 3766
rect 2874 3673 2877 3726
rect 2882 3723 2893 3726
rect 2898 3693 2901 3733
rect 2866 3533 2869 3606
rect 2890 3573 2893 3626
rect 2882 3533 2885 3556
rect 2890 3533 2893 3566
rect 2842 3433 2853 3436
rect 2834 3376 2837 3416
rect 2826 3373 2837 3376
rect 2826 3333 2829 3373
rect 2842 3333 2845 3346
rect 2802 3303 2805 3316
rect 2758 3243 2765 3246
rect 2674 3183 2685 3186
rect 2682 3136 2685 3183
rect 2674 3133 2685 3136
rect 2626 3103 2637 3106
rect 2582 2993 2589 2996
rect 2506 2983 2525 2986
rect 2450 2853 2461 2856
rect 2434 2833 2453 2836
rect 2426 2823 2445 2826
rect 2410 2796 2413 2806
rect 2418 2803 2421 2816
rect 2426 2796 2429 2823
rect 2434 2803 2437 2816
rect 2442 2813 2445 2823
rect 2450 2808 2453 2833
rect 2442 2805 2453 2808
rect 2458 2796 2461 2853
rect 2410 2793 2429 2796
rect 2450 2793 2461 2796
rect 2466 2853 2477 2856
rect 2402 2783 2413 2786
rect 2354 2683 2365 2686
rect 2330 2613 2349 2616
rect 2354 2613 2357 2626
rect 2362 2616 2365 2683
rect 2386 2636 2389 2706
rect 2410 2703 2413 2783
rect 2450 2776 2453 2793
rect 2446 2773 2453 2776
rect 2418 2713 2421 2726
rect 2426 2703 2429 2716
rect 2434 2673 2437 2726
rect 2446 2686 2449 2773
rect 2446 2683 2453 2686
rect 2450 2656 2453 2683
rect 2450 2653 2457 2656
rect 2386 2633 2413 2636
rect 2362 2613 2373 2616
rect 2378 2613 2381 2626
rect 2306 2603 2333 2606
rect 2298 2513 2301 2526
rect 2306 2405 2309 2566
rect 2314 2533 2325 2536
rect 2322 2386 2325 2526
rect 2330 2493 2333 2603
rect 2338 2583 2341 2606
rect 2362 2586 2365 2606
rect 2354 2583 2365 2586
rect 2338 2523 2341 2536
rect 2354 2526 2357 2583
rect 2370 2566 2373 2613
rect 2386 2583 2389 2633
rect 2394 2603 2397 2626
rect 2410 2613 2413 2633
rect 2370 2563 2381 2566
rect 2370 2533 2373 2556
rect 2378 2533 2381 2563
rect 2354 2523 2365 2526
rect 2362 2426 2365 2523
rect 2354 2413 2357 2426
rect 2362 2423 2373 2426
rect 2330 2403 2349 2406
rect 2322 2383 2341 2386
rect 2282 2373 2317 2376
rect 2290 2323 2293 2336
rect 2314 2296 2317 2373
rect 2306 2293 2317 2296
rect 2266 2283 2285 2286
rect 2282 2213 2285 2283
rect 2306 2236 2309 2293
rect 2306 2233 2317 2236
rect 2290 2213 2301 2216
rect 2314 2173 2317 2233
rect 2322 2213 2325 2336
rect 2330 2323 2333 2376
rect 2338 2176 2341 2383
rect 2346 2323 2349 2403
rect 2354 2296 2357 2406
rect 2362 2333 2365 2416
rect 2370 2366 2373 2423
rect 2378 2403 2381 2496
rect 2386 2473 2389 2526
rect 2370 2363 2381 2366
rect 2350 2293 2357 2296
rect 2350 2236 2353 2293
rect 2362 2243 2365 2326
rect 2378 2266 2381 2363
rect 2394 2313 2397 2546
rect 2402 2533 2405 2556
rect 2410 2543 2413 2606
rect 2418 2586 2421 2616
rect 2418 2583 2429 2586
rect 2402 2413 2405 2426
rect 2410 2276 2413 2536
rect 2418 2493 2421 2526
rect 2426 2453 2429 2583
rect 2454 2576 2457 2653
rect 2450 2573 2457 2576
rect 2434 2513 2437 2526
rect 2442 2493 2445 2536
rect 2450 2533 2453 2573
rect 2370 2263 2381 2266
rect 2402 2273 2413 2276
rect 2370 2236 2373 2263
rect 2350 2233 2357 2236
rect 2370 2233 2381 2236
rect 2354 2183 2357 2233
rect 2362 2203 2365 2216
rect 2370 2213 2373 2226
rect 2338 2173 2349 2176
rect 2274 2123 2277 2136
rect 2290 2123 2293 2136
rect 2306 2133 2309 2146
rect 2314 2143 2333 2146
rect 2298 2056 2301 2126
rect 2314 2123 2317 2143
rect 2294 2053 2301 2056
rect 2258 2003 2261 2026
rect 2266 2003 2269 2016
rect 2282 2013 2285 2026
rect 2258 1983 2261 1996
rect 2274 1966 2277 2006
rect 2294 1996 2297 2053
rect 2294 1993 2301 1996
rect 2298 1976 2301 1993
rect 2298 1973 2309 1976
rect 2274 1963 2285 1966
rect 2282 1946 2285 1963
rect 2242 1903 2245 1926
rect 2266 1846 2269 1946
rect 2282 1943 2293 1946
rect 2242 1843 2269 1846
rect 2218 1743 2229 1746
rect 2218 1666 2221 1743
rect 2242 1733 2245 1843
rect 2250 1813 2253 1836
rect 2250 1783 2253 1806
rect 2258 1666 2261 1726
rect 2218 1663 2237 1666
rect 2210 1653 2229 1656
rect 2170 1633 2181 1636
rect 2170 1596 2173 1616
rect 2178 1603 2181 1633
rect 2186 1613 2189 1653
rect 2162 1593 2173 1596
rect 2162 1546 2165 1593
rect 2202 1566 2205 1606
rect 2178 1563 2205 1566
rect 2162 1543 2173 1546
rect 2162 1503 2165 1526
rect 2154 1333 2157 1346
rect 2162 1326 2165 1496
rect 2170 1423 2173 1543
rect 2178 1533 2181 1563
rect 2146 1323 2165 1326
rect 2058 1053 2069 1056
rect 2050 1013 2053 1036
rect 2042 933 2045 956
rect 2066 953 2069 1053
rect 2026 803 2029 916
rect 2042 913 2045 926
rect 2050 866 2053 936
rect 2034 863 2053 866
rect 2034 813 2037 863
rect 2058 823 2061 926
rect 1954 753 1965 756
rect 1994 773 2021 776
rect 1954 723 1957 753
rect 1914 613 1933 616
rect 1914 603 1917 613
rect 1938 603 1941 616
rect 1898 583 1901 596
rect 1962 593 1965 746
rect 1986 723 1989 736
rect 1994 733 1997 773
rect 1970 606 1973 626
rect 1970 603 1981 606
rect 1906 543 1909 566
rect 1930 543 1949 546
rect 1914 526 1917 536
rect 1930 533 1933 543
rect 1906 513 1909 526
rect 1914 523 1933 526
rect 1938 523 1941 536
rect 1834 333 1853 336
rect 1858 333 1861 396
rect 1866 366 1869 406
rect 1874 393 1877 406
rect 1866 363 1877 366
rect 1802 253 1813 256
rect 1794 183 1797 216
rect 1802 203 1805 236
rect 1810 213 1813 253
rect 1818 213 1821 326
rect 1834 316 1837 333
rect 1866 326 1869 356
rect 1842 323 1853 326
rect 1858 323 1869 326
rect 1874 323 1877 363
rect 1882 353 1885 436
rect 1898 416 1901 456
rect 1922 453 1925 496
rect 1938 466 1941 516
rect 1946 503 1949 543
rect 1954 476 1957 586
rect 1962 513 1965 536
rect 1970 523 1973 596
rect 1978 493 1981 603
rect 1986 583 1989 716
rect 2002 703 2005 726
rect 2002 593 2005 606
rect 2010 523 2013 736
rect 2018 613 2021 726
rect 2026 723 2037 726
rect 2026 666 2029 686
rect 2026 663 2033 666
rect 2030 606 2033 663
rect 2026 603 2033 606
rect 2026 493 2029 603
rect 2042 583 2045 756
rect 2066 753 2069 936
rect 2074 933 2077 1126
rect 2090 1123 2101 1126
rect 2082 983 2085 1016
rect 2090 1013 2093 1036
rect 2090 966 2093 996
rect 2098 973 2101 1123
rect 2114 1103 2117 1196
rect 2130 1163 2133 1216
rect 2154 1213 2157 1226
rect 2162 1193 2165 1316
rect 2170 1293 2173 1416
rect 2106 1013 2109 1026
rect 2106 996 2109 1006
rect 2114 1003 2117 1046
rect 2122 996 2125 1016
rect 2106 993 2125 996
rect 2130 983 2133 1136
rect 2146 1063 2149 1186
rect 2170 1156 2173 1256
rect 2178 1183 2181 1516
rect 2186 1503 2189 1536
rect 2194 1523 2213 1526
rect 2186 1313 2189 1476
rect 2194 1386 2197 1426
rect 2210 1413 2213 1506
rect 2218 1476 2221 1576
rect 2226 1533 2229 1653
rect 2234 1573 2237 1663
rect 2250 1663 2261 1666
rect 2226 1483 2229 1516
rect 2218 1473 2229 1476
rect 2202 1393 2205 1406
rect 2194 1383 2205 1386
rect 2194 1193 2197 1336
rect 2202 1216 2205 1383
rect 2210 1223 2213 1336
rect 2226 1333 2229 1473
rect 2234 1326 2237 1536
rect 2242 1403 2245 1626
rect 2250 1613 2253 1663
rect 2266 1573 2269 1776
rect 2250 1513 2253 1556
rect 2274 1533 2277 1826
rect 2290 1803 2293 1943
rect 2298 1813 2301 1926
rect 2282 1613 2285 1786
rect 2290 1633 2293 1756
rect 2298 1713 2301 1746
rect 2306 1656 2309 1973
rect 2314 1753 2317 2086
rect 2322 2023 2325 2136
rect 2330 2133 2333 2143
rect 2330 2113 2333 2126
rect 2338 2013 2341 2126
rect 2346 2093 2349 2173
rect 2378 2166 2381 2233
rect 2386 2213 2389 2246
rect 2394 2193 2397 2206
rect 2370 2163 2381 2166
rect 2370 2086 2373 2163
rect 2386 2133 2389 2146
rect 2402 2136 2405 2273
rect 2418 2203 2421 2226
rect 2394 2133 2405 2136
rect 2410 2126 2413 2186
rect 2426 2183 2429 2326
rect 2434 2306 2437 2336
rect 2442 2323 2445 2406
rect 2458 2333 2461 2456
rect 2466 2443 2469 2853
rect 2474 2623 2477 2756
rect 2482 2673 2485 2966
rect 2490 2896 2493 2976
rect 2498 2913 2501 2926
rect 2522 2906 2525 2983
rect 2546 2933 2549 2946
rect 2522 2903 2533 2906
rect 2490 2893 2497 2896
rect 2494 2756 2497 2893
rect 2506 2813 2509 2836
rect 2490 2753 2497 2756
rect 2490 2663 2493 2753
rect 2514 2733 2517 2796
rect 2530 2793 2533 2903
rect 2570 2853 2573 2926
rect 2546 2813 2549 2826
rect 2582 2786 2585 2993
rect 2594 2813 2597 2966
rect 2610 2943 2613 3016
rect 2634 3003 2637 3103
rect 2650 3046 2653 3126
rect 2674 3056 2677 3133
rect 2706 3123 2709 3196
rect 2730 3146 2733 3206
rect 2746 3183 2749 3206
rect 2758 3176 2761 3243
rect 2770 3213 2773 3236
rect 2778 3213 2781 3246
rect 2786 3213 2789 3236
rect 2834 3223 2837 3326
rect 2850 3313 2853 3433
rect 2858 3413 2861 3526
rect 2874 3513 2877 3526
rect 2882 3403 2885 3456
rect 2898 3386 2901 3616
rect 2906 3563 2909 3726
rect 2914 3613 2917 3763
rect 2922 3733 2925 3756
rect 2930 3733 2933 3746
rect 2930 3686 2933 3726
rect 2938 3723 2941 3763
rect 2946 3733 2949 3746
rect 2954 3723 2957 3736
rect 2962 3733 2965 3756
rect 2922 3683 2933 3686
rect 2914 3576 2917 3606
rect 2922 3593 2925 3683
rect 2930 3613 2933 3676
rect 2946 3613 2949 3706
rect 2978 3683 2981 3773
rect 3002 3723 3005 3746
rect 3010 3733 3013 3916
rect 3026 3886 3029 3926
rect 3018 3883 3029 3886
rect 3018 3803 3021 3883
rect 3026 3766 3029 3826
rect 3034 3803 3037 3886
rect 3050 3803 3053 3856
rect 3074 3853 3077 3966
rect 3090 3933 3093 3976
rect 3098 3826 3101 4016
rect 3114 4013 3117 4140
rect 3306 4063 3309 4140
rect 3106 3933 3109 4006
rect 3162 4003 3165 4016
rect 3210 4003 3213 4016
rect 3250 3983 3253 4016
rect 3122 3933 3125 3956
rect 3082 3823 3101 3826
rect 3022 3763 3029 3766
rect 3022 3686 3025 3763
rect 3082 3756 3085 3823
rect 3098 3776 3101 3816
rect 3114 3786 3117 3926
rect 3138 3863 3141 3936
rect 3170 3926 3173 3946
rect 3218 3933 3237 3936
rect 3162 3886 3165 3926
rect 3170 3923 3181 3926
rect 3218 3923 3221 3933
rect 3154 3883 3165 3886
rect 3114 3783 3125 3786
rect 3098 3773 3117 3776
rect 3082 3753 3093 3756
rect 3058 3733 3077 3736
rect 3058 3723 3061 3733
rect 3066 3713 3069 3726
rect 3082 3693 3085 3736
rect 3090 3726 3093 3753
rect 3114 3733 3117 3773
rect 3090 3723 3097 3726
rect 3022 3683 3029 3686
rect 2970 3613 2973 3666
rect 2914 3573 2925 3576
rect 2914 3413 2917 3516
rect 2922 3513 2925 3573
rect 2930 3483 2933 3576
rect 2938 3513 2941 3606
rect 2954 3573 2957 3606
rect 2962 3593 2965 3606
rect 2978 3603 2981 3626
rect 2986 3613 2989 3656
rect 2994 3613 2997 3626
rect 3026 3616 3029 3683
rect 3018 3613 3029 3616
rect 3034 3616 3037 3646
rect 3034 3613 3045 3616
rect 2994 3573 2997 3606
rect 2938 3416 2941 3446
rect 2946 3423 2949 3526
rect 2938 3413 2949 3416
rect 2890 3383 2901 3386
rect 2866 3333 2869 3366
rect 2850 3213 2853 3226
rect 2866 3216 2869 3326
rect 2874 3313 2877 3326
rect 2882 3223 2885 3336
rect 2890 3306 2893 3383
rect 2922 3366 2925 3406
rect 2938 3393 2941 3406
rect 2954 3403 2957 3566
rect 2970 3533 2973 3566
rect 3002 3563 3005 3606
rect 2962 3523 2973 3526
rect 2962 3413 2965 3516
rect 2978 3473 2981 3556
rect 2994 3516 2997 3536
rect 3010 3533 3013 3606
rect 3018 3573 3021 3613
rect 2994 3513 3001 3516
rect 2986 3423 2989 3486
rect 2998 3436 3001 3513
rect 2994 3433 3001 3436
rect 2994 3416 2997 3433
rect 2986 3413 2997 3416
rect 2962 3393 2965 3406
rect 2986 3383 2989 3413
rect 3002 3403 3005 3416
rect 2922 3363 2933 3366
rect 2898 3323 2901 3346
rect 2922 3333 2925 3346
rect 2890 3303 2901 3306
rect 2898 3236 2901 3303
rect 2914 3286 2917 3326
rect 2930 3323 2933 3363
rect 2938 3333 2941 3366
rect 2914 3283 2925 3286
rect 2890 3233 2901 3236
rect 2866 3213 2885 3216
rect 2890 3213 2893 3233
rect 2914 3213 2917 3226
rect 2922 3213 2925 3283
rect 2758 3173 2765 3176
rect 2730 3143 2741 3146
rect 2730 3123 2733 3136
rect 2738 3116 2741 3143
rect 2722 3096 2725 3116
rect 2714 3093 2725 3096
rect 2730 3113 2741 3116
rect 2674 3053 2681 3056
rect 2650 3043 2669 3046
rect 2626 2923 2629 2986
rect 2634 2923 2637 2996
rect 2658 2963 2661 3026
rect 2666 2983 2669 3043
rect 2678 2976 2681 3053
rect 2714 3036 2717 3093
rect 2714 3033 2725 3036
rect 2722 3013 2725 3033
rect 2714 3003 2725 3006
rect 2730 2996 2733 3113
rect 2762 3063 2765 3173
rect 2770 3133 2773 3206
rect 2802 3193 2805 3206
rect 2786 3123 2789 3136
rect 2810 3133 2813 3146
rect 2738 3023 2749 3026
rect 2746 3013 2749 3023
rect 2674 2973 2681 2976
rect 2722 2973 2725 2996
rect 2730 2993 2741 2996
rect 2778 2993 2781 3006
rect 2786 2993 2789 3026
rect 2794 3003 2797 3036
rect 2674 2833 2677 2973
rect 2738 2946 2741 2993
rect 2714 2933 2717 2946
rect 2730 2943 2741 2946
rect 2810 2943 2813 3026
rect 2826 3003 2829 3146
rect 2842 3116 2845 3136
rect 2838 3113 2845 3116
rect 2838 3036 2841 3113
rect 2850 3096 2853 3126
rect 2866 3123 2869 3166
rect 2890 3163 2893 3206
rect 2954 3193 2957 3336
rect 2978 3323 2981 3346
rect 2986 3306 2989 3376
rect 3010 3366 3013 3526
rect 3002 3363 3013 3366
rect 3002 3326 3005 3363
rect 2982 3303 2989 3306
rect 2994 3323 3005 3326
rect 2982 3236 2985 3303
rect 2982 3233 2989 3236
rect 2946 3133 2949 3146
rect 2850 3093 2861 3096
rect 2858 3046 2861 3093
rect 2850 3043 2861 3046
rect 2838 3033 2845 3036
rect 2834 3003 2837 3016
rect 2842 2993 2845 3033
rect 2850 3013 2853 3043
rect 2858 3023 2877 3026
rect 2858 3013 2861 3023
rect 2850 3003 2861 3006
rect 2690 2886 2693 2926
rect 2690 2883 2697 2886
rect 2682 2813 2685 2856
rect 2694 2806 2697 2883
rect 2714 2856 2717 2926
rect 2730 2923 2733 2943
rect 2762 2903 2765 2926
rect 2810 2923 2813 2936
rect 2826 2933 2829 2946
rect 2834 2913 2837 2936
rect 2842 2933 2845 2946
rect 2714 2853 2721 2856
rect 2582 2783 2589 2786
rect 2586 2766 2589 2783
rect 2626 2766 2629 2806
rect 2650 2793 2653 2806
rect 2690 2803 2697 2806
rect 2586 2763 2597 2766
rect 2626 2763 2637 2766
rect 2530 2713 2533 2726
rect 2538 2653 2541 2726
rect 2546 2703 2549 2726
rect 2594 2686 2597 2763
rect 2634 2733 2637 2763
rect 2690 2753 2693 2803
rect 2718 2786 2721 2853
rect 2850 2836 2853 2936
rect 2858 2916 2861 3003
rect 2866 2996 2869 3023
rect 2874 3006 2877 3016
rect 2882 3013 2885 3026
rect 2874 3003 2893 3006
rect 2898 3003 2901 3016
rect 2866 2993 2877 2996
rect 2866 2923 2869 2936
rect 2874 2933 2877 2993
rect 2890 2933 2893 3003
rect 2858 2913 2869 2916
rect 2866 2893 2869 2913
rect 2714 2783 2721 2786
rect 2714 2766 2717 2783
rect 2706 2763 2717 2766
rect 2730 2766 2733 2816
rect 2770 2813 2773 2836
rect 2850 2833 2861 2836
rect 2810 2813 2829 2816
rect 2746 2793 2749 2806
rect 2794 2776 2797 2796
rect 2786 2773 2797 2776
rect 2730 2763 2737 2766
rect 2666 2733 2669 2746
rect 2610 2713 2613 2726
rect 2690 2723 2693 2736
rect 2590 2683 2597 2686
rect 2706 2686 2709 2763
rect 2734 2686 2737 2763
rect 2706 2683 2717 2686
rect 2474 2523 2477 2616
rect 2498 2586 2501 2606
rect 2522 2586 2525 2606
rect 2498 2583 2525 2586
rect 2522 2563 2525 2583
rect 2482 2533 2485 2556
rect 2506 2543 2525 2546
rect 2490 2486 2493 2536
rect 2506 2523 2509 2543
rect 2490 2483 2509 2486
rect 2506 2426 2509 2483
rect 2514 2453 2517 2536
rect 2522 2533 2525 2543
rect 2522 2513 2525 2526
rect 2530 2506 2533 2546
rect 2546 2523 2549 2616
rect 2554 2583 2557 2626
rect 2590 2576 2593 2683
rect 2586 2573 2593 2576
rect 2554 2533 2557 2556
rect 2586 2536 2589 2573
rect 2578 2533 2589 2536
rect 2594 2533 2597 2546
rect 2602 2533 2605 2616
rect 2618 2613 2621 2626
rect 2522 2503 2533 2506
rect 2506 2423 2513 2426
rect 2474 2373 2477 2406
rect 2434 2303 2441 2306
rect 2438 2216 2441 2303
rect 2438 2213 2445 2216
rect 2370 2083 2381 2086
rect 2378 2063 2381 2083
rect 2394 2076 2397 2126
rect 2402 2123 2413 2126
rect 2418 2123 2421 2146
rect 2442 2143 2445 2213
rect 2450 2126 2453 2316
rect 2458 2213 2461 2226
rect 2466 2193 2469 2216
rect 2402 2083 2405 2123
rect 2434 2113 2437 2126
rect 2446 2123 2453 2126
rect 2394 2073 2413 2076
rect 2410 2013 2413 2073
rect 2446 2066 2449 2123
rect 2418 2006 2421 2066
rect 2446 2063 2453 2066
rect 2362 1993 2365 2006
rect 2346 1906 2349 1926
rect 2338 1903 2349 1906
rect 2338 1836 2341 1903
rect 2338 1833 2349 1836
rect 2322 1813 2341 1816
rect 2322 1803 2325 1813
rect 2330 1766 2333 1806
rect 2346 1803 2349 1833
rect 2354 1796 2357 1976
rect 2370 1826 2373 1986
rect 2386 1983 2389 2006
rect 2410 2003 2421 2006
rect 2410 1973 2413 2003
rect 2450 1983 2453 2063
rect 2458 1986 2461 2156
rect 2474 2126 2477 2326
rect 2490 2313 2493 2336
rect 2498 2323 2501 2416
rect 2510 2346 2513 2423
rect 2506 2343 2513 2346
rect 2506 2323 2509 2343
rect 2514 2306 2517 2326
rect 2510 2303 2517 2306
rect 2498 2213 2501 2226
rect 2510 2216 2513 2303
rect 2510 2213 2517 2216
rect 2482 2133 2485 2146
rect 2490 2133 2493 2166
rect 2466 2013 2469 2126
rect 2474 2123 2485 2126
rect 2474 1996 2477 2056
rect 2482 2013 2485 2123
rect 2490 2053 2493 2126
rect 2498 2013 2501 2186
rect 2506 2136 2509 2196
rect 2514 2153 2517 2213
rect 2522 2196 2525 2503
rect 2570 2493 2573 2526
rect 2578 2456 2581 2533
rect 2586 2523 2597 2526
rect 2570 2453 2581 2456
rect 2538 2426 2541 2446
rect 2538 2423 2549 2426
rect 2546 2356 2549 2423
rect 2570 2406 2573 2453
rect 2602 2446 2605 2526
rect 2610 2523 2613 2606
rect 2626 2543 2629 2616
rect 2594 2443 2605 2446
rect 2570 2403 2589 2406
rect 2538 2353 2549 2356
rect 2538 2293 2541 2353
rect 2554 2276 2557 2326
rect 2546 2273 2557 2276
rect 2522 2193 2533 2196
rect 2506 2133 2513 2136
rect 2510 2026 2513 2133
rect 2530 2086 2533 2193
rect 2546 2133 2549 2273
rect 2562 2203 2565 2336
rect 2578 2333 2581 2396
rect 2586 2333 2589 2403
rect 2594 2396 2597 2443
rect 2602 2413 2605 2436
rect 2618 2413 2621 2426
rect 2626 2413 2629 2536
rect 2634 2413 2637 2536
rect 2650 2533 2653 2556
rect 2642 2513 2645 2526
rect 2658 2506 2661 2666
rect 2666 2613 2669 2626
rect 2674 2553 2677 2676
rect 2666 2513 2669 2536
rect 2594 2393 2601 2396
rect 2570 2313 2573 2326
rect 2578 2276 2581 2296
rect 2574 2273 2581 2276
rect 2574 2196 2577 2273
rect 2586 2213 2589 2326
rect 2598 2226 2601 2393
rect 2610 2343 2613 2406
rect 2594 2223 2601 2226
rect 2574 2193 2581 2196
rect 2586 2193 2589 2206
rect 2578 2176 2581 2193
rect 2506 2023 2513 2026
rect 2522 2083 2533 2086
rect 2546 2083 2549 2126
rect 2554 2113 2557 2126
rect 2490 1996 2493 2006
rect 2506 2003 2509 2023
rect 2474 1993 2485 1996
rect 2490 1993 2517 1996
rect 2458 1983 2477 1986
rect 2378 1903 2381 1926
rect 2370 1823 2377 1826
rect 2346 1793 2357 1796
rect 2322 1763 2333 1766
rect 2314 1726 2317 1736
rect 2322 1733 2325 1763
rect 2338 1733 2341 1786
rect 2346 1733 2349 1793
rect 2354 1726 2357 1776
rect 2314 1723 2333 1726
rect 2346 1723 2357 1726
rect 2362 1723 2365 1816
rect 2374 1766 2377 1823
rect 2386 1803 2389 1966
rect 2426 1933 2429 1946
rect 2442 1923 2445 1936
rect 2394 1896 2397 1916
rect 2394 1893 2405 1896
rect 2402 1846 2405 1893
rect 2394 1843 2405 1846
rect 2394 1773 2397 1843
rect 2370 1763 2377 1766
rect 2306 1653 2325 1656
rect 2298 1593 2301 1626
rect 2258 1523 2277 1526
rect 2274 1503 2277 1516
rect 2282 1493 2285 1536
rect 2218 1323 2237 1326
rect 2202 1213 2209 1216
rect 2162 1153 2173 1156
rect 2162 1133 2165 1153
rect 2170 1143 2197 1146
rect 2170 1133 2173 1143
rect 2162 1113 2165 1126
rect 2138 1013 2141 1036
rect 2090 963 2101 966
rect 2098 933 2101 963
rect 2090 906 2093 926
rect 2098 913 2101 926
rect 2090 903 2109 906
rect 2058 613 2061 716
rect 2074 613 2077 836
rect 2082 813 2085 826
rect 2090 823 2093 856
rect 2082 803 2093 806
rect 2098 803 2101 866
rect 2106 773 2109 903
rect 2114 863 2117 956
rect 2122 813 2125 926
rect 2130 823 2133 936
rect 2138 913 2141 926
rect 2146 923 2149 1006
rect 2154 1003 2157 1106
rect 2162 983 2165 1016
rect 2170 1013 2173 1096
rect 2178 1083 2181 1126
rect 2194 1113 2197 1136
rect 2170 963 2173 1006
rect 2178 996 2181 1066
rect 2186 1013 2189 1106
rect 2206 1036 2209 1213
rect 2206 1033 2213 1036
rect 2194 1013 2205 1016
rect 2178 993 2197 996
rect 2162 923 2165 936
rect 2186 923 2189 986
rect 2194 906 2197 993
rect 2190 903 2197 906
rect 2138 816 2141 866
rect 2130 813 2141 816
rect 2146 813 2165 816
rect 2130 806 2133 813
rect 2114 793 2117 806
rect 2122 803 2133 806
rect 2082 716 2085 736
rect 2082 713 2093 716
rect 2090 636 2093 713
rect 2114 656 2117 786
rect 2138 723 2141 806
rect 2146 793 2149 813
rect 2082 633 2093 636
rect 2106 653 2117 656
rect 2082 613 2085 633
rect 2066 593 2069 606
rect 2074 603 2085 606
rect 1954 473 1965 476
rect 1938 463 1949 466
rect 1906 423 1909 436
rect 1898 413 1909 416
rect 1906 393 1909 413
rect 1914 413 1933 416
rect 1914 403 1917 413
rect 1930 393 1933 406
rect 1938 403 1941 436
rect 1834 313 1845 316
rect 1826 213 1829 276
rect 1842 273 1845 313
rect 1834 196 1837 206
rect 1842 203 1845 216
rect 1850 196 1853 216
rect 1858 203 1861 316
rect 1866 213 1869 323
rect 1834 193 1853 196
rect 1794 113 1797 126
rect 1818 103 1821 136
rect 1834 133 1837 186
rect 1874 133 1877 206
rect 1882 203 1885 346
rect 1930 343 1933 366
rect 1946 353 1949 463
rect 1954 393 1957 446
rect 1962 416 1965 473
rect 1962 413 1973 416
rect 1946 343 1965 346
rect 1890 293 1893 326
rect 1898 323 1901 336
rect 1930 326 1933 336
rect 1946 333 1949 343
rect 1906 283 1909 326
rect 1922 313 1925 326
rect 1930 323 1949 326
rect 1954 323 1957 336
rect 1954 293 1957 316
rect 1962 313 1965 343
rect 1970 323 1973 413
rect 1978 393 1981 406
rect 1994 403 1997 476
rect 2050 473 2053 546
rect 2074 533 2077 546
rect 1978 333 1989 336
rect 1994 326 1997 356
rect 1890 133 1893 216
rect 1906 213 1909 266
rect 1914 213 1917 276
rect 1954 266 1957 286
rect 1914 156 1917 206
rect 1922 203 1925 216
rect 1930 183 1933 216
rect 1938 203 1941 216
rect 1946 213 1949 266
rect 1954 263 1965 266
rect 1954 213 1957 263
rect 1978 223 1981 326
rect 1986 323 1997 326
rect 1986 293 1989 323
rect 2002 273 2005 346
rect 2010 323 2013 336
rect 2018 333 2021 406
rect 2034 333 2037 416
rect 2026 316 2029 326
rect 2042 323 2045 396
rect 2050 333 2053 356
rect 2066 336 2069 496
rect 2090 393 2093 416
rect 2098 356 2101 586
rect 2106 543 2109 653
rect 2122 593 2125 616
rect 2114 413 2117 516
rect 2122 403 2125 526
rect 2138 486 2141 626
rect 2146 566 2149 786
rect 2154 753 2157 806
rect 2170 783 2173 866
rect 2190 836 2193 903
rect 2178 833 2193 836
rect 2178 716 2181 833
rect 2186 766 2189 806
rect 2186 763 2197 766
rect 2194 723 2197 763
rect 2202 723 2205 986
rect 2210 883 2213 1033
rect 2218 986 2221 1306
rect 2258 1256 2261 1436
rect 2282 1393 2285 1416
rect 2290 1366 2293 1546
rect 2306 1456 2309 1576
rect 2322 1543 2325 1653
rect 2330 1573 2333 1716
rect 2346 1666 2349 1723
rect 2338 1663 2349 1666
rect 2338 1533 2341 1663
rect 2346 1603 2349 1616
rect 2314 1523 2333 1526
rect 2330 1503 2333 1516
rect 2302 1453 2309 1456
rect 2302 1376 2305 1453
rect 2346 1436 2349 1536
rect 2362 1493 2365 1716
rect 2370 1696 2373 1763
rect 2402 1746 2405 1826
rect 2418 1756 2421 1906
rect 2466 1813 2469 1926
rect 2474 1903 2477 1983
rect 2482 1976 2485 1993
rect 2482 1973 2489 1976
rect 2486 1896 2489 1973
rect 2482 1893 2489 1896
rect 2418 1753 2425 1756
rect 2402 1743 2413 1746
rect 2370 1693 2377 1696
rect 2374 1636 2377 1693
rect 2370 1633 2377 1636
rect 2338 1433 2349 1436
rect 2370 1433 2373 1633
rect 2386 1623 2389 1736
rect 2378 1593 2381 1616
rect 2386 1603 2389 1616
rect 2402 1583 2405 1616
rect 2338 1376 2341 1433
rect 2354 1413 2357 1426
rect 2302 1373 2309 1376
rect 2338 1373 2349 1376
rect 2282 1363 2293 1366
rect 2282 1286 2285 1363
rect 2306 1346 2309 1373
rect 2302 1343 2309 1346
rect 2282 1283 2293 1286
rect 2242 1253 2261 1256
rect 2226 1213 2229 1236
rect 2226 993 2229 1196
rect 2242 1163 2245 1253
rect 2266 1243 2269 1266
rect 2266 1213 2269 1226
rect 2290 1206 2293 1283
rect 2302 1266 2305 1343
rect 2314 1326 2317 1336
rect 2314 1323 2325 1326
rect 2330 1323 2333 1356
rect 2302 1263 2309 1266
rect 2266 1203 2293 1206
rect 2218 983 2229 986
rect 2226 863 2229 983
rect 2226 813 2229 826
rect 2234 776 2237 1136
rect 2242 1063 2245 1136
rect 2258 1076 2261 1126
rect 2266 1093 2269 1203
rect 2274 1133 2277 1146
rect 2282 1143 2301 1146
rect 2282 1123 2285 1143
rect 2290 1113 2293 1136
rect 2298 1133 2301 1143
rect 2306 1086 2309 1263
rect 2314 1196 2317 1316
rect 2322 1306 2325 1323
rect 2322 1303 2329 1306
rect 2326 1246 2329 1303
rect 2322 1243 2329 1246
rect 2322 1213 2325 1243
rect 2338 1223 2341 1336
rect 2346 1326 2349 1373
rect 2362 1333 2365 1406
rect 2346 1323 2365 1326
rect 2370 1233 2373 1416
rect 2362 1213 2365 1226
rect 2314 1193 2321 1196
rect 2318 1136 2321 1193
rect 2338 1163 2341 1206
rect 2318 1133 2341 1136
rect 2314 1093 2317 1126
rect 2322 1113 2325 1126
rect 2330 1103 2333 1126
rect 2306 1083 2317 1086
rect 2258 1073 2269 1076
rect 2266 1013 2269 1073
rect 2242 923 2245 1006
rect 2250 883 2253 936
rect 2258 903 2261 926
rect 2242 836 2245 856
rect 2266 836 2269 976
rect 2274 933 2277 1026
rect 2282 1003 2285 1016
rect 2290 933 2293 986
rect 2306 973 2309 1076
rect 2314 1003 2317 1083
rect 2338 1036 2341 1133
rect 2362 1113 2365 1126
rect 2370 1096 2373 1186
rect 2322 1033 2341 1036
rect 2366 1093 2373 1096
rect 2322 936 2325 1033
rect 2346 1003 2349 1016
rect 2354 963 2357 1016
rect 2366 956 2369 1093
rect 2378 1066 2381 1576
rect 2386 1503 2389 1516
rect 2386 1073 2389 1496
rect 2394 1253 2397 1566
rect 2410 1533 2413 1743
rect 2422 1686 2425 1753
rect 2450 1726 2453 1806
rect 2458 1793 2461 1806
rect 2474 1803 2477 1816
rect 2434 1713 2437 1726
rect 2450 1723 2469 1726
rect 2474 1713 2477 1726
rect 2482 1686 2485 1893
rect 2422 1683 2429 1686
rect 2418 1603 2421 1616
rect 2426 1613 2429 1683
rect 2474 1683 2485 1686
rect 2474 1636 2477 1683
rect 2498 1676 2501 1816
rect 2506 1706 2509 1986
rect 2522 1973 2525 2083
rect 2570 2076 2573 2176
rect 2578 2173 2585 2176
rect 2582 2076 2585 2173
rect 2594 2133 2597 2223
rect 2602 2193 2605 2206
rect 2610 2173 2613 2336
rect 2618 2256 2621 2276
rect 2618 2253 2625 2256
rect 2622 2176 2625 2253
rect 2618 2173 2625 2176
rect 2554 2073 2573 2076
rect 2578 2073 2585 2076
rect 2530 1943 2533 2016
rect 2538 1963 2541 2016
rect 2546 1983 2549 2006
rect 2514 1923 2525 1926
rect 2514 1906 2517 1923
rect 2554 1916 2557 2073
rect 2562 2003 2565 2036
rect 2570 2003 2573 2066
rect 2578 2053 2581 2073
rect 2578 2013 2581 2026
rect 2586 1996 2589 2006
rect 2562 1993 2589 1996
rect 2594 1976 2597 2126
rect 2602 2013 2605 2136
rect 2610 2123 2613 2156
rect 2618 2133 2621 2173
rect 2626 2133 2629 2156
rect 2626 2113 2629 2126
rect 2634 2106 2637 2346
rect 2642 2326 2645 2446
rect 2650 2333 2653 2506
rect 2658 2503 2669 2506
rect 2674 2503 2677 2546
rect 2642 2323 2649 2326
rect 2646 2276 2649 2323
rect 2658 2283 2661 2496
rect 2666 2473 2669 2503
rect 2682 2443 2685 2646
rect 2714 2643 2717 2683
rect 2730 2683 2737 2686
rect 2706 2533 2709 2606
rect 2722 2603 2725 2636
rect 2730 2623 2733 2683
rect 2730 2583 2733 2616
rect 2738 2603 2741 2656
rect 2746 2586 2749 2756
rect 2754 2736 2757 2766
rect 2754 2733 2765 2736
rect 2754 2663 2757 2726
rect 2754 2603 2757 2646
rect 2762 2613 2765 2733
rect 2770 2713 2773 2736
rect 2786 2686 2789 2773
rect 2802 2733 2805 2746
rect 2802 2693 2805 2726
rect 2786 2683 2797 2686
rect 2794 2643 2797 2683
rect 2762 2593 2765 2606
rect 2742 2583 2749 2586
rect 2690 2513 2693 2526
rect 2730 2513 2733 2526
rect 2742 2496 2745 2583
rect 2738 2493 2745 2496
rect 2666 2323 2669 2426
rect 2646 2273 2653 2276
rect 2642 2123 2645 2216
rect 2618 2103 2637 2106
rect 2562 1923 2565 1966
rect 2554 1913 2561 1916
rect 2514 1903 2525 1906
rect 2522 1836 2525 1903
rect 2514 1833 2525 1836
rect 2514 1803 2517 1833
rect 2546 1816 2549 1906
rect 2558 1836 2561 1913
rect 2558 1833 2565 1836
rect 2538 1793 2541 1816
rect 2546 1813 2557 1816
rect 2514 1713 2517 1736
rect 2522 1733 2525 1756
rect 2546 1736 2549 1813
rect 2534 1733 2549 1736
rect 2506 1703 2525 1706
rect 2490 1673 2501 1676
rect 2474 1633 2485 1636
rect 2426 1593 2429 1606
rect 2402 1513 2405 1526
rect 2402 1356 2405 1436
rect 2410 1363 2413 1456
rect 2426 1423 2429 1536
rect 2458 1533 2461 1626
rect 2482 1613 2485 1633
rect 2490 1613 2493 1673
rect 2498 1613 2509 1616
rect 2466 1593 2469 1606
rect 2434 1523 2453 1526
rect 2466 1516 2469 1586
rect 2450 1503 2453 1516
rect 2462 1513 2469 1516
rect 2462 1436 2465 1513
rect 2462 1433 2469 1436
rect 2442 1413 2461 1416
rect 2402 1353 2421 1356
rect 2402 1296 2405 1336
rect 2418 1333 2421 1353
rect 2434 1346 2437 1406
rect 2450 1376 2453 1406
rect 2450 1373 2457 1376
rect 2434 1343 2445 1346
rect 2442 1323 2445 1343
rect 2454 1306 2457 1373
rect 2466 1313 2469 1433
rect 2474 1363 2477 1546
rect 2514 1536 2517 1656
rect 2522 1543 2525 1703
rect 2534 1656 2537 1733
rect 2546 1713 2549 1726
rect 2530 1653 2537 1656
rect 2454 1303 2461 1306
rect 2402 1293 2413 1296
rect 2410 1236 2413 1293
rect 2402 1233 2413 1236
rect 2402 1216 2405 1233
rect 2402 1213 2421 1216
rect 2434 1213 2437 1236
rect 2426 1183 2429 1206
rect 2410 1093 2413 1136
rect 2434 1133 2437 1196
rect 2442 1183 2445 1256
rect 2458 1226 2461 1303
rect 2458 1223 2477 1226
rect 2482 1216 2485 1426
rect 2490 1413 2493 1536
rect 2514 1533 2525 1536
rect 2498 1523 2517 1526
rect 2514 1503 2517 1516
rect 2522 1486 2525 1533
rect 2514 1483 2525 1486
rect 2498 1413 2501 1446
rect 2514 1426 2517 1483
rect 2506 1423 2517 1426
rect 2458 1213 2485 1216
rect 2490 1206 2493 1366
rect 2498 1323 2501 1406
rect 2450 1146 2453 1206
rect 2482 1203 2493 1206
rect 2450 1143 2461 1146
rect 2458 1123 2461 1143
rect 2434 1106 2437 1116
rect 2418 1103 2437 1106
rect 2402 1066 2405 1076
rect 2378 1063 2405 1066
rect 2378 983 2381 1016
rect 2386 1003 2389 1063
rect 2402 1023 2413 1026
rect 2402 1013 2405 1023
rect 2418 1016 2421 1103
rect 2410 1013 2421 1016
rect 2394 1003 2405 1006
rect 2366 953 2373 956
rect 2314 933 2325 936
rect 2274 853 2277 916
rect 2242 833 2249 836
rect 2266 833 2273 836
rect 2226 773 2237 776
rect 2178 713 2205 716
rect 2186 613 2189 626
rect 2146 563 2157 566
rect 2130 483 2141 486
rect 2130 386 2133 483
rect 2154 476 2157 563
rect 2170 543 2173 606
rect 2186 583 2189 606
rect 2170 513 2173 526
rect 2146 473 2157 476
rect 2090 353 2101 356
rect 2114 383 2133 386
rect 2058 333 2069 336
rect 2074 333 2077 346
rect 2050 323 2061 326
rect 2050 316 2053 323
rect 2026 313 2053 316
rect 1986 213 2005 216
rect 1946 193 1949 206
rect 1986 203 1989 213
rect 2002 196 2005 206
rect 2010 203 2013 216
rect 2018 213 2021 266
rect 2026 196 2029 286
rect 2042 223 2045 296
rect 2058 293 2061 323
rect 1986 163 1989 196
rect 2002 193 2029 196
rect 2034 193 2037 206
rect 1914 153 1925 156
rect 1834 113 1837 126
rect 1914 113 1917 126
rect 1922 123 1925 153
rect 2002 133 2005 166
rect 2018 133 2021 186
rect 1954 113 1957 126
rect 2034 113 2037 126
rect 2042 123 2045 216
rect 2050 183 2053 246
rect 2058 213 2061 276
rect 2066 223 2069 333
rect 2082 246 2085 336
rect 2090 263 2093 353
rect 2098 256 2101 326
rect 2098 253 2109 256
rect 2074 236 2077 246
rect 2082 243 2101 246
rect 2074 233 2085 236
rect 2074 203 2077 216
rect 2082 203 2085 233
rect 2074 173 2077 196
rect 2090 193 2093 216
rect 2098 213 2101 243
rect 2106 203 2109 253
rect 2114 213 2117 383
rect 2138 353 2141 416
rect 2146 396 2149 473
rect 2154 413 2157 426
rect 2178 423 2181 536
rect 2194 513 2197 696
rect 2202 603 2205 713
rect 2210 703 2213 726
rect 2226 696 2229 773
rect 2246 726 2249 833
rect 2270 766 2273 833
rect 2282 793 2285 866
rect 2266 763 2273 766
rect 2266 746 2269 763
rect 2290 753 2293 926
rect 2298 813 2301 886
rect 2314 863 2317 933
rect 2306 803 2309 826
rect 2314 776 2317 836
rect 2322 803 2325 926
rect 2330 833 2333 946
rect 2338 823 2341 936
rect 2370 933 2373 953
rect 2402 943 2405 976
rect 2410 963 2413 1006
rect 2330 813 2349 816
rect 2354 813 2357 906
rect 2370 856 2373 926
rect 2386 923 2389 936
rect 2418 873 2421 1013
rect 2426 1003 2429 1016
rect 2434 996 2437 1086
rect 2466 1083 2469 1186
rect 2482 1113 2485 1203
rect 2498 1086 2501 1316
rect 2506 1306 2509 1423
rect 2530 1416 2533 1653
rect 2538 1533 2541 1636
rect 2554 1616 2557 1806
rect 2562 1653 2565 1833
rect 2546 1613 2557 1616
rect 2546 1603 2549 1613
rect 2562 1593 2565 1606
rect 2546 1516 2549 1536
rect 2570 1526 2573 1976
rect 2590 1973 2597 1976
rect 2590 1916 2593 1973
rect 2602 1923 2605 1976
rect 2578 1896 2581 1916
rect 2590 1913 2597 1916
rect 2578 1893 2585 1896
rect 2582 1796 2585 1893
rect 2578 1793 2585 1796
rect 2578 1633 2581 1793
rect 2586 1723 2589 1776
rect 2594 1753 2597 1913
rect 2602 1716 2605 1916
rect 2594 1713 2605 1716
rect 2594 1696 2597 1713
rect 2590 1693 2597 1696
rect 2590 1636 2593 1693
rect 2590 1633 2597 1636
rect 2578 1613 2589 1616
rect 2594 1533 2597 1633
rect 2602 1533 2605 1676
rect 2610 1583 2613 2056
rect 2618 1993 2621 2103
rect 2626 2003 2629 2056
rect 2634 1946 2637 2016
rect 2642 2013 2645 2026
rect 2650 1966 2653 2273
rect 2666 2216 2669 2236
rect 2658 2213 2669 2216
rect 2674 2216 2677 2336
rect 2682 2323 2685 2436
rect 2698 2306 2701 2476
rect 2738 2436 2741 2493
rect 2754 2446 2757 2586
rect 2770 2563 2773 2616
rect 2778 2613 2781 2636
rect 2786 2533 2789 2606
rect 2794 2593 2797 2626
rect 2802 2593 2805 2606
rect 2778 2523 2789 2526
rect 2794 2493 2797 2566
rect 2802 2476 2805 2586
rect 2810 2563 2813 2813
rect 2834 2793 2837 2806
rect 2818 2713 2821 2726
rect 2826 2713 2829 2736
rect 2842 2723 2845 2816
rect 2858 2803 2861 2833
rect 2818 2703 2829 2706
rect 2798 2473 2805 2476
rect 2754 2443 2765 2446
rect 2706 2413 2709 2426
rect 2722 2413 2725 2436
rect 2738 2433 2749 2436
rect 2694 2303 2701 2306
rect 2682 2223 2685 2256
rect 2694 2226 2697 2303
rect 2714 2296 2717 2406
rect 2722 2386 2725 2406
rect 2746 2403 2749 2433
rect 2722 2383 2733 2386
rect 2730 2296 2733 2383
rect 2690 2223 2697 2226
rect 2706 2293 2717 2296
rect 2722 2293 2733 2296
rect 2674 2213 2685 2216
rect 2658 1973 2661 2156
rect 2666 2063 2669 2206
rect 2674 2193 2677 2206
rect 2618 1943 2637 1946
rect 2618 1933 2621 1943
rect 2626 1933 2637 1936
rect 2642 1926 2645 1966
rect 2650 1963 2661 1966
rect 2618 1796 2621 1926
rect 2626 1813 2629 1926
rect 2634 1923 2645 1926
rect 2634 1906 2637 1923
rect 2634 1903 2641 1906
rect 2638 1836 2641 1903
rect 2634 1833 2641 1836
rect 2618 1793 2625 1796
rect 2622 1636 2625 1793
rect 2618 1633 2625 1636
rect 2634 1633 2637 1833
rect 2642 1793 2645 1816
rect 2650 1803 2653 1926
rect 2658 1906 2661 1963
rect 2674 1913 2677 2176
rect 2682 2143 2685 2213
rect 2690 2136 2693 2223
rect 2698 2193 2701 2216
rect 2706 2163 2709 2293
rect 2714 2233 2717 2286
rect 2722 2226 2725 2293
rect 2714 2223 2725 2226
rect 2714 2173 2717 2223
rect 2722 2153 2725 2216
rect 2730 2203 2733 2226
rect 2738 2213 2741 2276
rect 2746 2203 2749 2336
rect 2754 2316 2757 2336
rect 2786 2333 2789 2416
rect 2798 2346 2801 2473
rect 2810 2456 2813 2556
rect 2818 2523 2821 2703
rect 2834 2623 2837 2636
rect 2842 2623 2845 2716
rect 2850 2636 2853 2796
rect 2866 2723 2869 2736
rect 2874 2716 2877 2926
rect 2898 2923 2901 2976
rect 2914 2916 2917 3016
rect 2922 3003 2925 3126
rect 2962 3113 2965 3136
rect 2898 2913 2917 2916
rect 2922 2913 2925 2926
rect 2922 2816 2925 2906
rect 2890 2793 2893 2806
rect 2906 2793 2909 2816
rect 2914 2813 2925 2816
rect 2914 2803 2917 2813
rect 2930 2796 2933 2926
rect 2938 2903 2941 3086
rect 2970 3073 2973 3146
rect 2978 3083 2981 3216
rect 2986 3133 2989 3233
rect 2994 3133 2997 3323
rect 3018 3303 3021 3536
rect 3026 3513 3029 3606
rect 3034 3533 3037 3606
rect 3042 3563 3045 3613
rect 3050 3556 3053 3646
rect 3094 3636 3097 3723
rect 3094 3633 3101 3636
rect 3058 3613 3061 3626
rect 3058 3593 3061 3606
rect 3066 3573 3069 3606
rect 3050 3553 3061 3556
rect 3074 3553 3077 3616
rect 3082 3593 3085 3606
rect 3026 3433 3029 3476
rect 3026 3366 3029 3406
rect 3034 3403 3037 3506
rect 3042 3493 3045 3536
rect 3058 3496 3061 3553
rect 3074 3513 3077 3536
rect 3090 3523 3093 3616
rect 3098 3533 3101 3633
rect 3106 3593 3109 3726
rect 3114 3613 3117 3666
rect 3122 3643 3125 3783
rect 3130 3743 3133 3816
rect 3146 3813 3149 3826
rect 3138 3793 3141 3806
rect 3154 3803 3157 3883
rect 3138 3733 3141 3756
rect 3146 3706 3149 3726
rect 3142 3703 3149 3706
rect 3122 3603 3125 3616
rect 3130 3613 3133 3656
rect 3142 3636 3145 3703
rect 3142 3633 3149 3636
rect 3138 3603 3141 3616
rect 3146 3593 3149 3633
rect 3154 3613 3157 3676
rect 3162 3613 3165 3876
rect 3178 3846 3181 3923
rect 3226 3873 3229 3926
rect 3242 3873 3245 3976
rect 3250 3923 3253 3956
rect 3258 3933 3261 3976
rect 3170 3843 3181 3846
rect 3170 3803 3173 3843
rect 3258 3826 3261 3926
rect 3266 3923 3269 3996
rect 3274 3933 3277 4016
rect 3282 3993 3285 4026
rect 3330 4006 3333 4066
rect 3338 4013 3341 4026
rect 3330 4003 3349 4006
rect 3298 3963 3301 3996
rect 3254 3823 3261 3826
rect 3186 3783 3189 3806
rect 3170 3733 3173 3746
rect 3178 3723 3181 3736
rect 3218 3733 3221 3766
rect 3234 3733 3237 3816
rect 3254 3776 3257 3823
rect 3254 3773 3261 3776
rect 3170 3613 3173 3636
rect 3162 3586 3165 3606
rect 3178 3603 3181 3616
rect 3186 3613 3189 3646
rect 3210 3613 3213 3636
rect 3106 3533 3109 3556
rect 3058 3493 3077 3496
rect 3050 3413 3053 3426
rect 3042 3403 3053 3406
rect 3026 3363 3037 3366
rect 3034 3323 3037 3363
rect 3042 3333 3045 3366
rect 3050 3256 3053 3346
rect 3058 3286 3061 3416
rect 3066 3323 3069 3336
rect 3074 3293 3077 3493
rect 3098 3433 3101 3526
rect 3114 3496 3117 3526
rect 3106 3493 3117 3496
rect 3106 3443 3109 3493
rect 3058 3283 3069 3286
rect 3042 3253 3053 3256
rect 3018 3156 3021 3206
rect 3042 3193 3045 3253
rect 3010 3153 3021 3156
rect 3010 3143 3013 3153
rect 2946 3013 2949 3026
rect 2962 3016 2965 3026
rect 2954 3013 2965 3016
rect 2970 3013 2973 3026
rect 2978 3013 2981 3036
rect 2986 3023 2989 3126
rect 2946 2913 2949 2996
rect 2954 2933 2957 3006
rect 2994 2993 2997 3006
rect 3002 3003 3005 3136
rect 3010 3113 3013 3126
rect 3002 2933 3005 2946
rect 3018 2916 3021 3016
rect 3034 3013 3037 3126
rect 3066 3096 3069 3283
rect 3082 3213 3085 3336
rect 3090 3203 3093 3426
rect 3114 3423 3117 3486
rect 3098 3383 3101 3416
rect 3122 3413 3125 3536
rect 3130 3453 3133 3526
rect 3138 3516 3141 3576
rect 3146 3533 3149 3586
rect 3158 3583 3165 3586
rect 3138 3513 3145 3516
rect 3142 3446 3145 3513
rect 3158 3486 3161 3583
rect 3186 3566 3189 3606
rect 3138 3443 3145 3446
rect 3154 3483 3161 3486
rect 3170 3563 3189 3566
rect 3098 3333 3101 3366
rect 3114 3333 3117 3346
rect 3098 3313 3101 3326
rect 3090 3116 3093 3126
rect 3058 3093 3069 3096
rect 3082 3113 3093 3116
rect 3058 3046 3061 3093
rect 3058 3043 3069 3046
rect 3066 3023 3069 3043
rect 3050 2933 3053 3006
rect 3074 2986 3077 3016
rect 3058 2983 3077 2986
rect 3026 2923 3053 2926
rect 3018 2913 3029 2916
rect 3034 2903 3037 2916
rect 3050 2903 3053 2916
rect 3058 2913 3061 2983
rect 3066 2923 3069 2936
rect 2914 2793 2933 2796
rect 2914 2746 2917 2793
rect 2890 2743 2909 2746
rect 2914 2743 2925 2746
rect 2866 2713 2877 2716
rect 2882 2713 2885 2726
rect 2866 2703 2869 2713
rect 2890 2673 2893 2743
rect 2906 2716 2909 2736
rect 2902 2713 2909 2716
rect 2902 2646 2905 2713
rect 2902 2643 2909 2646
rect 2850 2633 2869 2636
rect 2826 2613 2853 2616
rect 2858 2613 2861 2626
rect 2810 2453 2821 2456
rect 2818 2376 2821 2453
rect 2810 2373 2821 2376
rect 2798 2343 2805 2346
rect 2754 2313 2765 2316
rect 2778 2313 2781 2326
rect 2762 2256 2765 2313
rect 2794 2266 2797 2326
rect 2754 2253 2765 2256
rect 2786 2263 2797 2266
rect 2786 2253 2789 2263
rect 2802 2256 2805 2343
rect 2794 2253 2805 2256
rect 2754 2223 2757 2253
rect 2762 2213 2765 2236
rect 2770 2213 2773 2226
rect 2754 2193 2757 2206
rect 2778 2183 2781 2216
rect 2682 2133 2693 2136
rect 2682 1923 2685 2133
rect 2690 2013 2693 2126
rect 2658 1903 2677 1906
rect 2658 1766 2661 1806
rect 2666 1793 2669 1806
rect 2650 1763 2661 1766
rect 2618 1536 2621 1633
rect 2610 1533 2621 1536
rect 2554 1523 2565 1526
rect 2570 1523 2581 1526
rect 2546 1513 2557 1516
rect 2562 1513 2565 1523
rect 2554 1416 2557 1513
rect 2570 1503 2573 1516
rect 2514 1323 2517 1416
rect 2530 1413 2541 1416
rect 2554 1413 2573 1416
rect 2506 1303 2513 1306
rect 2510 1226 2513 1303
rect 2522 1253 2525 1406
rect 2530 1363 2533 1406
rect 2538 1346 2541 1413
rect 2530 1343 2541 1346
rect 2546 1343 2549 1406
rect 2530 1303 2533 1343
rect 2538 1266 2541 1336
rect 2554 1326 2557 1356
rect 2562 1333 2565 1406
rect 2578 1353 2581 1523
rect 2610 1516 2613 1533
rect 2602 1513 2613 1516
rect 2618 1513 2621 1526
rect 2602 1386 2605 1513
rect 2610 1393 2613 1406
rect 2602 1383 2621 1386
rect 2546 1313 2549 1326
rect 2554 1323 2565 1326
rect 2538 1263 2557 1266
rect 2490 1083 2501 1086
rect 2506 1223 2513 1226
rect 2506 1083 2509 1223
rect 2554 1213 2557 1263
rect 2514 1123 2517 1206
rect 2530 1193 2533 1206
rect 2562 1196 2565 1323
rect 2558 1193 2565 1196
rect 2426 993 2437 996
rect 2426 866 2429 993
rect 2434 923 2437 986
rect 2442 966 2445 1016
rect 2458 983 2461 1026
rect 2442 963 2453 966
rect 2450 866 2453 963
rect 2466 923 2469 1006
rect 2474 1003 2477 1016
rect 2482 1013 2485 1056
rect 2490 1006 2493 1083
rect 2514 1076 2517 1116
rect 2506 1073 2517 1076
rect 2482 1003 2493 1006
rect 2482 896 2485 1003
rect 2498 993 2501 1046
rect 2506 1013 2509 1073
rect 2522 1013 2525 1136
rect 2498 946 2501 966
rect 2418 863 2429 866
rect 2442 863 2453 866
rect 2466 893 2485 896
rect 2494 943 2501 946
rect 2362 846 2365 856
rect 2370 853 2389 856
rect 2362 843 2373 846
rect 2370 823 2373 843
rect 2362 813 2373 816
rect 2346 806 2349 813
rect 2362 806 2365 813
rect 2306 773 2317 776
rect 2210 693 2229 696
rect 2242 723 2249 726
rect 2258 743 2269 746
rect 2210 553 2213 693
rect 2242 633 2245 723
rect 2226 546 2229 606
rect 2234 593 2237 616
rect 2242 583 2245 606
rect 2250 603 2253 706
rect 2258 693 2261 743
rect 2266 723 2269 736
rect 2290 723 2293 736
rect 2306 723 2309 773
rect 2322 766 2325 796
rect 2314 763 2325 766
rect 2338 766 2341 806
rect 2346 803 2365 806
rect 2370 803 2381 806
rect 2386 803 2389 853
rect 2394 803 2397 826
rect 2338 763 2349 766
rect 2314 733 2317 763
rect 2322 733 2333 736
rect 2290 613 2293 626
rect 2314 623 2317 636
rect 2298 613 2317 616
rect 2266 593 2269 606
rect 2170 413 2181 416
rect 2170 403 2173 413
rect 2146 393 2153 396
rect 2130 323 2133 346
rect 2138 306 2141 326
rect 2134 303 2141 306
rect 2134 236 2137 303
rect 2150 296 2153 393
rect 2194 356 2197 406
rect 2210 366 2213 546
rect 2226 543 2237 546
rect 2234 523 2237 543
rect 2298 483 2301 556
rect 2306 523 2309 596
rect 2314 573 2317 606
rect 2322 603 2325 626
rect 2330 566 2333 646
rect 2338 623 2341 726
rect 2346 716 2349 763
rect 2346 713 2357 716
rect 2354 656 2357 713
rect 2378 683 2381 756
rect 2402 723 2405 816
rect 2410 813 2413 836
rect 2410 706 2413 806
rect 2418 796 2421 863
rect 2426 813 2429 826
rect 2418 793 2425 796
rect 2406 703 2413 706
rect 2346 653 2357 656
rect 2314 563 2333 566
rect 2314 536 2317 563
rect 2314 533 2325 536
rect 2314 466 2317 526
rect 2322 493 2325 533
rect 2306 463 2317 466
rect 2258 413 2261 426
rect 2306 416 2309 463
rect 2330 423 2333 536
rect 2338 533 2341 616
rect 2346 533 2349 653
rect 2354 553 2357 636
rect 2370 603 2373 616
rect 2378 593 2381 606
rect 2362 533 2365 566
rect 2338 496 2341 526
rect 2338 493 2349 496
rect 2346 436 2349 493
rect 2338 433 2349 436
rect 2306 413 2317 416
rect 2338 413 2341 433
rect 2202 363 2213 366
rect 2202 356 2205 363
rect 2194 353 2205 356
rect 2178 333 2181 346
rect 2150 293 2165 296
rect 2134 233 2141 236
rect 2098 133 2101 186
rect 2114 183 2117 206
rect 2114 163 2125 166
rect 2130 163 2133 206
rect 2138 173 2141 233
rect 2146 203 2149 266
rect 2154 213 2157 226
rect 2162 206 2165 293
rect 2170 213 2181 216
rect 2154 203 2165 206
rect 2074 113 2077 126
rect 2122 113 2125 163
rect 2146 133 2149 186
rect 2154 166 2157 203
rect 2170 193 2173 206
rect 2186 203 2189 266
rect 2154 163 2165 166
rect 2162 143 2165 163
rect 2170 123 2173 166
rect 2202 163 2205 353
rect 2250 323 2253 346
rect 2290 263 2293 336
rect 2306 333 2309 376
rect 2314 326 2317 413
rect 2362 356 2365 526
rect 2386 523 2389 616
rect 2394 583 2397 696
rect 2406 626 2409 703
rect 2422 696 2425 793
rect 2418 693 2425 696
rect 2418 643 2421 693
rect 2402 623 2409 626
rect 2402 576 2405 623
rect 2410 593 2413 616
rect 2402 573 2409 576
rect 2394 476 2397 556
rect 2386 473 2397 476
rect 2354 353 2365 356
rect 2322 333 2325 346
rect 2330 333 2341 336
rect 2298 306 2301 326
rect 2306 316 2309 326
rect 2314 323 2325 326
rect 2330 323 2349 326
rect 2330 316 2333 323
rect 2306 313 2333 316
rect 2298 303 2309 306
rect 2226 193 2229 216
rect 2290 213 2301 216
rect 2306 213 2309 303
rect 2298 203 2309 206
rect 2314 203 2317 266
rect 2354 216 2357 353
rect 2370 293 2373 336
rect 2378 326 2381 426
rect 2386 423 2389 473
rect 2386 403 2389 416
rect 2394 413 2397 456
rect 2406 436 2409 573
rect 2402 433 2409 436
rect 2386 333 2389 346
rect 2402 336 2405 433
rect 2410 376 2413 416
rect 2418 403 2421 436
rect 2410 373 2421 376
rect 2394 333 2405 336
rect 2418 333 2421 373
rect 2426 333 2429 616
rect 2434 533 2437 686
rect 2442 613 2445 863
rect 2450 606 2453 856
rect 2466 846 2469 893
rect 2494 876 2497 943
rect 2506 933 2509 1006
rect 2514 936 2517 1006
rect 2514 933 2525 936
rect 2494 873 2501 876
rect 2498 853 2501 873
rect 2458 843 2469 846
rect 2458 726 2461 843
rect 2466 733 2469 796
rect 2458 723 2477 726
rect 2458 706 2461 723
rect 2458 703 2465 706
rect 2462 636 2465 703
rect 2458 633 2465 636
rect 2458 613 2461 633
rect 2442 523 2445 606
rect 2450 603 2461 606
rect 2450 506 2453 536
rect 2446 503 2453 506
rect 2446 436 2449 503
rect 2458 453 2461 603
rect 2474 573 2477 626
rect 2482 556 2485 806
rect 2506 803 2509 916
rect 2514 813 2517 926
rect 2522 783 2525 933
rect 2514 743 2517 756
rect 2490 696 2493 716
rect 2490 693 2501 696
rect 2514 693 2517 736
rect 2498 636 2501 693
rect 2490 633 2501 636
rect 2490 613 2493 633
rect 2498 593 2501 606
rect 2506 603 2509 616
rect 2514 613 2517 666
rect 2522 643 2525 726
rect 2530 646 2533 1186
rect 2538 1113 2541 1126
rect 2538 883 2541 1036
rect 2546 1013 2549 1126
rect 2558 1106 2561 1193
rect 2570 1183 2573 1306
rect 2578 1193 2581 1336
rect 2602 1323 2605 1346
rect 2610 1293 2613 1376
rect 2618 1366 2621 1383
rect 2626 1373 2629 1606
rect 2634 1596 2637 1616
rect 2642 1603 2645 1736
rect 2650 1613 2653 1763
rect 2658 1656 2661 1756
rect 2674 1726 2677 1903
rect 2690 1836 2693 1856
rect 2686 1833 2693 1836
rect 2686 1746 2689 1833
rect 2686 1743 2693 1746
rect 2674 1723 2681 1726
rect 2666 1673 2669 1716
rect 2678 1666 2681 1723
rect 2674 1663 2681 1666
rect 2658 1653 2665 1656
rect 2650 1596 2653 1606
rect 2634 1593 2653 1596
rect 2662 1586 2665 1653
rect 2634 1513 2637 1586
rect 2658 1583 2665 1586
rect 2618 1363 2629 1366
rect 2618 1286 2621 1356
rect 2626 1323 2629 1363
rect 2602 1283 2621 1286
rect 2602 1246 2605 1283
rect 2602 1243 2613 1246
rect 2594 1176 2597 1236
rect 2610 1176 2613 1243
rect 2626 1213 2629 1306
rect 2586 1173 2597 1176
rect 2602 1173 2613 1176
rect 2578 1113 2581 1126
rect 2558 1103 2565 1106
rect 2546 773 2549 936
rect 2554 833 2557 1086
rect 2562 973 2565 1103
rect 2586 1096 2589 1173
rect 2582 1093 2589 1096
rect 2582 1026 2585 1093
rect 2582 1023 2589 1026
rect 2562 913 2565 936
rect 2570 933 2573 1016
rect 2578 983 2581 1006
rect 2586 963 2589 1023
rect 2594 956 2597 1146
rect 2602 963 2605 1173
rect 2634 1156 2637 1276
rect 2642 1233 2645 1346
rect 2650 1313 2653 1536
rect 2658 1486 2661 1583
rect 2674 1563 2677 1663
rect 2666 1503 2669 1526
rect 2658 1483 2665 1486
rect 2662 1406 2665 1483
rect 2682 1456 2685 1636
rect 2690 1533 2693 1743
rect 2698 1733 2701 2026
rect 2722 2023 2725 2126
rect 2730 2113 2733 2176
rect 2722 1973 2725 2006
rect 2706 1946 2709 1966
rect 2738 1963 2741 2096
rect 2746 2083 2749 2136
rect 2762 2043 2765 2106
rect 2770 2026 2773 2126
rect 2762 2023 2773 2026
rect 2746 2003 2749 2016
rect 2762 1966 2765 2023
rect 2762 1963 2773 1966
rect 2706 1943 2713 1946
rect 2710 1876 2713 1943
rect 2746 1933 2749 1946
rect 2706 1873 2713 1876
rect 2706 1853 2709 1873
rect 2722 1813 2725 1926
rect 2762 1923 2765 1936
rect 2730 1833 2733 1856
rect 2706 1733 2709 1766
rect 2698 1513 2701 1726
rect 2730 1656 2733 1746
rect 2746 1713 2749 1916
rect 2754 1703 2765 1706
rect 2706 1613 2709 1636
rect 2714 1613 2717 1656
rect 2726 1653 2733 1656
rect 2726 1546 2729 1653
rect 2770 1646 2773 1963
rect 2778 1943 2781 2166
rect 2786 2123 2789 2236
rect 2794 2166 2797 2253
rect 2810 2233 2813 2373
rect 2818 2313 2821 2336
rect 2810 2213 2813 2226
rect 2826 2206 2829 2536
rect 2834 2506 2837 2606
rect 2866 2583 2869 2633
rect 2834 2503 2841 2506
rect 2838 2426 2841 2503
rect 2850 2463 2853 2536
rect 2858 2523 2861 2536
rect 2866 2523 2869 2546
rect 2874 2503 2877 2616
rect 2882 2603 2885 2636
rect 2906 2623 2909 2643
rect 2914 2613 2917 2736
rect 2922 2723 2925 2743
rect 2930 2703 2933 2736
rect 2938 2723 2941 2816
rect 2946 2716 2949 2806
rect 2954 2803 2957 2826
rect 2970 2803 2973 2846
rect 2962 2723 2965 2746
rect 2938 2713 2949 2716
rect 2970 2713 2973 2736
rect 2978 2733 2981 2836
rect 2994 2823 2997 2836
rect 3010 2803 3013 2826
rect 3018 2813 3021 2846
rect 2882 2553 2885 2596
rect 2930 2593 2933 2606
rect 2890 2536 2893 2586
rect 2882 2533 2893 2536
rect 2914 2533 2917 2586
rect 2938 2536 2941 2713
rect 2946 2543 2949 2676
rect 2954 2583 2957 2656
rect 2986 2653 2989 2796
rect 3026 2723 3029 2836
rect 3034 2833 3037 2846
rect 3042 2823 3045 2856
rect 3066 2823 3069 2836
rect 3074 2826 3077 2936
rect 3082 2873 3085 3113
rect 3114 3046 3117 3306
rect 3138 3213 3141 3443
rect 3154 3413 3157 3483
rect 3162 3403 3165 3416
rect 3170 3366 3173 3563
rect 3154 3363 3173 3366
rect 3154 3316 3157 3363
rect 3162 3323 3165 3346
rect 3154 3313 3165 3316
rect 3178 3313 3181 3556
rect 3186 3493 3189 3536
rect 3194 3503 3197 3566
rect 3202 3553 3205 3606
rect 3226 3593 3229 3726
rect 3242 3723 3245 3736
rect 3250 3733 3253 3756
rect 3234 3613 3237 3646
rect 3250 3613 3253 3636
rect 3258 3623 3261 3773
rect 3266 3743 3269 3816
rect 3274 3813 3277 3826
rect 3282 3733 3285 3926
rect 3290 3813 3293 3956
rect 3298 3933 3301 3946
rect 3298 3756 3301 3926
rect 3314 3856 3317 3936
rect 3330 3926 3333 3936
rect 3338 3933 3341 3956
rect 3322 3913 3325 3926
rect 3330 3923 3341 3926
rect 3314 3853 3325 3856
rect 3322 3813 3325 3853
rect 3338 3793 3341 3923
rect 3354 3886 3357 4026
rect 3370 3993 3373 4006
rect 3394 3996 3397 4016
rect 3450 4006 3453 4016
rect 3458 4013 3461 4026
rect 3450 4003 3469 4006
rect 3386 3993 3397 3996
rect 3490 3993 3493 4006
rect 3346 3883 3357 3886
rect 3370 3883 3373 3946
rect 3386 3933 3389 3993
rect 3394 3916 3397 3926
rect 3402 3923 3405 3936
rect 3386 3913 3397 3916
rect 3394 3903 3397 3913
rect 3298 3753 3305 3756
rect 3290 3733 3293 3746
rect 3186 3346 3189 3406
rect 3186 3343 3197 3346
rect 3194 3323 3197 3343
rect 3202 3323 3205 3536
rect 3210 3523 3213 3536
rect 3218 3533 3221 3556
rect 3210 3403 3213 3456
rect 3218 3403 3221 3526
rect 3226 3513 3229 3526
rect 3226 3413 3229 3446
rect 3234 3403 3237 3606
rect 3242 3546 3245 3606
rect 3258 3603 3261 3616
rect 3266 3593 3269 3726
rect 3274 3613 3277 3666
rect 3290 3613 3293 3716
rect 3302 3636 3305 3753
rect 3314 3733 3317 3746
rect 3298 3633 3305 3636
rect 3314 3633 3317 3726
rect 3242 3543 3253 3546
rect 3242 3523 3245 3536
rect 3250 3523 3253 3543
rect 3266 3523 3269 3536
rect 3274 3533 3277 3556
rect 3282 3523 3285 3606
rect 3298 3603 3301 3633
rect 3322 3603 3325 3786
rect 3330 3653 3333 3736
rect 3338 3643 3341 3786
rect 3346 3733 3349 3883
rect 3370 3803 3373 3866
rect 3386 3803 3389 3886
rect 3370 3663 3373 3726
rect 3378 3656 3381 3736
rect 3394 3733 3397 3816
rect 3402 3803 3405 3916
rect 3410 3823 3413 3926
rect 3442 3913 3445 3926
rect 3418 3816 3421 3906
rect 3450 3836 3453 3986
rect 3442 3833 3453 3836
rect 3410 3813 3421 3816
rect 3410 3773 3413 3813
rect 3418 3793 3421 3806
rect 3426 3803 3429 3816
rect 3434 3803 3437 3826
rect 3386 3693 3389 3726
rect 3362 3636 3365 3656
rect 3378 3653 3389 3656
rect 3418 3653 3421 3736
rect 3358 3633 3365 3636
rect 3146 3213 3149 3246
rect 3154 3213 3157 3296
rect 3162 3213 3165 3313
rect 3202 3296 3205 3316
rect 3194 3293 3205 3296
rect 3194 3236 3197 3293
rect 3194 3233 3205 3236
rect 3122 3096 3125 3146
rect 3130 3116 3133 3126
rect 3138 3123 3141 3206
rect 3162 3163 3165 3206
rect 3186 3193 3189 3216
rect 3202 3213 3205 3233
rect 3210 3213 3213 3366
rect 3226 3333 3229 3346
rect 3234 3313 3237 3326
rect 3242 3323 3245 3336
rect 3250 3276 3253 3486
rect 3266 3483 3269 3516
rect 3266 3413 3269 3446
rect 3290 3423 3293 3526
rect 3298 3503 3301 3516
rect 3322 3436 3325 3526
rect 3330 3493 3333 3516
rect 3346 3506 3349 3626
rect 3358 3586 3361 3633
rect 3370 3593 3373 3616
rect 3358 3583 3365 3586
rect 3346 3503 3357 3506
rect 3318 3433 3325 3436
rect 3258 3333 3261 3376
rect 3274 3326 3277 3346
rect 3242 3273 3253 3276
rect 3266 3323 3277 3326
rect 3242 3226 3245 3273
rect 3242 3223 3253 3226
rect 3194 3176 3197 3206
rect 3218 3183 3221 3216
rect 3226 3176 3229 3206
rect 3234 3183 3237 3206
rect 3194 3173 3229 3176
rect 3226 3153 3229 3173
rect 3234 3126 3237 3146
rect 3250 3143 3253 3223
rect 3146 3116 3149 3126
rect 3234 3123 3245 3126
rect 3130 3113 3149 3116
rect 3122 3093 3133 3096
rect 3090 3013 3093 3046
rect 3110 3043 3117 3046
rect 3098 3013 3101 3026
rect 3110 2986 3113 3043
rect 3130 3036 3133 3093
rect 3122 3033 3133 3036
rect 3122 3003 3125 3033
rect 3110 2983 3117 2986
rect 3114 2963 3117 2983
rect 3098 2943 3101 2956
rect 3090 2933 3117 2936
rect 3090 2923 3093 2933
rect 3098 2913 3101 2926
rect 3122 2903 3125 2926
rect 3082 2833 3085 2846
rect 3122 2833 3125 2846
rect 3130 2826 3133 2936
rect 3138 2923 3141 3006
rect 3146 2986 3149 3016
rect 3162 3003 3165 3016
rect 3170 3013 3173 3046
rect 3170 2996 3173 3006
rect 3186 3003 3189 3106
rect 3242 3036 3245 3123
rect 3250 3113 3253 3136
rect 3258 3103 3261 3206
rect 3266 3133 3269 3323
rect 3282 3306 3285 3416
rect 3278 3303 3285 3306
rect 3278 3246 3281 3303
rect 3278 3243 3285 3246
rect 3274 3213 3277 3226
rect 3282 3206 3285 3243
rect 3290 3213 3293 3406
rect 3298 3306 3301 3326
rect 3306 3323 3309 3406
rect 3318 3366 3321 3433
rect 3330 3373 3333 3426
rect 3318 3363 3325 3366
rect 3322 3343 3325 3363
rect 3298 3303 3305 3306
rect 3302 3236 3305 3303
rect 3322 3283 3325 3336
rect 3354 3313 3357 3503
rect 3362 3496 3365 3583
rect 3386 3576 3389 3653
rect 3442 3643 3445 3833
rect 3458 3803 3461 3866
rect 3490 3863 3493 3986
rect 3506 3923 3509 3936
rect 3514 3883 3517 3956
rect 3522 3896 3525 3936
rect 3530 3933 3533 4016
rect 3546 3933 3549 3976
rect 3554 3933 3557 3956
rect 3570 3943 3573 4016
rect 3586 3983 3589 4006
rect 3634 3976 3637 4016
rect 3634 3973 3645 3976
rect 3554 3913 3557 3926
rect 3562 3896 3565 3926
rect 3522 3893 3541 3896
rect 3450 3706 3453 3776
rect 3466 3723 3469 3746
rect 3450 3703 3461 3706
rect 3458 3646 3461 3703
rect 3450 3643 3461 3646
rect 3378 3573 3389 3576
rect 3370 3516 3373 3536
rect 3378 3523 3381 3573
rect 3386 3543 3413 3546
rect 3386 3533 3389 3543
rect 3394 3533 3405 3536
rect 3410 3533 3413 3543
rect 3418 3533 3421 3616
rect 3426 3576 3429 3616
rect 3450 3613 3453 3643
rect 3442 3593 3445 3606
rect 3426 3573 3437 3576
rect 3386 3516 3389 3526
rect 3370 3513 3389 3516
rect 3362 3493 3373 3496
rect 3370 3436 3373 3493
rect 3362 3433 3373 3436
rect 3362 3413 3365 3433
rect 3394 3413 3397 3533
rect 3402 3523 3413 3526
rect 3418 3493 3421 3526
rect 3394 3393 3397 3406
rect 3370 3323 3373 3346
rect 3298 3233 3305 3236
rect 3298 3213 3301 3233
rect 3274 3203 3285 3206
rect 3258 3053 3261 3096
rect 3194 3023 3221 3026
rect 3194 3013 3197 3023
rect 3210 3013 3221 3016
rect 3170 2993 3181 2996
rect 3146 2983 3165 2986
rect 3146 2906 3149 2936
rect 3154 2923 3157 2946
rect 3162 2933 3165 2983
rect 3170 2943 3173 2993
rect 3194 2966 3197 3006
rect 3202 3003 3221 3006
rect 3202 2973 3205 3003
rect 3170 2923 3173 2936
rect 3178 2906 3181 2966
rect 3194 2963 3221 2966
rect 3186 2933 3189 2956
rect 3194 2906 3197 2936
rect 3146 2903 3157 2906
rect 3154 2826 3157 2903
rect 3170 2903 3181 2906
rect 3186 2903 3197 2906
rect 3202 2903 3205 2926
rect 3170 2836 3173 2903
rect 3170 2833 3181 2836
rect 3074 2823 3093 2826
rect 3114 2823 3133 2826
rect 3050 2803 3053 2816
rect 3058 2813 3085 2816
rect 3122 2813 3133 2816
rect 3042 2723 3061 2726
rect 3034 2703 3037 2716
rect 2970 2593 2973 2646
rect 2994 2613 2997 2626
rect 2922 2533 2941 2536
rect 2882 2513 2885 2533
rect 2890 2516 2893 2526
rect 2898 2523 2917 2526
rect 2890 2513 2917 2516
rect 2838 2423 2845 2426
rect 2834 2323 2837 2416
rect 2842 2353 2845 2423
rect 2882 2406 2885 2486
rect 2866 2373 2869 2406
rect 2882 2403 2893 2406
rect 2874 2336 2877 2356
rect 2870 2333 2877 2336
rect 2842 2273 2845 2326
rect 2850 2313 2853 2326
rect 2858 2293 2861 2326
rect 2870 2286 2873 2333
rect 2890 2313 2893 2326
rect 2870 2283 2877 2286
rect 2874 2226 2877 2283
rect 2898 2253 2901 2496
rect 2906 2436 2909 2506
rect 2906 2433 2917 2436
rect 2906 2413 2909 2433
rect 2922 2416 2925 2533
rect 2930 2523 2941 2526
rect 2946 2483 2949 2536
rect 2954 2493 2957 2556
rect 2962 2533 2965 2566
rect 3002 2536 3005 2666
rect 3042 2633 3045 2716
rect 3082 2703 3085 2716
rect 3114 2713 3117 2726
rect 3130 2723 3133 2813
rect 3138 2716 3141 2826
rect 3122 2713 3141 2716
rect 3146 2823 3157 2826
rect 3146 2713 3149 2823
rect 3178 2813 3181 2833
rect 3186 2813 3189 2903
rect 3194 2806 3197 2886
rect 3154 2776 3157 2806
rect 3186 2803 3197 2806
rect 3154 2773 3165 2776
rect 3122 2703 3125 2713
rect 3162 2706 3165 2773
rect 3186 2753 3189 2803
rect 3202 2776 3205 2876
rect 3210 2866 3213 2916
rect 3218 2883 3221 2963
rect 3226 2943 3229 3016
rect 3234 2966 3237 3036
rect 3242 3033 3253 3036
rect 3250 3013 3253 3033
rect 3258 3023 3261 3036
rect 3266 3013 3269 3126
rect 3274 3093 3277 3203
rect 3282 3113 3285 3126
rect 3314 3123 3317 3226
rect 3330 3213 3333 3226
rect 3322 3133 3325 3206
rect 3330 3153 3333 3206
rect 3346 3203 3349 3286
rect 3402 3283 3405 3466
rect 3410 3403 3413 3456
rect 3418 3416 3421 3446
rect 3426 3426 3429 3536
rect 3434 3473 3437 3573
rect 3450 3533 3453 3606
rect 3458 3586 3461 3606
rect 3474 3593 3477 3656
rect 3498 3623 3501 3816
rect 3506 3813 3509 3836
rect 3538 3786 3541 3893
rect 3554 3893 3565 3896
rect 3554 3846 3557 3893
rect 3554 3843 3565 3846
rect 3562 3813 3565 3843
rect 3570 3833 3573 3936
rect 3578 3923 3581 3936
rect 3522 3783 3541 3786
rect 3514 3736 3517 3776
rect 3522 3746 3525 3783
rect 3578 3766 3581 3846
rect 3586 3813 3589 3956
rect 3594 3933 3597 3946
rect 3594 3866 3597 3926
rect 3626 3893 3629 3936
rect 3634 3923 3637 3936
rect 3642 3933 3645 3973
rect 3658 3933 3661 3966
rect 3666 3933 3669 4016
rect 3682 3983 3685 4006
rect 3706 3996 3709 4016
rect 3698 3993 3709 3996
rect 3594 3863 3605 3866
rect 3522 3743 3533 3746
rect 3514 3733 3525 3736
rect 3514 3713 3517 3726
rect 3530 3656 3533 3743
rect 3538 3733 3541 3746
rect 3554 3736 3557 3766
rect 3570 3763 3581 3766
rect 3554 3733 3565 3736
rect 3522 3653 3533 3656
rect 3498 3603 3501 3616
rect 3458 3583 3469 3586
rect 3442 3513 3445 3526
rect 3426 3423 3437 3426
rect 3418 3413 3429 3416
rect 3418 3393 3421 3406
rect 3426 3303 3429 3356
rect 3434 3323 3437 3423
rect 3458 3416 3461 3576
rect 3466 3533 3469 3583
rect 3522 3573 3525 3653
rect 3474 3513 3477 3536
rect 3490 3533 3493 3546
rect 3482 3523 3493 3526
rect 3482 3436 3485 3523
rect 3450 3413 3461 3416
rect 3474 3433 3485 3436
rect 3474 3413 3477 3433
rect 3498 3413 3501 3526
rect 3506 3523 3509 3536
rect 3522 3533 3525 3566
rect 3530 3533 3533 3546
rect 3514 3513 3517 3526
rect 3538 3523 3541 3726
rect 3546 3713 3549 3726
rect 3554 3696 3557 3726
rect 3550 3693 3557 3696
rect 3550 3626 3553 3693
rect 3562 3673 3565 3733
rect 3570 3693 3573 3763
rect 3586 3743 3589 3806
rect 3594 3766 3597 3836
rect 3602 3803 3605 3863
rect 3610 3803 3613 3826
rect 3594 3763 3613 3766
rect 3546 3623 3553 3626
rect 3546 3516 3549 3623
rect 3554 3563 3557 3616
rect 3562 3613 3565 3666
rect 3538 3513 3549 3516
rect 3450 3366 3453 3413
rect 3450 3363 3461 3366
rect 3442 3333 3445 3346
rect 3458 3343 3461 3363
rect 3450 3333 3461 3336
rect 3450 3316 3453 3326
rect 3466 3323 3469 3406
rect 3450 3313 3461 3316
rect 3482 3313 3485 3326
rect 3362 3173 3365 3206
rect 3386 3146 3389 3216
rect 3458 3213 3461 3313
rect 3490 3256 3493 3396
rect 3498 3323 3501 3406
rect 3506 3393 3509 3406
rect 3530 3396 3533 3416
rect 3538 3413 3541 3513
rect 3562 3496 3565 3606
rect 3586 3593 3589 3736
rect 3610 3663 3613 3763
rect 3618 3703 3621 3816
rect 3554 3493 3565 3496
rect 3522 3393 3533 3396
rect 3506 3316 3509 3346
rect 3522 3326 3525 3393
rect 3538 3366 3541 3406
rect 3546 3393 3549 3416
rect 3530 3363 3541 3366
rect 3530 3333 3533 3363
rect 3474 3253 3493 3256
rect 3498 3313 3509 3316
rect 3466 3223 3469 3246
rect 3466 3193 3469 3206
rect 3474 3176 3477 3253
rect 3490 3223 3493 3246
rect 3498 3213 3501 3313
rect 3514 3213 3517 3326
rect 3522 3323 3541 3326
rect 3370 3126 3373 3146
rect 3378 3143 3389 3146
rect 3378 3133 3381 3143
rect 3370 3123 3381 3126
rect 3250 2983 3253 3006
rect 3274 2973 3277 3056
rect 3234 2963 3245 2966
rect 3210 2863 3217 2866
rect 3214 2786 3217 2863
rect 3226 2813 3229 2826
rect 3226 2793 3229 2806
rect 3194 2773 3205 2776
rect 3210 2783 3217 2786
rect 3178 2713 3181 2726
rect 3154 2703 3165 2706
rect 3098 2646 3101 2696
rect 3098 2643 3109 2646
rect 2986 2533 3005 2536
rect 2986 2503 2989 2526
rect 3002 2513 3005 2526
rect 3026 2523 3037 2526
rect 2918 2413 2925 2416
rect 2962 2413 2965 2426
rect 2874 2223 2893 2226
rect 2810 2203 2829 2206
rect 2794 2163 2801 2166
rect 2778 1923 2781 1936
rect 2786 1913 2789 2116
rect 2798 1956 2801 2163
rect 2794 1953 2801 1956
rect 2794 1916 2797 1953
rect 2810 1946 2813 2203
rect 2858 2193 2861 2206
rect 2874 2176 2877 2216
rect 2874 2173 2885 2176
rect 2826 2133 2829 2146
rect 2818 2113 2821 2126
rect 2834 2106 2837 2126
rect 2830 2103 2837 2106
rect 2830 2036 2833 2103
rect 2830 2033 2837 2036
rect 2818 2003 2821 2016
rect 2810 1943 2817 1946
rect 2802 1923 2805 1936
rect 2794 1913 2805 1916
rect 2794 1873 2797 1906
rect 2802 1866 2805 1913
rect 2786 1863 2805 1866
rect 2786 1846 2789 1863
rect 2814 1846 2817 1943
rect 2826 1933 2829 2016
rect 2834 1933 2837 2033
rect 2782 1843 2789 1846
rect 2810 1843 2817 1846
rect 2782 1746 2785 1843
rect 2794 1823 2805 1826
rect 2810 1823 2813 1843
rect 2802 1816 2805 1823
rect 2818 1816 2821 1826
rect 2802 1813 2821 1816
rect 2826 1806 2829 1916
rect 2782 1743 2789 1746
rect 2794 1743 2797 1806
rect 2818 1803 2829 1806
rect 2818 1746 2821 1803
rect 2814 1743 2821 1746
rect 2786 1723 2789 1743
rect 2762 1643 2773 1646
rect 2746 1613 2749 1636
rect 2762 1596 2765 1643
rect 2794 1613 2797 1716
rect 2802 1633 2805 1706
rect 2814 1606 2817 1743
rect 2834 1716 2837 1726
rect 2842 1723 2845 2116
rect 2850 2056 2853 2126
rect 2858 2123 2861 2146
rect 2866 2113 2869 2136
rect 2882 2133 2885 2173
rect 2890 2123 2893 2223
rect 2906 2116 2909 2406
rect 2918 2346 2921 2413
rect 2914 2343 2921 2346
rect 2914 2286 2917 2343
rect 2914 2283 2921 2286
rect 2918 2196 2921 2283
rect 2938 2276 2941 2376
rect 2954 2333 2957 2386
rect 2938 2273 2957 2276
rect 2914 2193 2921 2196
rect 2930 2196 2933 2216
rect 2930 2193 2941 2196
rect 2954 2193 2957 2273
rect 2962 2233 2965 2326
rect 2970 2313 2973 2346
rect 2986 2343 2989 2416
rect 3002 2413 3005 2436
rect 3018 2423 3021 2496
rect 3026 2405 3029 2426
rect 3034 2403 3037 2516
rect 3042 2413 3045 2506
rect 3050 2486 3053 2616
rect 3074 2593 3077 2606
rect 3106 2596 3109 2643
rect 3122 2613 3125 2626
rect 3154 2623 3157 2703
rect 3098 2593 3109 2596
rect 3058 2496 3061 2586
rect 3066 2513 3069 2526
rect 3082 2523 3085 2546
rect 3058 2493 3069 2496
rect 3050 2483 3061 2486
rect 3050 2403 3053 2426
rect 3058 2413 3061 2483
rect 3066 2413 3069 2493
rect 3090 2436 3093 2526
rect 3098 2523 3101 2593
rect 3106 2543 3125 2546
rect 3106 2533 3109 2543
rect 3114 2513 3117 2536
rect 3122 2523 3125 2543
rect 3130 2523 3133 2546
rect 3138 2526 3141 2606
rect 3154 2546 3157 2616
rect 3162 2553 3165 2616
rect 3194 2613 3197 2773
rect 3210 2766 3213 2783
rect 3202 2763 3213 2766
rect 3202 2723 3205 2763
rect 3202 2703 3205 2716
rect 3210 2693 3213 2756
rect 3234 2753 3237 2956
rect 3242 2923 3245 2963
rect 3258 2943 3261 2956
rect 3282 2936 3285 3016
rect 3298 3013 3301 3106
rect 3306 3013 3309 3036
rect 3290 2993 3293 3006
rect 3298 2963 3301 3006
rect 3314 3003 3317 3106
rect 3322 3016 3325 3096
rect 3322 3013 3329 3016
rect 3266 2933 3285 2936
rect 3290 2933 3293 2956
rect 3250 2913 3253 2926
rect 3298 2923 3301 2946
rect 3306 2916 3309 2926
rect 3290 2833 3293 2916
rect 3298 2913 3309 2916
rect 3306 2843 3309 2913
rect 3314 2833 3317 2976
rect 3326 2956 3329 3013
rect 3322 2953 3329 2956
rect 3322 2923 3325 2953
rect 3330 2836 3333 2936
rect 3338 2923 3341 3016
rect 3346 2996 3349 3106
rect 3354 3003 3357 3016
rect 3362 3003 3365 3016
rect 3370 3003 3373 3026
rect 3378 3013 3381 3123
rect 3386 3113 3389 3136
rect 3402 3133 3405 3176
rect 3470 3173 3477 3176
rect 3346 2993 3357 2996
rect 3346 2933 3349 2986
rect 3354 2973 3357 2993
rect 3362 2933 3365 2996
rect 3330 2833 3341 2836
rect 3242 2813 3245 2826
rect 3338 2816 3341 2833
rect 3234 2713 3237 2726
rect 3258 2706 3261 2726
rect 3266 2723 3269 2816
rect 3330 2813 3341 2816
rect 3346 2813 3349 2836
rect 3354 2823 3357 2926
rect 3330 2793 3333 2813
rect 3354 2808 3357 2816
rect 3362 2813 3365 2926
rect 3370 2813 3373 2976
rect 3378 2913 3381 2956
rect 3258 2703 3269 2706
rect 3274 2703 3277 2746
rect 3282 2723 3301 2726
rect 3146 2543 3157 2546
rect 3162 2543 3181 2546
rect 3146 2533 3149 2543
rect 3138 2523 3149 2526
rect 3082 2433 3093 2436
rect 3074 2413 3077 2426
rect 3066 2383 3069 2406
rect 3074 2393 3077 2406
rect 3082 2393 3085 2433
rect 3010 2336 3013 2376
rect 2994 2326 2997 2336
rect 3010 2333 3021 2336
rect 3050 2333 3053 2356
rect 2994 2323 3029 2326
rect 3026 2273 3029 2323
rect 3058 2313 3061 2326
rect 3066 2323 3069 2376
rect 3050 2236 3053 2256
rect 2914 2173 2917 2193
rect 2922 2133 2933 2136
rect 2938 2133 2941 2193
rect 2946 2126 2949 2166
rect 2978 2146 2981 2206
rect 2914 2123 2933 2126
rect 2942 2123 2949 2126
rect 2954 2143 2981 2146
rect 2906 2113 2917 2116
rect 2914 2066 2917 2113
rect 2914 2063 2925 2066
rect 2850 2053 2861 2056
rect 2858 1963 2861 2053
rect 2882 1993 2885 2016
rect 2906 1973 2909 2026
rect 2866 1936 2869 1956
rect 2850 1933 2869 1936
rect 2850 1923 2853 1933
rect 2858 1913 2861 1926
rect 2874 1923 2885 1926
rect 2866 1733 2869 1836
rect 2882 1833 2885 1923
rect 2890 1913 2893 1966
rect 2898 1936 2901 1946
rect 2898 1933 2909 1936
rect 2762 1593 2773 1596
rect 2794 1593 2797 1606
rect 2810 1603 2817 1606
rect 2826 1713 2837 1716
rect 2726 1543 2733 1546
rect 2682 1453 2693 1456
rect 2662 1403 2669 1406
rect 2658 1323 2661 1396
rect 2666 1353 2669 1403
rect 2674 1393 2677 1416
rect 2674 1306 2677 1376
rect 2690 1343 2693 1453
rect 2650 1303 2677 1306
rect 2650 1203 2653 1303
rect 2698 1286 2701 1506
rect 2714 1493 2717 1516
rect 2722 1446 2725 1526
rect 2714 1443 2725 1446
rect 2706 1313 2709 1436
rect 2682 1283 2701 1286
rect 2682 1266 2685 1283
rect 2714 1273 2717 1443
rect 2730 1436 2733 1543
rect 2738 1523 2741 1556
rect 2746 1533 2749 1546
rect 2754 1463 2757 1576
rect 2722 1433 2733 1436
rect 2722 1366 2725 1433
rect 2730 1413 2733 1426
rect 2738 1415 2741 1436
rect 2754 1416 2757 1436
rect 2746 1413 2757 1416
rect 2730 1386 2733 1406
rect 2738 1403 2749 1406
rect 2738 1393 2741 1403
rect 2754 1386 2757 1396
rect 2730 1383 2757 1386
rect 2722 1363 2741 1366
rect 2722 1323 2725 1346
rect 2678 1263 2685 1266
rect 2678 1156 2681 1263
rect 2690 1166 2693 1256
rect 2698 1193 2701 1216
rect 2690 1163 2697 1166
rect 2634 1153 2653 1156
rect 2678 1153 2685 1156
rect 2626 1123 2629 1136
rect 2578 953 2597 956
rect 2570 896 2573 926
rect 2562 893 2573 896
rect 2562 873 2565 893
rect 2570 816 2573 886
rect 2578 873 2581 953
rect 2586 943 2605 946
rect 2586 923 2589 943
rect 2594 923 2597 936
rect 2602 933 2605 943
rect 2610 923 2613 1006
rect 2618 1003 2621 1036
rect 2626 973 2629 1016
rect 2554 813 2565 816
rect 2570 813 2581 816
rect 2586 813 2589 916
rect 2618 886 2621 966
rect 2610 883 2621 886
rect 2634 883 2637 1106
rect 2642 1033 2645 1136
rect 2650 1126 2653 1153
rect 2650 1123 2661 1126
rect 2666 1123 2669 1146
rect 2658 1026 2661 1036
rect 2642 1023 2661 1026
rect 2642 1013 2645 1023
rect 2666 1016 2669 1106
rect 2674 1073 2677 1136
rect 2674 1036 2677 1056
rect 2682 1046 2685 1153
rect 2694 1076 2697 1163
rect 2706 1123 2717 1126
rect 2722 1103 2725 1306
rect 2738 1276 2741 1363
rect 2734 1273 2741 1276
rect 2734 1136 2737 1273
rect 2734 1133 2741 1136
rect 2738 1113 2741 1133
rect 2690 1073 2697 1076
rect 2690 1053 2693 1073
rect 2682 1043 2693 1046
rect 2674 1033 2681 1036
rect 2650 1003 2653 1016
rect 2658 1013 2669 1016
rect 2658 946 2661 1013
rect 2666 953 2669 996
rect 2678 976 2681 1033
rect 2678 973 2685 976
rect 2658 943 2669 946
rect 2642 913 2645 926
rect 2650 923 2661 926
rect 2666 916 2669 943
rect 2682 933 2685 973
rect 2650 913 2669 916
rect 2682 913 2685 926
rect 2602 813 2605 836
rect 2538 663 2541 766
rect 2546 716 2549 736
rect 2554 733 2557 813
rect 2562 806 2565 813
rect 2562 803 2573 806
rect 2546 713 2553 716
rect 2550 646 2553 713
rect 2530 643 2541 646
rect 2530 613 2533 636
rect 2538 606 2541 643
rect 2482 553 2493 556
rect 2482 533 2485 546
rect 2434 416 2437 436
rect 2446 433 2453 436
rect 2450 416 2453 433
rect 2434 413 2453 416
rect 2378 323 2389 326
rect 2378 216 2381 316
rect 2386 223 2389 323
rect 2394 223 2397 333
rect 2402 323 2421 326
rect 2402 303 2413 306
rect 2418 303 2421 323
rect 2330 213 2349 216
rect 2354 213 2373 216
rect 2378 213 2389 216
rect 2298 186 2301 203
rect 2290 183 2301 186
rect 2242 123 2245 176
rect 2258 133 2261 166
rect 2290 126 2293 183
rect 2322 166 2325 206
rect 2330 203 2341 206
rect 2306 163 2325 166
rect 2290 123 2301 126
rect 2306 123 2309 163
rect 2346 156 2349 206
rect 2386 203 2389 213
rect 2338 153 2349 156
rect 2338 123 2341 153
rect 2298 103 2301 123
rect 2354 113 2357 136
rect 2394 123 2397 216
rect 2402 63 2405 266
rect 2410 216 2413 303
rect 2426 286 2429 326
rect 2434 323 2437 406
rect 2466 403 2469 416
rect 2474 413 2477 516
rect 2482 513 2485 526
rect 2490 506 2493 553
rect 2522 543 2525 606
rect 2530 603 2541 606
rect 2546 643 2553 646
rect 2482 503 2493 506
rect 2442 333 2445 386
rect 2426 283 2437 286
rect 2410 213 2421 216
rect 2410 193 2413 206
rect 2418 183 2421 206
rect 2426 193 2429 216
rect 2434 123 2437 283
rect 2442 213 2445 326
rect 2450 303 2453 396
rect 2466 346 2469 386
rect 2458 343 2469 346
rect 2442 123 2445 206
rect 2450 183 2453 226
rect 2458 203 2461 343
rect 2466 323 2469 336
rect 2466 293 2469 316
rect 2482 293 2485 503
rect 2490 393 2493 456
rect 2514 386 2517 536
rect 2522 523 2525 536
rect 2530 506 2533 603
rect 2538 523 2541 596
rect 2546 586 2549 643
rect 2562 633 2565 776
rect 2570 733 2573 756
rect 2578 733 2581 813
rect 2586 733 2597 736
rect 2578 663 2581 726
rect 2554 603 2557 626
rect 2562 593 2565 616
rect 2570 603 2573 646
rect 2586 623 2589 726
rect 2594 703 2597 733
rect 2602 643 2605 806
rect 2610 773 2613 883
rect 2618 766 2621 876
rect 2650 873 2653 913
rect 2666 886 2669 896
rect 2634 823 2653 826
rect 2626 796 2629 816
rect 2634 803 2637 823
rect 2642 796 2645 806
rect 2626 793 2645 796
rect 2610 763 2621 766
rect 2610 626 2613 763
rect 2594 623 2613 626
rect 2546 583 2565 586
rect 2578 583 2581 606
rect 2530 503 2541 506
rect 2538 446 2541 503
rect 2530 443 2541 446
rect 2530 413 2533 443
rect 2562 436 2565 583
rect 2594 563 2597 623
rect 2602 536 2605 616
rect 2578 493 2581 536
rect 2586 533 2605 536
rect 2562 433 2581 436
rect 2514 383 2525 386
rect 2506 273 2509 356
rect 2466 196 2469 216
rect 2474 203 2477 226
rect 2482 196 2485 206
rect 2466 193 2485 196
rect 2490 123 2493 216
rect 2498 123 2501 216
rect 2522 113 2525 383
rect 2538 366 2541 406
rect 2546 403 2549 416
rect 2554 406 2557 416
rect 2562 413 2565 433
rect 2570 413 2573 426
rect 2554 403 2565 406
rect 2538 363 2557 366
rect 2530 303 2533 326
rect 2538 203 2541 226
rect 2546 93 2549 296
rect 2554 203 2557 363
rect 2562 323 2565 403
rect 2570 333 2573 406
rect 2578 333 2581 433
rect 2602 413 2605 526
rect 2610 423 2613 616
rect 2618 593 2621 606
rect 2626 583 2629 756
rect 2634 613 2637 726
rect 2642 596 2645 726
rect 2650 703 2653 823
rect 2658 753 2661 886
rect 2666 883 2677 886
rect 2666 803 2669 876
rect 2674 753 2677 883
rect 2682 783 2685 896
rect 2690 823 2693 1043
rect 2698 983 2701 996
rect 2674 696 2677 736
rect 2690 733 2693 816
rect 2698 743 2701 966
rect 2706 943 2709 976
rect 2714 953 2717 1006
rect 2722 996 2725 1096
rect 2730 1003 2733 1076
rect 2722 993 2733 996
rect 2706 893 2709 936
rect 2730 933 2733 993
rect 2738 973 2741 1016
rect 2746 933 2749 1376
rect 2762 1356 2765 1526
rect 2770 1373 2773 1593
rect 2810 1586 2813 1603
rect 2802 1583 2813 1586
rect 2778 1423 2781 1526
rect 2786 1426 2789 1566
rect 2794 1523 2797 1536
rect 2802 1523 2805 1583
rect 2794 1433 2797 1466
rect 2810 1433 2813 1536
rect 2818 1533 2821 1556
rect 2818 1513 2821 1526
rect 2826 1496 2829 1713
rect 2834 1683 2837 1706
rect 2822 1493 2829 1496
rect 2822 1426 2825 1493
rect 2786 1423 2805 1426
rect 2822 1423 2829 1426
rect 2754 1353 2765 1356
rect 2754 1296 2757 1353
rect 2778 1346 2781 1406
rect 2786 1393 2789 1416
rect 2786 1373 2789 1386
rect 2762 1343 2781 1346
rect 2762 1323 2765 1343
rect 2770 1333 2781 1336
rect 2786 1333 2789 1346
rect 2770 1313 2773 1326
rect 2794 1323 2797 1416
rect 2802 1386 2805 1423
rect 2802 1383 2813 1386
rect 2754 1293 2765 1296
rect 2762 1146 2765 1293
rect 2778 1213 2781 1226
rect 2786 1213 2789 1316
rect 2802 1266 2805 1376
rect 2810 1276 2813 1383
rect 2818 1333 2821 1406
rect 2826 1286 2829 1423
rect 2834 1373 2837 1636
rect 2842 1623 2845 1716
rect 2850 1633 2853 1646
rect 2858 1613 2861 1636
rect 2842 1323 2845 1556
rect 2866 1553 2869 1626
rect 2866 1533 2869 1546
rect 2850 1523 2861 1526
rect 2858 1503 2861 1523
rect 2850 1386 2853 1486
rect 2858 1403 2861 1446
rect 2866 1413 2869 1436
rect 2850 1383 2857 1386
rect 2854 1316 2857 1383
rect 2866 1333 2869 1346
rect 2874 1333 2877 1726
rect 2882 1533 2885 1796
rect 2882 1433 2885 1526
rect 2890 1483 2893 1826
rect 2882 1393 2885 1406
rect 2882 1333 2885 1356
rect 2890 1343 2893 1426
rect 2898 1413 2901 1926
rect 2906 1716 2909 1933
rect 2914 1906 2917 1946
rect 2922 1923 2925 2063
rect 2930 2003 2933 2096
rect 2942 2026 2945 2123
rect 2938 2023 2945 2026
rect 2954 2023 2957 2143
rect 2970 2106 2973 2136
rect 2966 2103 2973 2106
rect 2966 2026 2969 2103
rect 2966 2023 2973 2026
rect 2930 1926 2933 1936
rect 2938 1933 2941 2023
rect 2954 1953 2957 2016
rect 2962 1993 2965 2006
rect 2970 1986 2973 2023
rect 2978 2013 2981 2126
rect 2962 1983 2973 1986
rect 2954 1933 2957 1946
rect 2930 1923 2949 1926
rect 2914 1903 2925 1906
rect 2946 1903 2949 1923
rect 2922 1836 2925 1903
rect 2914 1833 2925 1836
rect 2914 1733 2917 1833
rect 2906 1713 2913 1716
rect 2910 1626 2913 1713
rect 2906 1623 2913 1626
rect 2922 1626 2925 1816
rect 2930 1733 2933 1806
rect 2946 1793 2949 1836
rect 2922 1623 2933 1626
rect 2906 1603 2909 1623
rect 2930 1603 2933 1623
rect 2938 1613 2941 1636
rect 2898 1386 2901 1406
rect 2898 1383 2909 1386
rect 2898 1336 2901 1376
rect 2906 1353 2909 1383
rect 2914 1353 2917 1536
rect 2938 1523 2941 1546
rect 2946 1443 2949 1736
rect 2954 1613 2957 1916
rect 2962 1723 2965 1983
rect 2970 1903 2973 1926
rect 2978 1856 2981 2006
rect 2970 1853 2981 1856
rect 2970 1766 2973 1853
rect 2986 1833 2989 2136
rect 2994 2023 2997 2176
rect 3002 2133 3005 2216
rect 3002 2096 3005 2126
rect 3010 2113 3013 2126
rect 3002 2093 3009 2096
rect 2986 1803 2989 1816
rect 2970 1763 2981 1766
rect 2978 1716 2981 1763
rect 2994 1723 2997 2016
rect 3006 1866 3009 2093
rect 3002 1863 3009 1866
rect 3002 1773 3005 1863
rect 3018 1846 3021 2146
rect 3026 2136 3029 2236
rect 3046 2233 3053 2236
rect 3026 2133 3037 2136
rect 3026 2113 3029 2126
rect 3034 2123 3037 2133
rect 3034 2033 3037 2066
rect 3046 2026 3049 2233
rect 3058 2133 3061 2216
rect 3066 2213 3069 2276
rect 3082 2256 3085 2336
rect 3090 2316 3093 2416
rect 3098 2383 3101 2466
rect 3106 2403 3109 2416
rect 3114 2403 3117 2436
rect 3122 2413 3125 2456
rect 3146 2406 3149 2523
rect 3154 2493 3157 2536
rect 3162 2523 3165 2543
rect 3170 2523 3173 2536
rect 3178 2533 3181 2543
rect 3186 2523 3189 2556
rect 3194 2543 3205 2546
rect 3194 2523 3197 2543
rect 3162 2423 3165 2506
rect 3138 2376 3141 2406
rect 3146 2403 3165 2406
rect 3162 2383 3165 2403
rect 3170 2376 3173 2486
rect 3202 2433 3205 2526
rect 3218 2463 3221 2536
rect 3242 2533 3245 2606
rect 3258 2546 3261 2696
rect 3266 2603 3269 2703
rect 3282 2656 3285 2723
rect 3306 2716 3309 2756
rect 3278 2653 3285 2656
rect 3298 2713 3309 2716
rect 3314 2716 3317 2736
rect 3330 2733 3333 2766
rect 3338 2756 3341 2806
rect 3346 2805 3357 2808
rect 3346 2763 3349 2805
rect 3338 2753 3357 2756
rect 3314 2713 3325 2716
rect 3278 2586 3281 2653
rect 3290 2613 3293 2646
rect 3290 2593 3293 2606
rect 3278 2583 3285 2586
rect 3258 2543 3269 2546
rect 3194 2413 3197 2426
rect 3226 2423 3229 2526
rect 3218 2413 3237 2416
rect 3218 2403 3229 2406
rect 3138 2373 3165 2376
rect 3170 2373 3181 2376
rect 3098 2333 3109 2336
rect 3138 2333 3141 2346
rect 3090 2313 3101 2316
rect 3078 2253 3085 2256
rect 3046 2023 3053 2026
rect 3026 1913 3029 1936
rect 3034 1873 3037 1976
rect 3010 1843 3021 1846
rect 3010 1743 3013 1843
rect 3034 1803 3037 1856
rect 3042 1833 3045 2006
rect 3050 1973 3053 2023
rect 3058 1966 3061 2126
rect 3050 1963 3061 1966
rect 3050 1903 3053 1963
rect 3066 1953 3069 2196
rect 3078 2136 3081 2253
rect 3098 2246 3101 2313
rect 3122 2256 3125 2326
rect 3162 2323 3165 2373
rect 3178 2316 3181 2373
rect 3218 2323 3221 2403
rect 3234 2396 3237 2413
rect 3226 2393 3237 2396
rect 3242 2396 3245 2516
rect 3266 2513 3269 2543
rect 3274 2516 3277 2556
rect 3282 2523 3285 2583
rect 3298 2566 3301 2713
rect 3322 2656 3325 2713
rect 3346 2703 3349 2726
rect 3354 2723 3357 2753
rect 3370 2723 3373 2806
rect 3378 2803 3381 2826
rect 3386 2813 3389 2936
rect 3394 2823 3397 2976
rect 3402 2913 3405 3126
rect 3426 3013 3429 3126
rect 3470 3116 3473 3173
rect 3482 3123 3485 3196
rect 3498 3133 3501 3206
rect 3470 3113 3477 3116
rect 3434 3013 3437 3036
rect 3434 2946 3437 2996
rect 3418 2936 3421 2946
rect 3434 2943 3445 2946
rect 3410 2933 3421 2936
rect 3442 2933 3445 2943
rect 3410 2896 3413 2933
rect 3418 2923 3437 2926
rect 3418 2913 3429 2916
rect 3434 2903 3437 2923
rect 3410 2893 3421 2896
rect 3394 2733 3397 2816
rect 3418 2813 3421 2893
rect 3434 2823 3437 2836
rect 3442 2813 3445 2926
rect 3450 2913 3453 3006
rect 3466 3003 3469 3026
rect 3474 2973 3477 3113
rect 3458 2906 3461 2936
rect 3466 2923 3469 2956
rect 3482 2916 3485 3016
rect 3490 2973 3493 3016
rect 3506 3013 3509 3026
rect 3522 3013 3525 3286
rect 3506 3003 3517 3006
rect 3522 2993 3525 3006
rect 3530 2966 3533 3316
rect 3538 3203 3541 3276
rect 3546 3206 3549 3336
rect 3554 3323 3557 3493
rect 3562 3403 3565 3416
rect 3570 3403 3573 3506
rect 3578 3483 3581 3556
rect 3578 3413 3581 3456
rect 3594 3413 3597 3446
rect 3586 3393 3589 3406
rect 3562 3273 3565 3346
rect 3554 3213 3557 3236
rect 3546 3203 3557 3206
rect 3538 2983 3541 3186
rect 3562 3166 3565 3206
rect 3546 3163 3565 3166
rect 3546 3123 3549 3163
rect 3546 3013 3549 3116
rect 3570 3083 3573 3386
rect 3602 3366 3605 3526
rect 3610 3506 3613 3526
rect 3610 3503 3617 3506
rect 3614 3416 3617 3503
rect 3614 3413 3621 3416
rect 3626 3413 3629 3806
rect 3634 3783 3637 3826
rect 3642 3803 3645 3816
rect 3650 3793 3653 3926
rect 3682 3883 3685 3936
rect 3698 3933 3701 3993
rect 3690 3913 3693 3926
rect 3706 3906 3709 3936
rect 3702 3903 3709 3906
rect 3658 3803 3661 3816
rect 3634 3723 3637 3746
rect 3634 3593 3637 3616
rect 3634 3493 3637 3516
rect 3650 3513 3653 3636
rect 3658 3583 3661 3736
rect 3666 3566 3669 3806
rect 3674 3763 3677 3826
rect 3690 3813 3693 3846
rect 3702 3836 3705 3903
rect 3714 3853 3717 3956
rect 3730 3933 3733 3946
rect 3746 3933 3749 3986
rect 3762 3943 3765 4016
rect 3778 3993 3781 4026
rect 3826 3993 3829 4016
rect 3858 4006 3861 4016
rect 3858 4003 3877 4006
rect 3850 3933 3853 3976
rect 3722 3836 3725 3926
rect 3702 3833 3709 3836
rect 3706 3813 3709 3833
rect 3714 3813 3717 3836
rect 3722 3833 3733 3836
rect 3674 3676 3677 3756
rect 3682 3713 3685 3806
rect 3690 3793 3693 3806
rect 3706 3753 3709 3806
rect 3690 3696 3693 3736
rect 3706 3733 3709 3746
rect 3698 3713 3701 3726
rect 3714 3723 3717 3806
rect 3722 3783 3725 3806
rect 3722 3733 3725 3746
rect 3730 3733 3733 3833
rect 3738 3733 3741 3826
rect 3746 3813 3749 3896
rect 3746 3743 3749 3806
rect 3754 3793 3757 3836
rect 3690 3693 3701 3696
rect 3674 3673 3685 3676
rect 3682 3606 3685 3673
rect 3662 3563 3669 3566
rect 3674 3603 3685 3606
rect 3698 3603 3701 3693
rect 3662 3516 3665 3563
rect 3674 3523 3677 3603
rect 3706 3543 3709 3616
rect 3714 3593 3717 3606
rect 3662 3513 3669 3516
rect 3642 3413 3645 3466
rect 3610 3393 3613 3406
rect 3594 3363 3605 3366
rect 3594 3346 3597 3363
rect 3590 3343 3597 3346
rect 3578 3203 3581 3306
rect 3590 3286 3593 3343
rect 3602 3333 3605 3356
rect 3602 3296 3605 3326
rect 3618 3313 3621 3413
rect 3602 3293 3613 3296
rect 3626 3293 3629 3386
rect 3642 3353 3645 3406
rect 3650 3373 3653 3496
rect 3666 3446 3669 3513
rect 3662 3443 3669 3446
rect 3662 3346 3665 3443
rect 3662 3343 3669 3346
rect 3666 3323 3669 3343
rect 3674 3306 3677 3436
rect 3690 3413 3693 3436
rect 3682 3326 3685 3406
rect 3698 3376 3701 3456
rect 3706 3403 3709 3536
rect 3714 3433 3717 3576
rect 3714 3413 3717 3426
rect 3722 3413 3725 3726
rect 3730 3703 3733 3726
rect 3730 3583 3733 3606
rect 3722 3376 3725 3406
rect 3730 3393 3733 3546
rect 3738 3533 3741 3716
rect 3746 3706 3749 3736
rect 3754 3723 3757 3766
rect 3762 3733 3765 3896
rect 3794 3876 3797 3926
rect 3786 3856 3789 3876
rect 3794 3873 3805 3876
rect 3770 3803 3773 3856
rect 3782 3853 3789 3856
rect 3782 3766 3785 3853
rect 3782 3763 3789 3766
rect 3746 3703 3757 3706
rect 3754 3636 3757 3703
rect 3746 3633 3757 3636
rect 3746 3533 3749 3633
rect 3754 3573 3757 3616
rect 3770 3603 3773 3736
rect 3778 3723 3781 3746
rect 3786 3616 3789 3763
rect 3794 3723 3797 3826
rect 3802 3803 3805 3873
rect 3810 3796 3813 3816
rect 3818 3803 3821 3886
rect 3842 3813 3845 3926
rect 3850 3893 3853 3926
rect 3858 3923 3861 3946
rect 3866 3933 3869 3996
rect 3882 3943 3885 4016
rect 3874 3923 3877 3936
rect 3882 3923 3885 3936
rect 3890 3933 3893 3976
rect 3898 3953 3901 4026
rect 3970 4023 3989 4026
rect 3922 3976 3925 4016
rect 3970 4006 3973 4023
rect 3906 3973 3925 3976
rect 3966 4003 3973 4006
rect 3978 4006 3981 4016
rect 3986 4013 3989 4023
rect 3978 4003 3997 4006
rect 3906 3933 3909 3973
rect 3866 3796 3869 3816
rect 3802 3793 3813 3796
rect 3802 3733 3805 3793
rect 3794 3683 3797 3716
rect 3802 3703 3805 3726
rect 3810 3693 3813 3736
rect 3778 3593 3781 3616
rect 3786 3613 3797 3616
rect 3818 3613 3821 3736
rect 3826 3663 3829 3796
rect 3850 3793 3869 3796
rect 3874 3793 3877 3806
rect 3834 3733 3837 3756
rect 3842 3733 3845 3766
rect 3842 3713 3845 3726
rect 3850 3723 3853 3793
rect 3882 3786 3885 3816
rect 3866 3783 3885 3786
rect 3858 3706 3861 3736
rect 3866 3723 3869 3783
rect 3890 3753 3893 3926
rect 3914 3876 3917 3926
rect 3922 3923 3925 3936
rect 3930 3933 3933 3966
rect 3966 3936 3969 4003
rect 3946 3916 3949 3936
rect 3966 3933 3973 3936
rect 3938 3913 3949 3916
rect 3914 3873 3925 3876
rect 3914 3803 3917 3816
rect 3922 3813 3925 3873
rect 3938 3846 3941 3913
rect 3938 3843 3949 3846
rect 3914 3773 3917 3796
rect 3930 3793 3933 3806
rect 3874 3723 3877 3736
rect 3882 3733 3885 3746
rect 3882 3713 3885 3726
rect 3898 3713 3901 3736
rect 3906 3723 3909 3736
rect 3914 3733 3917 3756
rect 3922 3733 3925 3746
rect 3938 3743 3941 3826
rect 3946 3803 3949 3843
rect 3954 3786 3957 3926
rect 3970 3913 3973 3933
rect 3978 3886 3981 3986
rect 3986 3923 3989 3936
rect 3994 3933 3997 3996
rect 4010 3983 4013 4006
rect 4034 3993 4037 4016
rect 4090 4006 4093 4016
rect 4090 4003 4109 4006
rect 4002 3906 4005 3946
rect 4010 3916 4013 3936
rect 4010 3913 4021 3916
rect 3970 3883 3981 3886
rect 3998 3903 4005 3906
rect 3970 3803 3973 3883
rect 3998 3836 4001 3903
rect 4018 3866 4021 3913
rect 4010 3863 4021 3866
rect 3998 3833 4005 3836
rect 3994 3803 3997 3816
rect 3954 3783 3965 3786
rect 3858 3703 3869 3706
rect 3786 3556 3789 3606
rect 3794 3583 3797 3613
rect 3770 3553 3789 3556
rect 3754 3533 3757 3546
rect 3770 3533 3773 3553
rect 3786 3546 3789 3553
rect 3778 3533 3781 3546
rect 3786 3543 3797 3546
rect 3698 3373 3709 3376
rect 3722 3373 3733 3376
rect 3690 3333 3693 3346
rect 3682 3323 3693 3326
rect 3706 3323 3709 3373
rect 3714 3333 3717 3346
rect 3722 3323 3725 3336
rect 3730 3333 3733 3373
rect 3738 3333 3741 3446
rect 3746 3413 3749 3526
rect 3762 3443 3765 3526
rect 3666 3303 3677 3306
rect 3590 3283 3597 3286
rect 3594 3213 3597 3283
rect 3610 3226 3613 3293
rect 3602 3223 3613 3226
rect 3666 3226 3669 3303
rect 3666 3223 3677 3226
rect 3578 3123 3581 3196
rect 3602 3183 3605 3223
rect 3618 3193 3621 3206
rect 3594 3133 3597 3146
rect 3634 3046 3637 3126
rect 3642 3123 3645 3136
rect 3658 3126 3661 3206
rect 3674 3196 3677 3223
rect 3682 3203 3685 3216
rect 3690 3213 3693 3323
rect 3706 3213 3709 3296
rect 3722 3256 3725 3276
rect 3718 3253 3725 3256
rect 3674 3193 3693 3196
rect 3658 3123 3677 3126
rect 3682 3123 3685 3166
rect 3690 3093 3693 3193
rect 3698 3133 3701 3206
rect 3718 3176 3721 3253
rect 3730 3183 3733 3326
rect 3738 3213 3741 3326
rect 3746 3323 3749 3356
rect 3754 3333 3757 3346
rect 3762 3303 3765 3416
rect 3770 3403 3773 3526
rect 3786 3523 3789 3536
rect 3794 3506 3797 3543
rect 3790 3503 3797 3506
rect 3778 3413 3781 3446
rect 3790 3436 3793 3503
rect 3790 3433 3797 3436
rect 3794 3413 3797 3433
rect 3802 3423 3805 3596
rect 3810 3493 3813 3516
rect 3810 3413 3813 3436
rect 3746 3213 3749 3236
rect 3762 3213 3765 3246
rect 3770 3206 3773 3336
rect 3778 3233 3781 3406
rect 3786 3353 3789 3406
rect 3794 3393 3797 3406
rect 3826 3403 3829 3606
rect 3850 3553 3853 3686
rect 3866 3626 3869 3703
rect 3858 3623 3869 3626
rect 3858 3603 3861 3623
rect 3866 3593 3869 3606
rect 3842 3533 3845 3546
rect 3850 3446 3853 3536
rect 3850 3443 3861 3446
rect 3834 3413 3837 3426
rect 3786 3296 3789 3336
rect 3786 3293 3793 3296
rect 3790 3236 3793 3293
rect 3786 3233 3793 3236
rect 3786 3213 3789 3233
rect 3754 3193 3757 3206
rect 3762 3203 3773 3206
rect 3718 3173 3725 3176
rect 3634 3043 3645 3046
rect 3578 3006 3581 3016
rect 3578 3003 3589 3006
rect 3514 2963 3533 2966
rect 3490 2923 3501 2926
rect 3466 2913 3477 2916
rect 3482 2913 3493 2916
rect 3458 2903 3469 2906
rect 3458 2853 3461 2903
rect 3458 2823 3461 2846
rect 3466 2813 3469 2836
rect 3442 2743 3445 2806
rect 3474 2796 3477 2826
rect 3470 2793 3477 2796
rect 3470 2736 3473 2793
rect 3482 2743 3485 2826
rect 3498 2813 3501 2923
rect 3506 2903 3509 2916
rect 3514 2856 3517 2963
rect 3522 2916 3525 2926
rect 3530 2923 3533 2956
rect 3554 2936 3557 2946
rect 3538 2916 3541 2936
rect 3522 2913 3541 2916
rect 3538 2896 3541 2913
rect 3530 2893 3541 2896
rect 3546 2933 3557 2936
rect 3562 2933 3565 2946
rect 3514 2853 3521 2856
rect 3506 2833 3509 2846
rect 3490 2753 3493 2766
rect 3498 2746 3501 2806
rect 3490 2743 3501 2746
rect 3458 2713 3461 2736
rect 3470 2733 3477 2736
rect 3314 2653 3325 2656
rect 3306 2613 3309 2646
rect 3314 2633 3317 2653
rect 3298 2563 3309 2566
rect 3306 2546 3309 2563
rect 3306 2543 3313 2546
rect 3274 2513 3285 2516
rect 3250 2408 3253 2486
rect 3282 2433 3285 2513
rect 3310 2486 3313 2543
rect 3306 2483 3313 2486
rect 3322 2536 3325 2596
rect 3394 2593 3397 2616
rect 3402 2603 3405 2626
rect 3410 2613 3413 2706
rect 3474 2633 3477 2733
rect 3490 2703 3493 2743
rect 3498 2673 3501 2726
rect 3506 2693 3509 2826
rect 3518 2786 3521 2853
rect 3530 2836 3533 2893
rect 3530 2833 3541 2836
rect 3538 2813 3541 2833
rect 3546 2816 3549 2933
rect 3570 2926 3573 2996
rect 3586 2993 3589 3003
rect 3634 2993 3637 3006
rect 3586 2933 3589 2966
rect 3594 2933 3597 2986
rect 3554 2913 3557 2926
rect 3562 2923 3573 2926
rect 3562 2823 3565 2923
rect 3546 2813 3565 2816
rect 3570 2813 3573 2826
rect 3514 2783 3521 2786
rect 3530 2783 3533 2806
rect 3538 2793 3541 2806
rect 3562 2805 3565 2813
rect 3578 2793 3581 2926
rect 3602 2823 3605 2936
rect 3610 2913 3613 2946
rect 3626 2903 3629 2956
rect 3634 2933 3637 2966
rect 3634 2913 3637 2926
rect 3642 2893 3645 3043
rect 3650 3003 3653 3026
rect 3658 3016 3661 3066
rect 3722 3033 3725 3173
rect 3762 3133 3765 3156
rect 3738 3113 3741 3126
rect 3778 3123 3781 3146
rect 3802 3143 3805 3336
rect 3826 3323 3829 3346
rect 3842 3313 3845 3406
rect 3858 3403 3861 3443
rect 3850 3246 3853 3346
rect 3866 3263 3869 3556
rect 3874 3543 3877 3606
rect 3882 3576 3885 3616
rect 3890 3593 3893 3606
rect 3882 3573 3889 3576
rect 3874 3523 3877 3536
rect 3886 3516 3889 3573
rect 3898 3523 3901 3686
rect 3906 3533 3909 3626
rect 3914 3526 3917 3616
rect 3906 3523 3917 3526
rect 3882 3513 3889 3516
rect 3874 3306 3877 3416
rect 3882 3403 3885 3513
rect 3906 3506 3909 3523
rect 3922 3516 3925 3716
rect 3930 3693 3933 3726
rect 3938 3656 3941 3736
rect 3954 3733 3957 3756
rect 3962 3733 3965 3783
rect 3946 3663 3949 3726
rect 3962 3693 3965 3726
rect 3970 3683 3973 3776
rect 4002 3773 4005 3833
rect 4010 3813 4013 3863
rect 4042 3796 4045 3956
rect 4066 3933 4069 3956
rect 4114 3933 4117 4016
rect 4050 3806 4053 3816
rect 4058 3813 4061 3826
rect 4082 3813 4085 3836
rect 4050 3803 4069 3806
rect 4010 3736 4013 3796
rect 4042 3793 4053 3796
rect 3938 3653 3949 3656
rect 3930 3623 3933 3636
rect 3946 3613 3949 3653
rect 3962 3623 3965 3636
rect 3930 3523 3933 3606
rect 3938 3533 3941 3546
rect 3898 3503 3909 3506
rect 3898 3376 3901 3503
rect 3914 3383 3917 3516
rect 3922 3513 3933 3516
rect 3898 3373 3909 3376
rect 3922 3373 3925 3506
rect 3930 3413 3933 3513
rect 3938 3503 3941 3526
rect 3946 3426 3949 3556
rect 3954 3533 3957 3606
rect 3962 3603 3965 3616
rect 3978 3613 3981 3736
rect 3986 3733 3997 3736
rect 4002 3733 4013 3736
rect 4018 3733 4021 3746
rect 3994 3726 3997 3733
rect 3986 3713 3989 3726
rect 3994 3723 4005 3726
rect 4002 3713 4005 3723
rect 3986 3566 3989 3606
rect 3994 3603 3997 3706
rect 4010 3673 4013 3733
rect 4026 3656 4029 3776
rect 4034 3733 4037 3786
rect 4050 3733 4053 3793
rect 4074 3763 4077 3806
rect 4090 3803 4093 3926
rect 4146 3876 4149 3926
rect 4138 3873 4149 3876
rect 4138 3826 4141 3873
rect 4138 3823 4149 3826
rect 4098 3756 4101 3816
rect 4106 3793 4109 3806
rect 4146 3803 4149 3823
rect 4090 3753 4101 3756
rect 4074 3723 4077 3746
rect 4130 3733 4149 3736
rect 4130 3723 4133 3733
rect 4138 3713 4141 3726
rect 4026 3653 4045 3656
rect 4002 3573 4005 3616
rect 4010 3613 4013 3626
rect 3986 3563 4005 3566
rect 3962 3533 3965 3546
rect 3978 3533 3981 3546
rect 3986 3533 3989 3556
rect 3970 3446 3973 3526
rect 3938 3423 3949 3426
rect 3962 3443 3973 3446
rect 3882 3333 3901 3336
rect 3882 3323 3885 3333
rect 3890 3313 3893 3326
rect 3898 3306 3901 3326
rect 3874 3303 3881 3306
rect 3842 3243 3853 3246
rect 3818 3193 3821 3216
rect 3842 3183 3845 3243
rect 3878 3236 3881 3303
rect 3890 3303 3901 3306
rect 3878 3233 3885 3236
rect 3866 3186 3869 3206
rect 3882 3203 3885 3233
rect 3890 3203 3893 3303
rect 3906 3223 3909 3373
rect 3922 3343 3933 3346
rect 3938 3343 3941 3423
rect 3930 3336 3933 3343
rect 3914 3313 3917 3326
rect 3898 3213 3909 3216
rect 3914 3213 3917 3246
rect 3922 3233 3925 3336
rect 3930 3333 3941 3336
rect 3930 3303 3933 3326
rect 3922 3213 3933 3216
rect 3938 3213 3941 3326
rect 3946 3313 3949 3416
rect 3962 3406 3965 3443
rect 3970 3413 3973 3436
rect 3954 3396 3957 3406
rect 3962 3403 3973 3406
rect 3978 3403 3981 3526
rect 3986 3433 3989 3526
rect 3994 3516 3997 3536
rect 4002 3533 4005 3563
rect 4010 3533 4013 3606
rect 4026 3596 4029 3616
rect 4018 3593 4029 3596
rect 4034 3593 4037 3606
rect 4018 3526 4021 3593
rect 4042 3553 4045 3653
rect 4050 3563 4053 3626
rect 4066 3576 4069 3646
rect 4090 3593 4093 3616
rect 4066 3573 4093 3576
rect 4034 3533 4037 3546
rect 3994 3513 4001 3516
rect 3986 3413 3989 3426
rect 3998 3416 4001 3513
rect 4010 3423 4013 3526
rect 4018 3523 4029 3526
rect 4050 3523 4053 3536
rect 3998 3413 4013 3416
rect 4034 3413 4037 3426
rect 3954 3393 3965 3396
rect 3954 3323 3957 3376
rect 3962 3333 3965 3393
rect 3970 3323 3973 3403
rect 3994 3336 3997 3406
rect 3978 3333 3997 3336
rect 3986 3313 3989 3326
rect 4002 3273 4005 3336
rect 4010 3333 4013 3413
rect 4042 3403 4045 3506
rect 4074 3503 4077 3526
rect 4082 3496 4085 3566
rect 4074 3493 4085 3496
rect 4050 3413 4061 3416
rect 4018 3323 4021 3366
rect 4026 3333 4029 3346
rect 4042 3333 4045 3356
rect 4050 3326 4053 3406
rect 4058 3353 4061 3406
rect 4066 3363 4069 3416
rect 4074 3393 4077 3493
rect 4090 3426 4093 3573
rect 4114 3536 4117 3556
rect 4114 3533 4121 3536
rect 4118 3486 4121 3533
rect 4114 3483 4121 3486
rect 4114 3436 4117 3483
rect 4114 3433 4121 3436
rect 4082 3413 4085 3426
rect 4090 3423 4109 3426
rect 4090 3363 4093 3406
rect 4034 3293 4037 3326
rect 4042 3323 4053 3326
rect 4066 3323 4069 3336
rect 4090 3323 4093 3346
rect 3866 3183 3877 3186
rect 3794 3133 3813 3136
rect 3842 3133 3853 3136
rect 3658 3013 3669 3016
rect 3658 2993 3661 3006
rect 3666 2966 3669 3013
rect 3674 3003 3677 3016
rect 3770 3013 3773 3036
rect 3778 3016 3781 3116
rect 3794 3113 3797 3126
rect 3802 3073 3805 3116
rect 3810 3103 3813 3133
rect 3818 3113 3821 3126
rect 3826 3123 3837 3126
rect 3826 3113 3829 3123
rect 3842 3113 3845 3126
rect 3858 3113 3861 3136
rect 3874 3133 3877 3183
rect 3778 3013 3789 3016
rect 3770 3003 3781 3006
rect 3786 3003 3789 3013
rect 3650 2963 3669 2966
rect 3650 2913 3653 2963
rect 3674 2956 3677 2996
rect 3658 2943 3661 2956
rect 3666 2953 3677 2956
rect 3658 2923 3661 2936
rect 3666 2846 3669 2953
rect 3674 2933 3685 2936
rect 3698 2933 3701 2956
rect 3714 2933 3717 2996
rect 3746 2943 3749 2956
rect 3754 2936 3757 2976
rect 3762 2946 3765 2996
rect 3762 2943 3773 2946
rect 3674 2923 3693 2926
rect 3706 2903 3709 2926
rect 3714 2893 3717 2926
rect 3658 2843 3669 2846
rect 3594 2813 3605 2816
rect 3514 2763 3517 2783
rect 3602 2743 3605 2786
rect 3610 2743 3613 2806
rect 3618 2803 3637 2806
rect 3642 2753 3645 2816
rect 3514 2713 3517 2726
rect 3642 2713 3645 2736
rect 3650 2723 3653 2816
rect 3658 2766 3661 2843
rect 3666 2823 3669 2836
rect 3666 2783 3669 2806
rect 3674 2803 3677 2826
rect 3698 2813 3701 2836
rect 3722 2813 3725 2936
rect 3754 2933 3765 2936
rect 3770 2923 3773 2943
rect 3786 2936 3789 2996
rect 3778 2906 3781 2936
rect 3786 2933 3797 2936
rect 3786 2913 3789 2926
rect 3794 2923 3797 2933
rect 3770 2903 3781 2906
rect 3794 2903 3797 2916
rect 3802 2913 3805 2996
rect 3810 2933 3813 2976
rect 3858 2956 3861 3016
rect 3874 3003 3877 3016
rect 3858 2953 3865 2956
rect 3826 2936 3829 2946
rect 3842 2943 3853 2946
rect 3818 2933 3829 2936
rect 3674 2773 3677 2796
rect 3658 2763 3677 2766
rect 3410 2553 3413 2606
rect 3418 2566 3421 2616
rect 3426 2613 3429 2626
rect 3522 2616 3525 2706
rect 3514 2613 3525 2616
rect 3418 2563 3445 2566
rect 3322 2533 3333 2536
rect 3378 2533 3381 2546
rect 3322 2483 3325 2533
rect 3306 2433 3309 2483
rect 3330 2473 3333 2526
rect 3258 2423 3277 2426
rect 3258 2413 3261 2423
rect 3250 2405 3261 2408
rect 3242 2393 3261 2396
rect 3226 2323 3229 2393
rect 3170 2313 3181 2316
rect 3170 2293 3173 2313
rect 3122 2253 3141 2256
rect 3090 2243 3101 2246
rect 3090 2176 3093 2243
rect 3098 2183 3101 2206
rect 3114 2193 3117 2206
rect 3138 2176 3141 2253
rect 3258 2226 3261 2393
rect 3266 2333 3269 2416
rect 3274 2413 3277 2423
rect 3306 2333 3309 2416
rect 3362 2393 3365 2406
rect 3370 2403 3373 2426
rect 3378 2413 3381 2526
rect 3394 2523 3397 2536
rect 3322 2323 3325 2336
rect 3354 2233 3357 2246
rect 3362 2226 3365 2326
rect 3378 2323 3381 2406
rect 3386 2403 3389 2496
rect 3394 2413 3397 2516
rect 3402 2403 3405 2526
rect 3410 2523 3413 2546
rect 3418 2513 3421 2536
rect 3426 2523 3429 2536
rect 3434 2523 3437 2556
rect 3410 2413 3413 2476
rect 3418 2413 3421 2446
rect 3442 2433 3445 2563
rect 3474 2433 3477 2586
rect 3498 2563 3501 2596
rect 3514 2593 3517 2613
rect 3530 2603 3533 2626
rect 3538 2613 3541 2696
rect 3546 2573 3549 2606
rect 3554 2586 3557 2616
rect 3562 2613 3565 2626
rect 3658 2616 3661 2746
rect 3666 2723 3669 2736
rect 3674 2733 3677 2763
rect 3682 2703 3685 2806
rect 3738 2803 3741 2846
rect 3770 2836 3773 2903
rect 3818 2896 3821 2933
rect 3826 2903 3829 2926
rect 3770 2833 3781 2836
rect 3778 2816 3781 2833
rect 3706 2783 3709 2796
rect 3754 2793 3757 2816
rect 3762 2813 3781 2816
rect 3794 2813 3797 2896
rect 3818 2893 3829 2896
rect 3762 2803 3781 2806
rect 3762 2783 3765 2796
rect 3778 2743 3781 2796
rect 3802 2743 3805 2806
rect 3810 2743 3813 2826
rect 3826 2803 3829 2893
rect 3834 2813 3837 2926
rect 3842 2823 3845 2936
rect 3850 2803 3853 2926
rect 3862 2796 3865 2953
rect 3874 2803 3877 2966
rect 3882 2923 3885 3086
rect 3890 2923 3893 3096
rect 3898 2816 3901 3206
rect 3906 3123 3909 3206
rect 3922 3183 3925 3206
rect 3946 3196 3949 3226
rect 4002 3213 4005 3236
rect 3942 3193 3949 3196
rect 3942 3126 3945 3193
rect 3942 3123 3949 3126
rect 3954 3123 3957 3206
rect 3978 3193 3981 3206
rect 3970 3133 3973 3156
rect 3994 3123 3997 3136
rect 3906 2993 3909 3106
rect 3946 3103 3949 3123
rect 4018 3106 4021 3126
rect 4010 3103 4021 3106
rect 4010 3046 4013 3103
rect 4010 3043 4021 3046
rect 3922 3013 3925 3026
rect 3922 2943 3933 2946
rect 3906 2923 3909 2936
rect 3922 2856 3925 2943
rect 3882 2813 3901 2816
rect 3906 2853 3925 2856
rect 3938 2853 3941 2996
rect 3962 2933 3973 2936
rect 3858 2793 3865 2796
rect 3906 2793 3909 2853
rect 3930 2833 3941 2836
rect 3922 2813 3925 2826
rect 3938 2823 3941 2833
rect 3690 2723 3693 2736
rect 3786 2733 3797 2736
rect 3802 2726 3805 2736
rect 3858 2733 3861 2793
rect 3906 2733 3909 2746
rect 3914 2733 3917 2756
rect 3938 2743 3941 2806
rect 3946 2803 3949 2926
rect 3954 2823 3957 2926
rect 3962 2923 3965 2933
rect 3970 2913 3973 2926
rect 3970 2823 3973 2836
rect 3978 2823 3981 2986
rect 3994 2933 3997 2956
rect 3986 2833 3989 2926
rect 4010 2923 4013 2996
rect 4018 2983 4021 3043
rect 4026 3033 4029 3086
rect 4026 3003 4029 3026
rect 4034 3013 4037 3116
rect 3954 2813 3965 2816
rect 3978 2743 3981 2806
rect 3922 2733 3941 2736
rect 3794 2723 3805 2726
rect 3794 2706 3797 2723
rect 3730 2686 3733 2706
rect 3730 2683 3741 2686
rect 3650 2613 3661 2616
rect 3650 2593 3653 2613
rect 3682 2603 3685 2626
rect 3722 2613 3725 2676
rect 3738 2606 3741 2683
rect 3698 2593 3701 2606
rect 3730 2603 3741 2606
rect 3770 2603 3773 2686
rect 3554 2583 3573 2586
rect 3514 2533 3517 2566
rect 3490 2513 3493 2526
rect 3530 2426 3533 2526
rect 3538 2463 3541 2536
rect 3554 2533 3557 2546
rect 3538 2433 3541 2446
rect 3546 2426 3549 2506
rect 3554 2433 3557 2526
rect 3562 2523 3565 2576
rect 3570 2566 3573 2583
rect 3570 2563 3577 2566
rect 3410 2333 3413 2356
rect 3258 2223 3269 2226
rect 3346 2223 3365 2226
rect 3090 2173 3109 2176
rect 3074 2133 3081 2136
rect 3074 2093 3077 2133
rect 3082 2016 3085 2126
rect 3090 2113 3093 2136
rect 3074 2013 3085 2016
rect 3066 1923 3069 1946
rect 3074 1913 3077 2013
rect 3082 1966 3085 2006
rect 3090 1983 3093 2036
rect 3098 2013 3101 2126
rect 3106 1993 3109 2173
rect 3114 2173 3141 2176
rect 3114 2123 3117 2173
rect 3122 2123 3125 2136
rect 3130 2063 3133 2166
rect 3146 2133 3149 2216
rect 3194 2143 3205 2146
rect 3194 2136 3197 2143
rect 3138 2113 3141 2126
rect 3154 2043 3157 2136
rect 3162 2133 3197 2136
rect 3114 2013 3117 2036
rect 3082 1963 3089 1966
rect 3086 1906 3089 1963
rect 3082 1903 3089 1906
rect 2970 1713 2981 1716
rect 3018 1713 3021 1726
rect 2970 1606 2973 1713
rect 2962 1603 2973 1606
rect 2962 1566 2965 1603
rect 2986 1576 2989 1636
rect 2994 1603 2997 1676
rect 3026 1656 3029 1736
rect 3034 1673 3037 1726
rect 3050 1713 3053 1726
rect 3010 1603 3013 1656
rect 3026 1653 3037 1656
rect 3058 1653 3061 1876
rect 3082 1846 3085 1903
rect 3114 1853 3117 1946
rect 3130 1896 3133 2026
rect 3138 2003 3141 2026
rect 3146 2013 3149 2026
rect 3162 1996 3165 2133
rect 3138 1913 3141 1996
rect 3154 1993 3165 1996
rect 3170 2123 3181 2126
rect 3154 1926 3157 1993
rect 3154 1923 3165 1926
rect 3126 1893 3133 1896
rect 3082 1843 3089 1846
rect 3086 1796 3089 1843
rect 3082 1793 3089 1796
rect 3074 1733 3077 1746
rect 3082 1716 3085 1793
rect 3078 1713 3085 1716
rect 3034 1613 3037 1653
rect 3078 1626 3081 1713
rect 3078 1623 3085 1626
rect 2986 1573 2997 1576
rect 2958 1563 2965 1566
rect 2958 1486 2961 1563
rect 2978 1546 2981 1566
rect 2978 1543 2985 1546
rect 2982 1486 2985 1543
rect 2958 1483 2965 1486
rect 2938 1393 2941 1416
rect 2946 1366 2949 1416
rect 2926 1363 2949 1366
rect 2898 1333 2905 1336
rect 2866 1323 2877 1326
rect 2826 1283 2833 1286
rect 2810 1273 2821 1276
rect 2802 1263 2813 1266
rect 2802 1213 2805 1226
rect 2754 1143 2765 1146
rect 2754 1023 2757 1143
rect 2762 1053 2765 1126
rect 2778 1093 2781 1206
rect 2794 1193 2797 1206
rect 2810 1193 2813 1263
rect 2818 1203 2821 1273
rect 2830 1196 2833 1283
rect 2842 1213 2845 1316
rect 2854 1313 2869 1316
rect 2866 1236 2869 1313
rect 2866 1233 2877 1236
rect 2826 1193 2833 1196
rect 2818 1133 2821 1146
rect 2786 1113 2789 1126
rect 2762 973 2765 1016
rect 2770 1003 2773 1016
rect 2778 1013 2781 1026
rect 2778 956 2781 996
rect 2786 963 2789 1106
rect 2810 1103 2813 1116
rect 2794 983 2797 1016
rect 2802 966 2805 1016
rect 2810 1003 2813 1096
rect 2818 1023 2821 1126
rect 2826 1016 2829 1193
rect 2834 1103 2837 1126
rect 2818 1013 2829 1016
rect 2834 1013 2837 1096
rect 2842 1013 2845 1206
rect 2858 1146 2861 1216
rect 2866 1203 2869 1216
rect 2874 1213 2877 1233
rect 2882 1203 2885 1226
rect 2890 1213 2893 1326
rect 2902 1226 2905 1333
rect 2898 1223 2905 1226
rect 2890 1186 2893 1206
rect 2886 1183 2893 1186
rect 2850 1133 2853 1146
rect 2858 1143 2877 1146
rect 2850 1103 2853 1126
rect 2858 1093 2861 1136
rect 2866 1036 2869 1126
rect 2874 1103 2877 1143
rect 2886 1086 2889 1183
rect 2898 1113 2901 1223
rect 2906 1103 2909 1206
rect 2914 1176 2917 1336
rect 2926 1246 2929 1363
rect 2922 1243 2929 1246
rect 2922 1186 2925 1243
rect 2938 1203 2941 1356
rect 2946 1303 2949 1346
rect 2954 1323 2957 1436
rect 2962 1343 2965 1483
rect 2978 1483 2985 1486
rect 2978 1456 2981 1483
rect 2978 1453 2985 1456
rect 2982 1376 2985 1453
rect 2978 1373 2985 1376
rect 2962 1213 2965 1336
rect 2978 1333 2981 1373
rect 2970 1213 2973 1326
rect 2986 1323 2989 1336
rect 2994 1316 2997 1573
rect 2978 1313 2997 1316
rect 2922 1183 2933 1186
rect 2914 1173 2925 1176
rect 2914 1093 2917 1126
rect 2922 1086 2925 1173
rect 2930 1123 2933 1183
rect 2978 1163 2981 1313
rect 2946 1113 2949 1126
rect 2886 1083 2893 1086
rect 2890 1066 2893 1083
rect 2914 1083 2925 1086
rect 2890 1063 2909 1066
rect 2850 1033 2869 1036
rect 2818 993 2821 1013
rect 2826 1003 2837 1006
rect 2802 963 2813 966
rect 2778 953 2805 956
rect 2754 933 2765 936
rect 2706 833 2709 846
rect 2714 813 2717 826
rect 2722 823 2725 856
rect 2730 823 2733 926
rect 2746 883 2749 926
rect 2762 853 2765 926
rect 2770 836 2773 946
rect 2778 943 2797 946
rect 2802 943 2805 953
rect 2778 933 2781 943
rect 2778 873 2781 926
rect 2786 923 2789 936
rect 2794 913 2797 943
rect 2738 813 2741 836
rect 2754 833 2773 836
rect 2690 703 2693 726
rect 2706 723 2709 786
rect 2722 723 2725 736
rect 2674 693 2685 696
rect 2634 593 2645 596
rect 2618 533 2621 566
rect 2634 536 2637 593
rect 2658 586 2661 626
rect 2682 603 2685 693
rect 2690 613 2693 626
rect 2626 533 2637 536
rect 2642 583 2661 586
rect 2642 533 2645 583
rect 2666 543 2693 546
rect 2618 513 2621 526
rect 2626 393 2629 533
rect 2650 413 2653 536
rect 2666 533 2669 543
rect 2658 436 2661 526
rect 2658 433 2669 436
rect 2650 393 2653 406
rect 2666 366 2669 433
rect 2586 333 2589 346
rect 2594 333 2597 366
rect 2658 363 2669 366
rect 2602 343 2629 346
rect 2570 303 2573 326
rect 2602 296 2605 336
rect 2594 293 2605 296
rect 2562 196 2565 216
rect 2570 213 2581 216
rect 2586 213 2589 226
rect 2594 203 2597 293
rect 2610 213 2613 336
rect 2626 333 2629 343
rect 2618 263 2621 326
rect 2634 323 2637 336
rect 2562 193 2573 196
rect 2570 123 2573 193
rect 2610 166 2613 206
rect 2618 176 2621 206
rect 2626 196 2629 216
rect 2634 203 2637 236
rect 2642 223 2645 336
rect 2642 196 2645 206
rect 2626 193 2645 196
rect 2650 176 2653 336
rect 2658 303 2661 363
rect 2666 333 2669 356
rect 2674 306 2677 526
rect 2682 476 2685 536
rect 2690 486 2693 536
rect 2698 533 2701 676
rect 2706 593 2709 646
rect 2722 576 2725 686
rect 2730 663 2733 806
rect 2738 653 2741 756
rect 2746 733 2749 806
rect 2754 743 2757 833
rect 2762 803 2765 826
rect 2802 813 2805 936
rect 2810 893 2813 963
rect 2826 933 2829 946
rect 2818 913 2821 926
rect 2778 753 2781 806
rect 2762 586 2765 666
rect 2770 643 2773 746
rect 2786 733 2789 776
rect 2770 613 2773 626
rect 2722 573 2733 576
rect 2706 523 2709 546
rect 2714 513 2717 526
rect 2730 496 2733 573
rect 2730 493 2741 496
rect 2690 483 2709 486
rect 2682 473 2693 476
rect 2682 413 2685 436
rect 2670 303 2677 306
rect 2658 193 2661 236
rect 2618 173 2653 176
rect 2670 176 2673 303
rect 2682 233 2685 406
rect 2690 366 2693 473
rect 2698 396 2701 416
rect 2706 403 2709 483
rect 2714 396 2717 406
rect 2698 393 2717 396
rect 2690 363 2701 366
rect 2690 333 2693 346
rect 2698 316 2701 363
rect 2714 333 2717 346
rect 2694 313 2701 316
rect 2694 236 2697 313
rect 2694 233 2701 236
rect 2670 173 2677 176
rect 2610 163 2629 166
rect 2626 123 2629 163
rect 2634 123 2637 173
rect 2674 153 2677 173
rect 2682 123 2685 216
rect 2690 203 2693 216
rect 2698 146 2701 233
rect 2706 213 2709 326
rect 2722 236 2725 476
rect 2730 333 2733 416
rect 2738 403 2741 493
rect 2746 396 2749 576
rect 2754 473 2757 586
rect 2762 583 2769 586
rect 2766 496 2769 583
rect 2762 493 2769 496
rect 2738 393 2749 396
rect 2738 333 2741 393
rect 2746 343 2749 356
rect 2730 323 2741 326
rect 2754 323 2757 416
rect 2762 403 2765 493
rect 2770 383 2773 476
rect 2778 413 2781 526
rect 2786 473 2789 726
rect 2794 663 2797 736
rect 2802 723 2805 806
rect 2810 773 2813 886
rect 2834 883 2837 976
rect 2842 906 2845 1006
rect 2850 923 2853 1033
rect 2858 973 2861 1016
rect 2874 1003 2877 1046
rect 2842 903 2849 906
rect 2802 676 2805 706
rect 2810 696 2813 736
rect 2818 723 2821 876
rect 2826 703 2829 846
rect 2846 786 2849 903
rect 2858 813 2861 936
rect 2842 783 2849 786
rect 2842 763 2845 783
rect 2842 733 2845 746
rect 2810 693 2821 696
rect 2802 673 2809 676
rect 2794 406 2797 656
rect 2806 586 2809 673
rect 2818 613 2821 693
rect 2802 583 2809 586
rect 2802 423 2805 583
rect 2810 533 2813 566
rect 2810 496 2813 526
rect 2818 513 2821 526
rect 2826 523 2829 656
rect 2834 613 2837 646
rect 2842 603 2845 626
rect 2866 616 2869 896
rect 2874 703 2877 986
rect 2890 976 2893 996
rect 2882 973 2893 976
rect 2882 843 2885 973
rect 2898 923 2901 1006
rect 2906 873 2909 1063
rect 2914 983 2917 1083
rect 2938 1056 2941 1086
rect 2938 1053 2949 1056
rect 2922 1003 2925 1016
rect 2946 976 2949 1053
rect 2962 983 2965 1136
rect 2970 1113 2973 1126
rect 2914 973 2949 976
rect 2890 813 2893 826
rect 2882 783 2885 806
rect 2914 803 2917 973
rect 2922 863 2925 946
rect 2946 856 2949 936
rect 2922 853 2949 856
rect 2882 653 2885 766
rect 2890 723 2893 776
rect 2906 686 2909 726
rect 2898 683 2909 686
rect 2922 683 2925 853
rect 2970 816 2973 1036
rect 2978 923 2981 1136
rect 2986 1076 2989 1306
rect 2994 1083 2997 1166
rect 3002 1123 3005 1216
rect 3010 1203 3013 1596
rect 3042 1533 3053 1536
rect 3074 1533 3077 1606
rect 3018 1503 3021 1526
rect 3026 1493 3029 1516
rect 3050 1503 3053 1533
rect 3018 1413 3021 1426
rect 3034 1403 3037 1416
rect 3034 1333 3037 1396
rect 3042 1323 3045 1346
rect 3050 1333 3053 1376
rect 3058 1313 3061 1516
rect 3066 1393 3069 1416
rect 3066 1226 3069 1336
rect 3074 1323 3077 1516
rect 3082 1513 3085 1623
rect 3090 1603 3093 1736
rect 3098 1716 3101 1836
rect 3106 1733 3109 1816
rect 3126 1766 3129 1893
rect 3126 1763 3133 1766
rect 3122 1733 3125 1746
rect 3130 1743 3133 1763
rect 3114 1723 3133 1726
rect 3098 1713 3105 1716
rect 3102 1596 3105 1713
rect 3114 1613 3117 1676
rect 3098 1593 3105 1596
rect 3098 1546 3101 1593
rect 3090 1503 3093 1546
rect 3098 1543 3109 1546
rect 3098 1413 3101 1536
rect 3082 1333 3085 1356
rect 3090 1333 3093 1346
rect 3106 1336 3109 1543
rect 3114 1423 3117 1606
rect 3122 1586 3125 1716
rect 3130 1603 3133 1723
rect 3138 1713 3141 1906
rect 3154 1883 3157 1906
rect 3138 1613 3141 1636
rect 3146 1593 3149 1876
rect 3162 1833 3165 1923
rect 3154 1733 3157 1816
rect 3162 1753 3165 1816
rect 3162 1716 3165 1746
rect 3158 1713 3165 1716
rect 3158 1636 3161 1713
rect 3158 1633 3165 1636
rect 3122 1583 3149 1586
rect 3122 1523 3125 1576
rect 3138 1523 3141 1536
rect 3146 1533 3149 1583
rect 3154 1543 3157 1616
rect 3102 1333 3109 1336
rect 3122 1336 3125 1516
rect 3146 1473 3149 1526
rect 3154 1513 3157 1536
rect 3162 1523 3165 1633
rect 3170 1466 3173 2123
rect 3178 2023 3181 2116
rect 3202 2113 3205 2136
rect 3210 2113 3213 2216
rect 3226 2193 3229 2206
rect 3250 2176 3253 2216
rect 3234 2173 3253 2176
rect 3234 2133 3237 2173
rect 3266 2156 3269 2223
rect 3258 2153 3269 2156
rect 3250 2133 3253 2146
rect 3258 2133 3261 2153
rect 3218 2116 3221 2126
rect 3234 2123 3245 2126
rect 3218 2113 3229 2116
rect 3258 2113 3261 2126
rect 3186 2103 3197 2106
rect 3186 1916 3189 2096
rect 3218 2073 3221 2113
rect 3266 2056 3269 2136
rect 3298 2133 3301 2146
rect 3306 2133 3317 2136
rect 3306 2123 3325 2126
rect 3330 2123 3333 2216
rect 3362 2186 3365 2206
rect 3354 2183 3365 2186
rect 3242 2053 3269 2056
rect 3202 2013 3213 2016
rect 3202 1933 3205 2013
rect 3210 1983 3213 2006
rect 3218 2003 3221 2016
rect 3226 2013 3229 2026
rect 3218 1933 3221 1946
rect 3178 1913 3189 1916
rect 3178 1573 3181 1913
rect 3186 1563 3189 1906
rect 3202 1883 3205 1916
rect 3242 1873 3245 2053
rect 3250 1986 3253 2016
rect 3258 2003 3261 2026
rect 3266 2013 3269 2046
rect 3266 1993 3269 2006
rect 3250 1983 3257 1986
rect 3254 1876 3257 1983
rect 3274 1963 3277 2016
rect 3290 2013 3293 2026
rect 3282 2003 3293 2006
rect 3298 1993 3301 2066
rect 3306 2013 3309 2123
rect 3354 2066 3357 2183
rect 3370 2166 3373 2226
rect 3386 2183 3389 2326
rect 3426 2323 3429 2416
rect 3434 2413 3437 2426
rect 3530 2423 3541 2426
rect 3546 2423 3557 2426
rect 3458 2306 3461 2416
rect 3474 2386 3477 2406
rect 3522 2393 3525 2416
rect 3530 2413 3549 2416
rect 3554 2413 3557 2423
rect 3530 2403 3533 2413
rect 3470 2383 3477 2386
rect 3470 2326 3473 2383
rect 3470 2323 3477 2326
rect 3458 2303 3465 2306
rect 3434 2193 3437 2216
rect 3450 2206 3453 2286
rect 3462 2246 3465 2303
rect 3474 2283 3477 2323
rect 3458 2243 3465 2246
rect 3458 2226 3461 2243
rect 3482 2233 3485 2366
rect 3506 2283 3509 2356
rect 3530 2333 3533 2386
rect 3458 2223 3477 2226
rect 3450 2203 3457 2206
rect 3366 2163 3373 2166
rect 3366 2086 3369 2163
rect 3386 2123 3389 2146
rect 3434 2133 3437 2186
rect 3454 2106 3457 2203
rect 3466 2133 3469 2216
rect 3490 2146 3493 2206
rect 3474 2143 3493 2146
rect 3450 2103 3457 2106
rect 3366 2083 3373 2086
rect 3354 2063 3365 2066
rect 3266 1923 3269 1946
rect 3250 1873 3257 1876
rect 3250 1853 3253 1873
rect 3202 1816 3205 1836
rect 3202 1813 3213 1816
rect 3210 1766 3213 1813
rect 3202 1763 3213 1766
rect 3194 1733 3197 1756
rect 3202 1656 3205 1763
rect 3218 1726 3221 1746
rect 3194 1653 3205 1656
rect 3214 1723 3221 1726
rect 3214 1656 3217 1723
rect 3214 1653 3221 1656
rect 3194 1573 3197 1653
rect 3210 1613 3213 1636
rect 3218 1613 3221 1653
rect 3202 1593 3205 1606
rect 3210 1603 3221 1606
rect 3226 1603 3229 1816
rect 3250 1803 3253 1836
rect 3266 1823 3269 1886
rect 3274 1786 3277 1856
rect 3282 1833 3285 1986
rect 3330 1983 3333 2006
rect 3354 2003 3357 2016
rect 3290 1816 3293 1916
rect 3306 1903 3317 1906
rect 3258 1783 3277 1786
rect 3286 1813 3293 1816
rect 3298 1813 3301 1836
rect 3306 1813 3309 1903
rect 3322 1886 3325 1956
rect 3330 1946 3333 1966
rect 3330 1943 3337 1946
rect 3318 1883 3325 1886
rect 3234 1593 3237 1726
rect 3178 1533 3181 1556
rect 3178 1493 3181 1526
rect 3162 1463 3173 1466
rect 3130 1343 3133 1416
rect 3138 1413 3141 1436
rect 3146 1343 3149 1426
rect 3122 1333 3133 1336
rect 3102 1246 3105 1333
rect 3114 1253 3117 1326
rect 3130 1323 3133 1333
rect 3146 1313 3149 1326
rect 3154 1283 3157 1416
rect 3162 1323 3165 1463
rect 3186 1456 3189 1536
rect 3202 1533 3205 1546
rect 3170 1453 3189 1456
rect 3102 1243 3109 1246
rect 3066 1223 3077 1226
rect 3018 1133 3021 1216
rect 2986 1073 2997 1076
rect 2986 933 2989 1006
rect 2994 1003 2997 1073
rect 3002 933 3005 1006
rect 3010 993 3013 1016
rect 3018 1003 3021 1026
rect 3026 1013 3029 1146
rect 3050 1066 3053 1136
rect 3066 1133 3069 1216
rect 3074 1206 3077 1223
rect 3074 1203 3081 1206
rect 3078 1146 3081 1203
rect 3106 1176 3109 1243
rect 3074 1143 3081 1146
rect 3090 1173 3109 1176
rect 3074 1123 3077 1143
rect 3042 1063 3053 1066
rect 3034 986 3037 1056
rect 3042 1013 3045 1063
rect 3074 1013 3077 1026
rect 2930 813 2949 816
rect 2930 803 2933 813
rect 2938 746 2941 806
rect 2946 766 2949 813
rect 2954 773 2957 806
rect 2946 763 2957 766
rect 2934 743 2941 746
rect 2898 626 2901 683
rect 2934 646 2937 743
rect 2934 643 2941 646
rect 2890 623 2901 626
rect 2866 613 2877 616
rect 2850 603 2861 606
rect 2834 526 2837 536
rect 2834 523 2853 526
rect 2810 493 2821 496
rect 2794 403 2805 406
rect 2818 396 2821 493
rect 2858 446 2861 556
rect 2866 523 2869 606
rect 2874 596 2877 613
rect 2874 593 2881 596
rect 2878 486 2881 593
rect 2890 576 2893 623
rect 2930 616 2933 626
rect 2890 573 2901 576
rect 2878 483 2893 486
rect 2834 433 2837 446
rect 2858 443 2869 446
rect 2842 413 2845 426
rect 2810 393 2821 396
rect 2810 346 2813 393
rect 2850 353 2853 426
rect 2866 403 2869 443
rect 2890 386 2893 483
rect 2722 233 2733 236
rect 2714 166 2717 216
rect 2722 193 2725 226
rect 2730 176 2733 233
rect 2738 203 2741 216
rect 2754 213 2757 226
rect 2762 213 2765 346
rect 2802 343 2813 346
rect 2786 323 2789 336
rect 2802 296 2805 343
rect 2802 293 2813 296
rect 2794 213 2797 226
rect 2810 203 2813 293
rect 2834 276 2837 346
rect 2858 333 2861 386
rect 2886 383 2893 386
rect 2886 296 2889 383
rect 2874 293 2889 296
rect 2898 293 2901 573
rect 2906 393 2909 616
rect 2914 613 2933 616
rect 2938 613 2941 643
rect 2946 613 2949 756
rect 2954 723 2957 763
rect 2962 753 2965 816
rect 2970 813 2981 816
rect 2970 756 2973 806
rect 2978 763 2981 813
rect 2986 803 2989 866
rect 2994 813 2997 926
rect 3010 853 3013 936
rect 2994 773 2997 806
rect 3002 786 3005 826
rect 3018 813 3021 986
rect 3034 983 3045 986
rect 3026 806 3029 966
rect 3034 813 3037 936
rect 3042 896 3045 983
rect 3050 913 3053 936
rect 3058 933 3069 936
rect 3074 933 3077 946
rect 3042 893 3053 896
rect 3050 876 3053 893
rect 3050 873 3057 876
rect 3010 803 3021 806
rect 3026 803 3037 806
rect 3002 783 3013 786
rect 2970 753 2997 756
rect 2970 733 2973 746
rect 2962 703 2965 726
rect 2922 603 2941 606
rect 2946 603 2957 606
rect 2914 453 2917 536
rect 2922 523 2925 603
rect 2914 413 2917 446
rect 2906 323 2909 346
rect 2938 323 2941 486
rect 2946 383 2949 596
rect 2970 536 2973 726
rect 2978 723 2981 736
rect 2986 623 2989 736
rect 2994 676 2997 753
rect 3002 683 3005 736
rect 2994 673 3005 676
rect 2994 613 2997 666
rect 3002 653 3005 673
rect 2986 583 2989 606
rect 3002 603 3005 626
rect 3010 546 3013 783
rect 3018 733 3021 756
rect 3026 726 3029 746
rect 3034 736 3037 803
rect 3042 773 3045 856
rect 3034 733 3045 736
rect 2954 403 2957 456
rect 2962 413 2965 536
rect 2970 533 2981 536
rect 2986 526 2989 546
rect 3002 543 3013 546
rect 2970 523 2989 526
rect 2994 443 2997 536
rect 2978 413 2981 426
rect 3002 413 3005 543
rect 3010 413 3013 536
rect 2954 393 2965 396
rect 2834 273 2845 276
rect 2730 173 2741 176
rect 2714 163 2733 166
rect 2690 143 2701 146
rect 2690 43 2693 143
rect 2714 123 2717 136
rect 2730 133 2733 163
rect 2738 23 2741 173
rect 2746 113 2749 126
rect 2754 123 2757 196
rect 2842 176 2845 273
rect 2874 213 2877 293
rect 2890 213 2909 216
rect 2930 213 2933 296
rect 2946 213 2949 356
rect 2962 333 2965 393
rect 2970 326 2973 396
rect 2986 383 2989 406
rect 3002 356 3005 406
rect 3010 393 3013 406
rect 3018 386 3021 726
rect 3026 723 3045 726
rect 3054 716 3057 873
rect 3066 723 3069 926
rect 3082 923 3085 996
rect 3090 916 3093 1173
rect 3114 1133 3117 1196
rect 3122 1173 3125 1216
rect 3146 1203 3149 1246
rect 3154 1133 3157 1176
rect 3130 1123 3149 1126
rect 3162 1123 3165 1236
rect 3170 1183 3173 1453
rect 3178 1416 3181 1426
rect 3194 1416 3197 1526
rect 3210 1506 3213 1526
rect 3206 1503 3213 1506
rect 3206 1436 3209 1503
rect 3218 1436 3221 1526
rect 3226 1453 3229 1576
rect 3242 1533 3245 1736
rect 3258 1733 3261 1783
rect 3274 1666 3277 1726
rect 3258 1663 3277 1666
rect 3250 1613 3253 1626
rect 3250 1583 3253 1606
rect 3206 1433 3213 1436
rect 3218 1433 3225 1436
rect 3178 1413 3189 1416
rect 3194 1413 3205 1416
rect 3178 1333 3181 1406
rect 3194 1373 3197 1406
rect 3210 1366 3213 1433
rect 3222 1376 3225 1433
rect 3194 1363 3213 1366
rect 3218 1373 3225 1376
rect 3170 1133 3173 1166
rect 3170 1046 3173 1126
rect 3178 1113 3181 1326
rect 3186 1216 3189 1346
rect 3194 1233 3197 1363
rect 3202 1306 3205 1336
rect 3218 1333 3221 1373
rect 3234 1353 3237 1426
rect 3242 1403 3245 1526
rect 3242 1323 3245 1336
rect 3202 1303 3213 1306
rect 3186 1213 3197 1216
rect 3210 1213 3213 1303
rect 3218 1286 3221 1316
rect 3250 1306 3253 1566
rect 3258 1456 3261 1663
rect 3266 1633 3269 1646
rect 3266 1476 3269 1616
rect 3274 1613 3277 1656
rect 3286 1646 3289 1813
rect 3318 1776 3321 1883
rect 3334 1876 3337 1943
rect 3346 1933 3349 1986
rect 3346 1916 3349 1926
rect 3354 1923 3357 1966
rect 3362 1953 3365 2063
rect 3370 2043 3373 2083
rect 3426 2013 3429 2026
rect 3434 2023 3437 2046
rect 3378 1946 3381 1996
rect 3402 1946 3405 1956
rect 3362 1933 3365 1946
rect 3378 1943 3405 1946
rect 3378 1933 3381 1943
rect 3386 1926 3389 1936
rect 3362 1923 3389 1926
rect 3362 1916 3365 1923
rect 3346 1913 3365 1916
rect 3394 1913 3397 1926
rect 3402 1906 3405 1943
rect 3418 1926 3421 1936
rect 3426 1933 3429 1946
rect 3298 1773 3321 1776
rect 3330 1873 3337 1876
rect 3386 1903 3405 1906
rect 3410 1903 3413 1926
rect 3418 1923 3429 1926
rect 3298 1706 3301 1773
rect 3306 1733 3317 1736
rect 3322 1723 3325 1766
rect 3330 1743 3333 1873
rect 3330 1723 3333 1736
rect 3298 1703 3309 1706
rect 3306 1656 3309 1703
rect 3338 1673 3341 1826
rect 3346 1803 3357 1806
rect 3346 1666 3349 1756
rect 3354 1716 3357 1803
rect 3362 1793 3365 1806
rect 3370 1733 3373 1816
rect 3354 1713 3365 1716
rect 3298 1653 3309 1656
rect 3338 1663 3349 1666
rect 3286 1643 3293 1646
rect 3282 1603 3285 1626
rect 3290 1613 3293 1643
rect 3298 1633 3301 1653
rect 3290 1573 3293 1606
rect 3282 1523 3285 1546
rect 3290 1506 3293 1536
rect 3286 1503 3293 1506
rect 3266 1473 3277 1476
rect 3258 1453 3265 1456
rect 3262 1396 3265 1453
rect 3246 1303 3253 1306
rect 3258 1393 3265 1396
rect 3218 1283 3225 1286
rect 3222 1226 3225 1283
rect 3222 1223 3229 1226
rect 3186 1156 3189 1206
rect 3194 1163 3197 1213
rect 3202 1203 3213 1206
rect 3218 1183 3221 1206
rect 3226 1173 3229 1223
rect 3234 1193 3237 1266
rect 3246 1236 3249 1303
rect 3242 1233 3249 1236
rect 3186 1153 3197 1156
rect 3170 1043 3177 1046
rect 3122 976 3125 1006
rect 3146 1003 3149 1016
rect 3174 996 3177 1043
rect 3082 913 3093 916
rect 3106 973 3125 976
rect 3170 993 3177 996
rect 3082 866 3085 913
rect 3106 896 3109 973
rect 3130 923 3133 936
rect 3074 863 3085 866
rect 3098 893 3109 896
rect 3050 713 3057 716
rect 3026 513 3029 706
rect 3034 603 3037 686
rect 3042 613 3045 646
rect 3042 513 3045 526
rect 3034 493 3037 506
rect 3050 486 3053 713
rect 3074 703 3077 863
rect 3098 836 3101 893
rect 3098 833 3109 836
rect 3090 803 3093 816
rect 3090 723 3093 746
rect 3058 636 3061 656
rect 3058 633 3069 636
rect 3066 546 3069 633
rect 3098 613 3101 626
rect 3106 606 3109 833
rect 3034 483 3053 486
rect 3058 543 3069 546
rect 3098 603 3109 606
rect 3026 413 3029 456
rect 2994 353 3005 356
rect 3010 383 3021 386
rect 2978 333 2981 346
rect 2954 323 2973 326
rect 2986 323 2989 336
rect 2994 276 2997 353
rect 2986 273 2997 276
rect 2962 213 2965 266
rect 2970 213 2973 226
rect 2866 193 2869 206
rect 2834 173 2845 176
rect 2834 133 2837 173
rect 2786 113 2789 126
rect 2858 123 2861 166
rect 2882 123 2885 206
rect 2890 203 2901 206
rect 2898 183 2901 203
rect 2914 163 2917 206
rect 2970 173 2973 206
rect 2978 203 2981 236
rect 2986 193 2989 273
rect 3002 233 3005 336
rect 3010 296 3013 383
rect 3018 333 3021 356
rect 3026 323 3029 346
rect 3034 303 3037 483
rect 3058 453 3061 543
rect 3098 533 3101 603
rect 3114 533 3117 886
rect 3170 876 3173 993
rect 3162 873 3173 876
rect 3154 813 3157 856
rect 3162 806 3165 873
rect 3178 836 3181 946
rect 3186 883 3189 1146
rect 3194 1133 3197 1153
rect 3242 1143 3245 1233
rect 3258 1213 3261 1393
rect 3274 1376 3277 1473
rect 3266 1373 3277 1376
rect 3266 1263 3269 1373
rect 3286 1316 3289 1503
rect 3298 1413 3301 1616
rect 3306 1593 3309 1606
rect 3306 1476 3309 1566
rect 3314 1553 3317 1616
rect 3322 1563 3325 1606
rect 3338 1603 3341 1663
rect 3362 1646 3365 1713
rect 3378 1653 3381 1726
rect 3362 1643 3381 1646
rect 3362 1593 3365 1616
rect 3330 1523 3333 1536
rect 3354 1513 3357 1526
rect 3306 1473 3317 1476
rect 3314 1416 3317 1473
rect 3306 1413 3317 1416
rect 3298 1323 3301 1406
rect 3306 1393 3309 1413
rect 3286 1313 3293 1316
rect 3330 1313 3333 1486
rect 3258 1153 3261 1206
rect 3282 1203 3285 1216
rect 3290 1196 3293 1313
rect 3338 1296 3341 1456
rect 3362 1416 3365 1536
rect 3370 1523 3373 1606
rect 3378 1483 3381 1643
rect 3386 1583 3389 1903
rect 3394 1733 3397 1786
rect 3402 1753 3405 1836
rect 3426 1793 3429 1816
rect 3418 1756 3421 1776
rect 3434 1763 3437 1976
rect 3442 1896 3445 2066
rect 3450 2026 3453 2103
rect 3458 2033 3461 2046
rect 3474 2036 3477 2143
rect 3482 2133 3493 2136
rect 3498 2133 3501 2226
rect 3522 2216 3525 2326
rect 3546 2323 3549 2413
rect 3562 2405 3565 2516
rect 3574 2476 3577 2563
rect 3570 2473 3577 2476
rect 3570 2323 3573 2473
rect 3578 2413 3581 2456
rect 3586 2403 3589 2436
rect 3594 2383 3597 2576
rect 3602 2546 3605 2566
rect 3602 2543 3609 2546
rect 3606 2456 3609 2543
rect 3642 2533 3645 2566
rect 3658 2533 3661 2546
rect 3706 2533 3709 2576
rect 3602 2453 3609 2456
rect 3602 2353 3605 2453
rect 3610 2413 3613 2426
rect 3618 2403 3621 2526
rect 3706 2513 3709 2526
rect 3722 2523 3725 2546
rect 3634 2413 3637 2456
rect 3642 2403 3645 2426
rect 3650 2396 3653 2416
rect 3658 2403 3661 2466
rect 3674 2413 3677 2426
rect 3682 2406 3685 2416
rect 3690 2413 3693 2496
rect 3674 2403 3685 2406
rect 3706 2405 3709 2436
rect 3634 2393 3653 2396
rect 3674 2393 3677 2403
rect 3634 2343 3637 2393
rect 3730 2373 3733 2603
rect 3738 2523 3741 2536
rect 3746 2513 3749 2526
rect 3754 2483 3757 2536
rect 3762 2493 3765 2526
rect 3770 2523 3773 2536
rect 3778 2523 3781 2616
rect 3786 2613 3789 2706
rect 3794 2703 3805 2706
rect 3802 2606 3805 2703
rect 3890 2633 3893 2726
rect 3898 2703 3901 2726
rect 3810 2613 3813 2626
rect 3786 2506 3789 2606
rect 3794 2583 3797 2606
rect 3802 2603 3813 2606
rect 3794 2533 3805 2536
rect 3778 2503 3789 2506
rect 3778 2456 3781 2503
rect 3778 2453 3789 2456
rect 3642 2333 3645 2346
rect 3658 2333 3661 2356
rect 3546 2233 3549 2316
rect 3706 2313 3709 2326
rect 3738 2323 3741 2396
rect 3754 2393 3757 2416
rect 3786 2413 3789 2453
rect 3794 2423 3797 2526
rect 3802 2503 3805 2516
rect 3810 2496 3813 2603
rect 3898 2593 3901 2616
rect 3906 2603 3909 2626
rect 3914 2613 3917 2726
rect 3922 2706 3925 2726
rect 3946 2723 3949 2736
rect 3994 2733 3997 2836
rect 4002 2813 4005 2826
rect 4010 2823 4013 2836
rect 4018 2816 4021 2936
rect 4026 2913 4029 2926
rect 4034 2896 4037 3006
rect 4042 2933 4045 3323
rect 4058 3213 4061 3276
rect 4066 3213 4069 3306
rect 4098 3303 4101 3416
rect 4106 3323 4109 3423
rect 4118 3376 4121 3433
rect 4114 3373 4121 3376
rect 4090 3223 4093 3256
rect 4114 3246 4117 3373
rect 4130 3313 4133 3526
rect 4106 3243 4117 3246
rect 4106 3213 4109 3243
rect 4050 3203 4069 3206
rect 4050 3123 4053 3203
rect 4066 3133 4069 3156
rect 4090 3113 4093 3126
rect 4138 3083 4141 3576
rect 4146 3526 4149 3616
rect 4146 3523 4153 3526
rect 4150 3376 4153 3523
rect 4150 3373 4157 3376
rect 4146 3323 4149 3366
rect 4154 3333 4157 3373
rect 4146 3123 4149 3206
rect 4050 3013 4053 3026
rect 4066 2983 4069 3016
rect 4138 3003 4149 3006
rect 4050 2933 4053 2946
rect 4042 2916 4045 2926
rect 4074 2923 4077 2936
rect 4042 2913 4069 2916
rect 4034 2893 4045 2896
rect 4010 2813 4021 2816
rect 3922 2703 3933 2706
rect 3930 2646 3933 2703
rect 3922 2643 3933 2646
rect 3914 2593 3917 2606
rect 3802 2493 3813 2496
rect 3762 2333 3765 2376
rect 3746 2306 3749 2326
rect 3770 2313 3773 2336
rect 3786 2313 3789 2406
rect 3794 2393 3797 2406
rect 3802 2316 3805 2493
rect 3810 2323 3813 2456
rect 3818 2403 3821 2476
rect 3826 2423 3829 2506
rect 3826 2403 3829 2416
rect 3834 2406 3837 2516
rect 3842 2413 3845 2526
rect 3858 2513 3861 2586
rect 3922 2556 3925 2643
rect 3954 2633 3957 2726
rect 4002 2643 4005 2736
rect 4010 2723 4013 2776
rect 4018 2726 4021 2756
rect 4026 2733 4029 2856
rect 4042 2793 4045 2893
rect 4058 2813 4061 2836
rect 4066 2823 4069 2846
rect 4090 2833 4093 2926
rect 4106 2913 4109 2986
rect 4138 2933 4141 2996
rect 4154 2916 4157 3266
rect 4146 2913 4157 2916
rect 4098 2886 4101 2906
rect 4098 2883 4109 2886
rect 4106 2826 4109 2883
rect 4074 2813 4077 2826
rect 4098 2823 4109 2826
rect 4050 2753 4053 2806
rect 4098 2773 4101 2823
rect 4130 2743 4133 2796
rect 4146 2756 4149 2913
rect 4146 2753 4157 2756
rect 4018 2723 4029 2726
rect 4026 2716 4029 2723
rect 4018 2703 4021 2716
rect 4026 2713 4037 2716
rect 4042 2713 4045 2726
rect 3930 2613 3933 2626
rect 4026 2616 4029 2636
rect 4018 2613 4029 2616
rect 4034 2616 4037 2713
rect 4138 2706 4141 2736
rect 4130 2703 4141 2706
rect 4034 2613 4045 2616
rect 3914 2553 3925 2556
rect 3834 2403 3845 2406
rect 3850 2403 3853 2486
rect 3866 2413 3869 2536
rect 3874 2413 3877 2526
rect 3882 2513 3885 2536
rect 3890 2523 3893 2536
rect 3898 2476 3901 2526
rect 3894 2473 3901 2476
rect 3894 2426 3897 2473
rect 3882 2413 3885 2426
rect 3894 2423 3901 2426
rect 3826 2333 3829 2396
rect 3834 2333 3837 2403
rect 3874 2383 3877 2406
rect 3882 2393 3885 2406
rect 3890 2393 3893 2406
rect 3898 2383 3901 2423
rect 3906 2403 3909 2466
rect 3914 2403 3917 2553
rect 3962 2533 3965 2596
rect 4018 2593 4021 2613
rect 4026 2603 4037 2606
rect 4042 2593 4045 2613
rect 3986 2543 4005 2546
rect 3938 2513 3941 2526
rect 3962 2513 3965 2526
rect 3970 2483 3973 2536
rect 3986 2523 3989 2543
rect 3994 2523 3997 2536
rect 4002 2533 4005 2543
rect 4026 2536 4029 2546
rect 4018 2533 4029 2536
rect 4010 2513 4013 2526
rect 4018 2523 4021 2533
rect 4026 2473 4029 2526
rect 4042 2463 4045 2536
rect 3922 2403 3925 2436
rect 4050 2416 4053 2526
rect 4058 2513 4061 2526
rect 3930 2396 3933 2416
rect 3930 2393 3941 2396
rect 3802 2313 3813 2316
rect 3842 2313 3845 2326
rect 3850 2323 3853 2346
rect 3938 2343 3941 2393
rect 3946 2326 3949 2416
rect 3954 2333 3957 2416
rect 4042 2413 4053 2416
rect 4058 2413 4061 2426
rect 4098 2413 4101 2616
rect 4130 2613 4133 2703
rect 4146 2613 4149 2706
rect 4114 2523 4117 2556
rect 4146 2553 4149 2606
rect 3946 2323 3957 2326
rect 3742 2303 3749 2306
rect 3506 2213 3525 2216
rect 3562 2213 3565 2236
rect 3586 2203 3589 2286
rect 3602 2223 3605 2296
rect 3610 2233 3613 2266
rect 3506 2133 3509 2196
rect 3530 2156 3533 2176
rect 3526 2153 3533 2156
rect 3482 2123 3501 2126
rect 3474 2033 3485 2036
rect 3450 2023 3461 2026
rect 3450 1913 3453 1986
rect 3458 1913 3461 2023
rect 3466 2013 3469 2026
rect 3466 1973 3469 2006
rect 3474 1956 3477 2026
rect 3470 1953 3477 1956
rect 3442 1893 3453 1896
rect 3418 1753 3425 1756
rect 3394 1713 3397 1726
rect 3402 1723 3405 1746
rect 3402 1593 3405 1636
rect 3386 1473 3389 1526
rect 3362 1413 3381 1416
rect 3330 1293 3341 1296
rect 3250 1143 3269 1146
rect 3250 1136 3253 1143
rect 3242 1133 3253 1136
rect 3202 1113 3205 1126
rect 3194 1063 3197 1106
rect 3210 1103 3213 1116
rect 3218 1076 3221 1126
rect 3226 1086 3229 1126
rect 3234 1096 3237 1126
rect 3250 1113 3253 1126
rect 3258 1096 3261 1136
rect 3234 1093 3245 1096
rect 3226 1083 3237 1086
rect 3218 1073 3229 1076
rect 3194 1003 3197 1016
rect 3226 1013 3229 1073
rect 3234 1013 3237 1083
rect 3242 1013 3245 1093
rect 3254 1093 3261 1096
rect 3254 1026 3257 1093
rect 3254 1023 3261 1026
rect 3218 933 3229 936
rect 3234 933 3237 1006
rect 3194 923 3205 926
rect 3210 866 3213 926
rect 3242 923 3245 1006
rect 3258 1003 3261 1023
rect 3250 896 3253 936
rect 3242 893 3253 896
rect 3202 863 3213 866
rect 3178 833 3189 836
rect 3178 813 3181 826
rect 3138 686 3141 806
rect 3154 803 3165 806
rect 3170 763 3173 806
rect 3162 733 3165 746
rect 3186 733 3189 833
rect 3194 783 3197 826
rect 3202 813 3205 863
rect 3218 856 3221 866
rect 3210 853 3221 856
rect 3194 723 3197 766
rect 3202 733 3205 806
rect 3210 803 3213 853
rect 3122 683 3141 686
rect 3074 523 3109 526
rect 3122 523 3125 683
rect 3130 533 3133 546
rect 3042 413 3045 436
rect 3074 426 3077 516
rect 3050 403 3053 416
rect 3058 413 3061 426
rect 3074 423 3085 426
rect 3130 423 3133 526
rect 3082 406 3085 423
rect 3066 403 3085 406
rect 3010 293 3021 296
rect 2938 123 2941 166
rect 2962 123 2965 136
rect 2994 123 2997 206
rect 3002 163 3005 216
rect 3018 213 3021 293
rect 3010 183 3013 206
rect 3018 193 3021 206
rect 3026 173 3029 216
rect 3042 163 3045 336
rect 3050 323 3053 376
rect 3066 323 3069 403
rect 3122 383 3125 416
rect 3146 393 3149 606
rect 3170 603 3173 636
rect 3210 633 3213 786
rect 3218 763 3221 816
rect 3226 803 3229 826
rect 3234 813 3237 836
rect 3234 776 3237 796
rect 3230 773 3237 776
rect 3230 716 3233 773
rect 3242 753 3245 893
rect 3258 886 3261 936
rect 3250 883 3261 886
rect 3250 813 3253 883
rect 3266 833 3269 1143
rect 3274 1116 3277 1196
rect 3282 1193 3293 1196
rect 3282 1123 3285 1193
rect 3274 1113 3285 1116
rect 3274 1013 3277 1096
rect 3282 1056 3285 1113
rect 3290 1076 3293 1136
rect 3298 1133 3301 1256
rect 3306 1086 3309 1216
rect 3330 1196 3333 1293
rect 3330 1193 3341 1196
rect 3338 1173 3341 1193
rect 3314 1123 3317 1136
rect 3306 1083 3313 1086
rect 3290 1073 3301 1076
rect 3282 1053 3289 1056
rect 3274 933 3277 1006
rect 3286 956 3289 1053
rect 3282 953 3289 956
rect 3274 853 3277 926
rect 3282 893 3285 953
rect 3290 833 3293 936
rect 3298 926 3301 1073
rect 3310 1036 3313 1083
rect 3306 1033 3313 1036
rect 3306 1013 3309 1033
rect 3322 1013 3325 1136
rect 3330 1123 3333 1146
rect 3346 1133 3349 1376
rect 3354 1333 3357 1406
rect 3370 1393 3373 1406
rect 3378 1323 3381 1406
rect 3354 1213 3357 1226
rect 3362 1186 3365 1216
rect 3370 1213 3373 1236
rect 3354 1183 3365 1186
rect 3330 1013 3333 1036
rect 3314 993 3317 1006
rect 3322 1003 3333 1006
rect 3338 1003 3341 1116
rect 3346 1103 3349 1126
rect 3354 1086 3357 1183
rect 3362 1133 3365 1176
rect 3362 1103 3365 1126
rect 3370 1123 3373 1206
rect 3346 1083 3357 1086
rect 3346 1013 3349 1083
rect 3378 1056 3381 1316
rect 3386 1176 3389 1446
rect 3394 1286 3397 1536
rect 3402 1373 3405 1516
rect 3410 1346 3413 1736
rect 3422 1546 3425 1753
rect 3434 1733 3437 1746
rect 3442 1733 3445 1816
rect 3434 1653 3437 1716
rect 3450 1713 3453 1893
rect 3470 1886 3473 1953
rect 3482 1913 3485 2033
rect 3490 1956 3493 2116
rect 3498 2036 3501 2123
rect 3514 2113 3517 2126
rect 3526 2086 3529 2153
rect 3526 2083 3533 2086
rect 3498 2033 3525 2036
rect 3498 1983 3501 2006
rect 3506 2003 3509 2016
rect 3514 2013 3517 2026
rect 3522 2003 3525 2033
rect 3530 2013 3533 2083
rect 3538 2013 3541 2126
rect 3490 1953 3501 1956
rect 3498 1926 3501 1953
rect 3506 1936 3509 1976
rect 3538 1943 3541 2006
rect 3546 1963 3549 2126
rect 3562 2113 3565 2136
rect 3554 2013 3565 2016
rect 3554 1993 3557 2006
rect 3570 1953 3573 2166
rect 3602 2103 3605 2156
rect 3610 2123 3613 2136
rect 3618 2123 3621 2206
rect 3586 1946 3589 2006
rect 3610 1993 3613 2016
rect 3506 1933 3517 1936
rect 3482 1893 3485 1906
rect 3470 1883 3477 1886
rect 3466 1773 3469 1856
rect 3474 1753 3477 1883
rect 3482 1743 3485 1816
rect 3490 1813 3493 1926
rect 3498 1923 3509 1926
rect 3498 1873 3501 1916
rect 3506 1856 3509 1923
rect 3498 1853 3509 1856
rect 3498 1813 3501 1853
rect 3514 1826 3517 1933
rect 3522 1833 3525 1936
rect 3530 1926 3533 1936
rect 3530 1923 3549 1926
rect 3506 1823 3517 1826
rect 3506 1813 3509 1823
rect 3538 1816 3541 1916
rect 3554 1913 3557 1936
rect 3546 1823 3549 1896
rect 3554 1833 3557 1866
rect 3562 1816 3565 1936
rect 3570 1853 3573 1946
rect 3586 1943 3597 1946
rect 3586 1916 3589 1936
rect 3582 1913 3589 1916
rect 3582 1836 3585 1913
rect 3582 1833 3589 1836
rect 3514 1813 3533 1816
rect 3538 1813 3549 1816
rect 3490 1793 3493 1806
rect 3498 1743 3501 1766
rect 3442 1703 3453 1706
rect 3458 1686 3461 1726
rect 3482 1723 3485 1736
rect 3506 1723 3509 1806
rect 3514 1783 3517 1813
rect 3522 1793 3525 1806
rect 3514 1716 3517 1756
rect 3450 1683 3461 1686
rect 3434 1553 3437 1616
rect 3450 1606 3453 1683
rect 3466 1633 3469 1716
rect 3510 1713 3517 1716
rect 3482 1616 3485 1706
rect 3446 1603 3453 1606
rect 3418 1543 3425 1546
rect 3418 1413 3421 1543
rect 3410 1343 3421 1346
rect 3410 1323 3413 1336
rect 3394 1283 3405 1286
rect 3402 1213 3405 1283
rect 3418 1253 3421 1343
rect 3434 1336 3437 1526
rect 3446 1466 3449 1603
rect 3458 1476 3461 1616
rect 3478 1613 3485 1616
rect 3498 1613 3501 1676
rect 3510 1636 3513 1713
rect 3522 1703 3525 1776
rect 3530 1713 3533 1806
rect 3538 1763 3541 1806
rect 3546 1676 3549 1813
rect 3542 1673 3549 1676
rect 3554 1813 3565 1816
rect 3570 1813 3573 1826
rect 3586 1816 3589 1833
rect 3578 1813 3589 1816
rect 3506 1633 3513 1636
rect 3466 1533 3469 1566
rect 3478 1526 3481 1613
rect 3506 1606 3509 1633
rect 3522 1623 3525 1636
rect 3490 1533 3493 1606
rect 3498 1603 3509 1606
rect 3466 1503 3469 1526
rect 3478 1523 3485 1526
rect 3458 1473 3465 1476
rect 3446 1463 3453 1466
rect 3450 1443 3453 1463
rect 3462 1406 3465 1473
rect 3458 1403 3465 1406
rect 3458 1383 3461 1403
rect 3426 1333 3437 1336
rect 3458 1333 3461 1346
rect 3394 1193 3397 1206
rect 3410 1186 3413 1206
rect 3402 1183 3413 1186
rect 3386 1173 3393 1176
rect 3426 1173 3429 1333
rect 3474 1303 3477 1486
rect 3482 1443 3485 1523
rect 3482 1393 3485 1416
rect 3482 1256 3485 1386
rect 3490 1313 3493 1336
rect 3498 1323 3501 1603
rect 3498 1276 3501 1296
rect 3466 1253 3485 1256
rect 3494 1273 3501 1276
rect 3450 1193 3453 1216
rect 3466 1176 3469 1253
rect 3494 1186 3497 1273
rect 3494 1183 3501 1186
rect 3466 1173 3477 1176
rect 3370 1053 3381 1056
rect 3306 933 3309 986
rect 3322 943 3325 966
rect 3298 923 3317 926
rect 3306 846 3309 896
rect 3322 856 3325 936
rect 3330 863 3333 1003
rect 3338 923 3341 976
rect 3346 933 3349 1006
rect 3354 1003 3357 1046
rect 3362 996 3365 1016
rect 3354 993 3365 996
rect 3354 926 3357 993
rect 3362 933 3365 946
rect 3370 933 3373 1053
rect 3390 1046 3393 1173
rect 3410 1113 3413 1126
rect 3386 1043 3393 1046
rect 3354 923 3373 926
rect 3378 886 3381 1016
rect 3386 1013 3389 1043
rect 3394 1013 3397 1026
rect 3410 1006 3413 1016
rect 3386 933 3389 1006
rect 3394 1003 3413 1006
rect 3394 933 3397 1003
rect 3402 933 3405 966
rect 3378 883 3389 886
rect 3322 853 3349 856
rect 3302 843 3309 846
rect 3282 813 3285 826
rect 3302 796 3305 843
rect 3302 793 3309 796
rect 3306 776 3309 793
rect 3330 783 3333 846
rect 3346 813 3349 853
rect 3378 813 3381 836
rect 3306 773 3325 776
rect 3242 723 3245 736
rect 3230 713 3237 716
rect 3210 613 3213 626
rect 3162 513 3165 526
rect 3170 383 3173 526
rect 3186 516 3189 536
rect 3194 533 3197 546
rect 3202 523 3205 536
rect 3182 513 3189 516
rect 3182 446 3185 513
rect 3182 443 3189 446
rect 3186 423 3189 443
rect 3194 433 3197 506
rect 3218 436 3221 596
rect 3234 593 3237 713
rect 3242 496 3245 636
rect 3250 533 3253 726
rect 3214 433 3221 436
rect 3234 493 3245 496
rect 3202 413 3205 426
rect 3074 333 3077 346
rect 3050 213 3061 216
rect 3050 193 3053 206
rect 3066 203 3069 306
rect 3082 263 3085 326
rect 3154 323 3157 356
rect 3202 286 3205 396
rect 3214 376 3217 433
rect 3214 373 3221 376
rect 3218 353 3221 373
rect 3226 343 3229 426
rect 3234 413 3237 493
rect 3242 403 3245 416
rect 3250 413 3253 426
rect 3258 373 3261 656
rect 3274 616 3277 766
rect 3266 603 3269 616
rect 3274 613 3285 616
rect 3274 593 3277 606
rect 3290 603 3293 626
rect 3298 603 3301 736
rect 3306 723 3309 736
rect 3314 706 3317 756
rect 3310 703 3317 706
rect 3310 626 3313 703
rect 3322 633 3325 773
rect 3310 623 3317 626
rect 3314 603 3317 623
rect 3266 513 3269 526
rect 3314 523 3317 546
rect 3266 413 3269 456
rect 3274 406 3277 416
rect 3266 403 3277 406
rect 3266 393 3269 403
rect 3226 323 3229 336
rect 3250 296 3253 346
rect 3258 323 3261 356
rect 3274 323 3277 346
rect 3306 323 3309 406
rect 3314 403 3317 446
rect 3322 396 3325 616
rect 3330 613 3333 736
rect 3338 676 3341 746
rect 3346 713 3349 786
rect 3362 723 3365 736
rect 3378 733 3381 746
rect 3386 726 3389 883
rect 3394 763 3397 926
rect 3402 776 3405 926
rect 3410 923 3413 986
rect 3418 943 3421 1006
rect 3418 883 3421 936
rect 3426 926 3429 996
rect 3434 983 3437 1146
rect 3474 1143 3477 1173
rect 3458 1093 3461 1136
rect 3474 1023 3477 1136
rect 3482 1123 3485 1136
rect 3498 1133 3501 1183
rect 3490 1123 3501 1126
rect 3506 1056 3509 1596
rect 3514 1453 3517 1616
rect 3514 1293 3517 1446
rect 3522 1316 3525 1556
rect 3530 1413 3533 1606
rect 3542 1576 3545 1673
rect 3542 1573 3549 1576
rect 3546 1553 3549 1573
rect 3530 1366 3533 1386
rect 3538 1373 3541 1546
rect 3546 1466 3549 1526
rect 3554 1483 3557 1813
rect 3562 1783 3565 1806
rect 3562 1723 3565 1766
rect 3578 1733 3581 1746
rect 3594 1743 3597 1943
rect 3610 1846 3613 1916
rect 3618 1856 3621 2116
rect 3626 1913 3629 2226
rect 3634 2223 3637 2236
rect 3642 2203 3645 2236
rect 3650 2183 3653 2216
rect 3658 2176 3661 2226
rect 3742 2216 3745 2303
rect 3674 2193 3677 2206
rect 3650 2173 3661 2176
rect 3634 1933 3637 2126
rect 3650 2113 3653 2173
rect 3682 2133 3685 2156
rect 3658 2083 3661 2106
rect 3666 2103 3669 2126
rect 3674 2066 3677 2116
rect 3682 2083 3685 2126
rect 3666 2063 3677 2066
rect 3666 1996 3669 2063
rect 3666 1993 3677 1996
rect 3674 1973 3677 1993
rect 3690 1946 3693 2186
rect 3698 2133 3701 2216
rect 3738 2213 3745 2216
rect 3714 2153 3717 2186
rect 3706 2113 3709 2126
rect 3714 2123 3717 2146
rect 3722 2083 3725 2126
rect 3738 2113 3741 2213
rect 3754 2146 3757 2306
rect 3810 2246 3813 2313
rect 3994 2293 3997 2406
rect 4042 2393 4045 2413
rect 4042 2283 4045 2346
rect 4058 2313 4061 2326
rect 4090 2323 4093 2376
rect 4138 2333 4141 2536
rect 4154 2296 4157 2753
rect 4146 2293 4157 2296
rect 3810 2243 3821 2246
rect 3770 2186 3773 2216
rect 3770 2183 3781 2186
rect 3746 2143 3757 2146
rect 3746 2103 3749 2143
rect 3770 2133 3773 2176
rect 3754 2123 3765 2126
rect 3698 2013 3701 2026
rect 3690 1943 3697 1946
rect 3634 1903 3637 1926
rect 3642 1903 3645 1926
rect 3618 1853 3637 1856
rect 3650 1853 3653 1916
rect 3666 1906 3669 1936
rect 3662 1903 3669 1906
rect 3610 1843 3621 1846
rect 3610 1813 3613 1836
rect 3618 1793 3621 1843
rect 3562 1676 3565 1716
rect 3562 1673 3573 1676
rect 3570 1586 3573 1673
rect 3602 1636 3605 1726
rect 3562 1583 3573 1586
rect 3594 1633 3605 1636
rect 3546 1463 3553 1466
rect 3550 1366 3553 1463
rect 3562 1403 3565 1583
rect 3586 1523 3589 1566
rect 3594 1533 3597 1633
rect 3610 1586 3613 1786
rect 3634 1776 3637 1853
rect 3662 1846 3665 1903
rect 3694 1896 3697 1943
rect 3690 1893 3697 1896
rect 3706 1893 3709 2046
rect 3722 1986 3725 2016
rect 3738 1993 3741 2006
rect 3746 1996 3749 2066
rect 3754 2023 3757 2116
rect 3762 2063 3765 2123
rect 3770 2086 3773 2126
rect 3778 2113 3781 2183
rect 3786 2153 3789 2206
rect 3818 2196 3821 2243
rect 3834 2203 3837 2216
rect 3802 2193 3821 2196
rect 3786 2123 3789 2136
rect 3770 2083 3781 2086
rect 3762 2033 3765 2056
rect 3770 2013 3773 2026
rect 3746 1993 3757 1996
rect 3722 1983 3741 1986
rect 3714 1923 3717 1946
rect 3658 1843 3665 1846
rect 3658 1786 3661 1843
rect 3674 1823 3677 1876
rect 3690 1873 3693 1893
rect 3682 1833 3685 1846
rect 3690 1813 3693 1836
rect 3658 1783 3677 1786
rect 3634 1773 3649 1776
rect 3618 1633 3621 1696
rect 3646 1636 3649 1773
rect 3646 1633 3653 1636
rect 3626 1613 3637 1616
rect 3610 1583 3621 1586
rect 3602 1523 3605 1536
rect 3610 1533 3613 1576
rect 3570 1413 3581 1416
rect 3586 1413 3589 1426
rect 3570 1403 3581 1406
rect 3570 1393 3573 1403
rect 3594 1396 3597 1406
rect 3578 1393 3597 1396
rect 3530 1363 3541 1366
rect 3530 1323 3533 1336
rect 3538 1333 3541 1363
rect 3546 1363 3553 1366
rect 3522 1313 3533 1316
rect 3514 1153 3517 1256
rect 3514 1103 3517 1126
rect 3522 1113 3525 1306
rect 3482 1053 3509 1056
rect 3458 1003 3461 1016
rect 3434 933 3437 976
rect 3426 923 3445 926
rect 3466 893 3469 1016
rect 3426 793 3429 806
rect 3402 773 3421 776
rect 3410 733 3413 746
rect 3378 723 3389 726
rect 3394 723 3405 726
rect 3354 693 3357 706
rect 3338 673 3349 676
rect 3330 523 3333 606
rect 3330 403 3333 516
rect 3338 413 3341 546
rect 3346 503 3349 673
rect 3354 496 3357 526
rect 3346 493 3357 496
rect 3314 393 3325 396
rect 3314 333 3317 393
rect 3322 333 3325 356
rect 3330 323 3333 396
rect 3346 353 3349 493
rect 3362 413 3365 626
rect 3370 603 3373 616
rect 3378 613 3381 723
rect 3386 703 3389 716
rect 3418 706 3421 773
rect 3426 773 3445 776
rect 3450 773 3453 816
rect 3474 813 3477 886
rect 3482 783 3485 1053
rect 3522 1013 3525 1026
rect 3506 993 3509 1006
rect 3530 1003 3533 1313
rect 3538 1293 3541 1326
rect 3546 1303 3549 1363
rect 3554 1333 3557 1346
rect 3562 1313 3565 1386
rect 3570 1333 3573 1376
rect 3570 1296 3573 1326
rect 3562 1293 3573 1296
rect 3562 1246 3565 1293
rect 3562 1243 3573 1246
rect 3538 1213 3541 1226
rect 3546 1213 3549 1236
rect 3570 1213 3573 1243
rect 3546 1163 3549 1206
rect 3562 1163 3565 1206
rect 3578 1183 3581 1393
rect 3602 1383 3605 1416
rect 3594 1333 3597 1376
rect 3618 1276 3621 1583
rect 3642 1563 3645 1616
rect 3626 1523 3629 1536
rect 3642 1473 3645 1526
rect 3650 1463 3653 1633
rect 3658 1533 3661 1726
rect 3674 1723 3677 1783
rect 3698 1746 3701 1826
rect 3706 1813 3709 1826
rect 3714 1823 3717 1836
rect 3722 1803 3725 1816
rect 3730 1763 3733 1826
rect 3738 1813 3741 1983
rect 3754 1896 3757 1993
rect 3778 1986 3781 2083
rect 3802 2043 3805 2193
rect 3810 2133 3813 2176
rect 3818 2133 3821 2146
rect 3810 2106 3813 2126
rect 3810 2103 3817 2106
rect 3826 2103 3829 2126
rect 3834 2113 3837 2136
rect 3850 2133 3861 2136
rect 3866 2133 3869 2206
rect 3882 2176 3885 2216
rect 3898 2183 3901 2206
rect 3874 2173 3885 2176
rect 3814 2036 3817 2103
rect 3810 2033 3817 2036
rect 3786 1993 3789 2016
rect 3778 1983 3789 1986
rect 3778 1913 3781 1926
rect 3750 1893 3757 1896
rect 3750 1806 3753 1893
rect 3746 1803 3753 1806
rect 3746 1776 3749 1803
rect 3742 1773 3749 1776
rect 3698 1743 3709 1746
rect 3706 1696 3709 1743
rect 3722 1713 3725 1726
rect 3698 1693 3709 1696
rect 3666 1593 3669 1626
rect 3626 1413 3629 1436
rect 3626 1323 3629 1346
rect 3634 1333 3637 1406
rect 3610 1273 3621 1276
rect 3586 1213 3589 1226
rect 3610 1186 3613 1273
rect 3610 1183 3621 1186
rect 3538 1123 3541 1136
rect 3554 1133 3557 1146
rect 3538 973 3541 1116
rect 3546 1013 3549 1036
rect 3546 956 3549 996
rect 3542 953 3549 956
rect 3490 913 3493 936
rect 3426 733 3429 773
rect 3442 766 3445 773
rect 3410 703 3421 706
rect 3410 646 3413 703
rect 3410 643 3421 646
rect 3386 606 3389 636
rect 3418 623 3421 643
rect 3402 613 3421 616
rect 3426 613 3429 726
rect 3378 603 3389 606
rect 3378 593 3381 603
rect 3378 533 3381 566
rect 3394 546 3397 606
rect 3410 593 3413 606
rect 3418 603 3421 613
rect 3434 566 3437 766
rect 3442 763 3453 766
rect 3442 633 3445 763
rect 3474 723 3477 746
rect 3450 613 3453 706
rect 3442 583 3445 606
rect 3458 603 3461 626
rect 3466 613 3469 656
rect 3466 566 3469 606
rect 3474 603 3477 636
rect 3482 603 3485 616
rect 3490 613 3493 896
rect 3506 876 3509 936
rect 3530 923 3533 936
rect 3498 873 3509 876
rect 3498 793 3501 873
rect 3514 763 3517 876
rect 3530 813 3533 916
rect 3542 846 3545 953
rect 3554 873 3557 1116
rect 3578 1106 3581 1156
rect 3586 1123 3589 1166
rect 3578 1103 3585 1106
rect 3562 983 3565 1006
rect 3570 1003 3573 1056
rect 3582 1026 3585 1103
rect 3578 1023 3585 1026
rect 3578 996 3581 1023
rect 3594 1013 3597 1126
rect 3570 993 3581 996
rect 3586 993 3589 1006
rect 3542 843 3549 846
rect 3522 733 3525 796
rect 3546 656 3549 843
rect 3570 696 3573 993
rect 3578 906 3581 976
rect 3586 923 3589 986
rect 3594 913 3597 1006
rect 3578 903 3585 906
rect 3538 653 3549 656
rect 3562 693 3573 696
rect 3498 613 3501 626
rect 3514 613 3517 626
rect 3410 563 3437 566
rect 3458 563 3469 566
rect 3410 546 3413 563
rect 3394 543 3405 546
rect 3410 543 3421 546
rect 3378 473 3381 526
rect 3402 523 3405 543
rect 3386 413 3397 416
rect 3338 333 3341 346
rect 3346 323 3349 336
rect 3198 283 3205 286
rect 3058 123 3061 166
rect 3066 123 3069 176
rect 3074 133 3077 216
rect 3114 193 3117 216
rect 3130 183 3133 216
rect 3178 213 3181 226
rect 3098 123 3101 136
rect 3146 123 3149 196
rect 3162 183 3165 206
rect 3186 173 3189 276
rect 3198 226 3201 283
rect 3194 223 3201 226
rect 3194 183 3197 223
rect 3202 193 3205 206
rect 3210 196 3213 216
rect 3218 203 3221 216
rect 3226 213 3229 296
rect 3242 293 3253 296
rect 3242 213 3245 293
rect 3258 213 3261 266
rect 3226 196 3229 206
rect 3266 203 3269 226
rect 3274 213 3277 236
rect 3282 206 3285 276
rect 3354 273 3357 406
rect 3378 333 3381 406
rect 3386 393 3389 406
rect 3402 403 3405 506
rect 3418 446 3421 543
rect 3458 506 3461 563
rect 3474 523 3477 586
rect 3490 543 3493 606
rect 3506 553 3509 606
rect 3458 503 3469 506
rect 3466 486 3469 503
rect 3466 483 3473 486
rect 3410 443 3421 446
rect 3410 336 3413 443
rect 3426 383 3429 406
rect 3450 393 3453 416
rect 3458 343 3461 466
rect 3470 336 3473 483
rect 3490 393 3493 536
rect 3514 523 3517 546
rect 3522 533 3525 606
rect 3538 563 3541 653
rect 3562 646 3565 693
rect 3582 686 3585 903
rect 3602 883 3605 1166
rect 3610 1003 3613 1046
rect 3610 903 3613 956
rect 3594 793 3597 816
rect 3618 776 3621 1183
rect 3626 1053 3629 1296
rect 3642 1213 3645 1416
rect 3658 1403 3661 1426
rect 3666 1413 3669 1436
rect 3674 1346 3677 1656
rect 3698 1633 3701 1693
rect 3698 1613 3717 1616
rect 3690 1543 3693 1606
rect 3666 1343 3677 1346
rect 3666 1276 3669 1343
rect 3674 1323 3677 1336
rect 3658 1273 3669 1276
rect 3634 1123 3637 1206
rect 3642 1173 3653 1176
rect 3650 1133 3653 1173
rect 3658 1166 3661 1273
rect 3682 1223 3685 1436
rect 3690 1216 3693 1536
rect 3698 1523 3701 1606
rect 3706 1573 3709 1606
rect 3714 1533 3717 1613
rect 3722 1603 3725 1636
rect 3714 1436 3717 1526
rect 3706 1433 3717 1436
rect 3698 1413 3701 1426
rect 3698 1223 3701 1406
rect 3706 1306 3709 1433
rect 3714 1403 3717 1426
rect 3714 1323 3717 1336
rect 3722 1323 3725 1596
rect 3730 1506 3733 1646
rect 3742 1626 3745 1773
rect 3742 1623 3749 1626
rect 3738 1523 3741 1606
rect 3730 1503 3737 1506
rect 3734 1426 3737 1503
rect 3746 1433 3749 1623
rect 3730 1423 3737 1426
rect 3730 1343 3733 1423
rect 3754 1416 3757 1766
rect 3762 1643 3765 1876
rect 3786 1813 3789 1983
rect 3794 1813 3797 2026
rect 3802 2003 3805 2016
rect 3810 2013 3813 2033
rect 3826 2013 3829 2026
rect 3802 1903 3805 1926
rect 3818 1886 3821 1996
rect 3834 1993 3837 2036
rect 3842 2013 3845 2126
rect 3850 2016 3853 2126
rect 3874 2113 3877 2173
rect 3898 2136 3901 2156
rect 3850 2013 3861 2016
rect 3842 1983 3845 2006
rect 3850 1993 3853 2006
rect 3826 1933 3829 1956
rect 3834 1906 3837 1966
rect 3850 1933 3853 1946
rect 3842 1913 3845 1926
rect 3810 1883 3821 1886
rect 3826 1903 3837 1906
rect 3770 1783 3773 1806
rect 3778 1733 3781 1796
rect 3794 1726 3797 1806
rect 3802 1803 3805 1816
rect 3770 1603 3773 1726
rect 3778 1723 3797 1726
rect 3802 1713 3805 1736
rect 3810 1646 3813 1883
rect 3818 1783 3821 1816
rect 3826 1773 3829 1903
rect 3834 1756 3837 1856
rect 3842 1803 3845 1816
rect 3830 1753 3837 1756
rect 3802 1643 3813 1646
rect 3770 1523 3773 1546
rect 3778 1506 3781 1556
rect 3774 1503 3781 1506
rect 3746 1413 3757 1416
rect 3738 1393 3741 1406
rect 3706 1303 3717 1306
rect 3714 1226 3717 1303
rect 3706 1223 3717 1226
rect 3682 1213 3701 1216
rect 3658 1163 3669 1166
rect 3666 1153 3669 1163
rect 3674 1123 3677 1206
rect 3634 1003 3637 1096
rect 3658 993 3661 1016
rect 3626 926 3629 986
rect 3666 983 3669 1076
rect 3674 976 3677 1056
rect 3682 983 3685 1206
rect 3690 1183 3693 1206
rect 3690 1073 3693 1156
rect 3698 1076 3701 1206
rect 3706 1163 3709 1223
rect 3730 1213 3733 1336
rect 3738 1293 3741 1376
rect 3754 1366 3757 1406
rect 3762 1373 3765 1476
rect 3774 1436 3777 1503
rect 3774 1433 3781 1436
rect 3770 1393 3773 1416
rect 3754 1363 3765 1366
rect 3746 1303 3749 1356
rect 3754 1283 3757 1346
rect 3762 1236 3765 1363
rect 3778 1356 3781 1433
rect 3786 1413 3789 1576
rect 3794 1523 3797 1566
rect 3802 1553 3805 1643
rect 3810 1613 3813 1636
rect 3818 1563 3821 1736
rect 3830 1666 3833 1753
rect 3842 1743 3845 1796
rect 3830 1663 3837 1666
rect 3818 1533 3821 1546
rect 3834 1536 3837 1663
rect 3842 1573 3845 1736
rect 3850 1653 3853 1856
rect 3858 1723 3861 2013
rect 3866 1993 3869 2006
rect 3874 1983 3877 2016
rect 3882 1963 3885 2136
rect 3898 2133 3905 2136
rect 3914 2133 3925 2136
rect 3930 2133 3933 2216
rect 3890 2093 3893 2126
rect 3902 2086 3905 2133
rect 3914 2113 3917 2126
rect 3898 2083 3905 2086
rect 3898 2003 3901 2083
rect 3922 2026 3925 2133
rect 3938 2126 3941 2146
rect 3946 2133 3949 2166
rect 3978 2133 3981 2216
rect 3938 2123 3957 2126
rect 3922 2023 3941 2026
rect 3922 1993 3925 2016
rect 3938 1966 3941 2023
rect 3962 2016 3965 2036
rect 3962 2013 3969 2016
rect 3874 1933 3877 1946
rect 3906 1943 3909 1966
rect 3930 1963 3941 1966
rect 3890 1923 3893 1936
rect 3866 1896 3869 1916
rect 3914 1913 3917 1926
rect 3866 1893 3877 1896
rect 3874 1836 3877 1893
rect 3930 1886 3933 1963
rect 3930 1883 3949 1886
rect 3866 1833 3877 1836
rect 3866 1803 3869 1833
rect 3890 1816 3893 1826
rect 3874 1813 3893 1816
rect 3898 1816 3901 1846
rect 3898 1813 3909 1816
rect 3914 1813 3917 1836
rect 3882 1776 3885 1806
rect 3890 1803 3893 1813
rect 3882 1773 3893 1776
rect 3874 1706 3877 1736
rect 3890 1733 3893 1773
rect 3866 1703 3877 1706
rect 3882 1706 3885 1726
rect 3882 1703 3889 1706
rect 3866 1656 3869 1703
rect 3866 1653 3877 1656
rect 3874 1633 3877 1653
rect 3886 1636 3889 1703
rect 3882 1633 3889 1636
rect 3882 1613 3885 1633
rect 3834 1533 3845 1536
rect 3794 1406 3797 1516
rect 3818 1433 3821 1526
rect 3834 1513 3837 1526
rect 3802 1413 3821 1416
rect 3786 1373 3789 1406
rect 3794 1403 3805 1406
rect 3810 1403 3821 1406
rect 3826 1403 3829 1506
rect 3842 1493 3845 1533
rect 3810 1356 3813 1403
rect 3770 1353 3781 1356
rect 3802 1353 3813 1356
rect 3770 1303 3773 1353
rect 3778 1333 3781 1346
rect 3802 1333 3805 1353
rect 3818 1333 3821 1386
rect 3834 1353 3837 1416
rect 3842 1413 3845 1426
rect 3842 1356 3845 1406
rect 3850 1383 3853 1546
rect 3858 1403 3861 1586
rect 3874 1503 3877 1526
rect 3866 1403 3869 1436
rect 3858 1356 3861 1376
rect 3874 1373 3877 1446
rect 3842 1353 3853 1356
rect 3858 1353 3865 1356
rect 3778 1323 3789 1326
rect 3842 1323 3845 1346
rect 3786 1313 3789 1323
rect 3850 1306 3853 1353
rect 3746 1213 3749 1236
rect 3754 1233 3765 1236
rect 3714 1126 3717 1206
rect 3722 1183 3725 1206
rect 3738 1193 3741 1206
rect 3746 1133 3749 1176
rect 3754 1163 3757 1233
rect 3770 1143 3773 1206
rect 3794 1193 3797 1216
rect 3802 1176 3805 1266
rect 3778 1173 3805 1176
rect 3778 1136 3781 1173
rect 3770 1133 3781 1136
rect 3714 1123 3733 1126
rect 3698 1073 3705 1076
rect 3674 973 3693 976
rect 3634 933 3653 936
rect 3658 933 3661 946
rect 3666 933 3669 956
rect 3626 923 3645 926
rect 3626 913 3637 916
rect 3626 893 3629 906
rect 3634 866 3637 886
rect 3630 863 3637 866
rect 3630 786 3633 863
rect 3630 783 3637 786
rect 3614 773 3621 776
rect 3594 723 3597 746
rect 3614 706 3617 773
rect 3626 713 3629 766
rect 3614 703 3621 706
rect 3578 683 3585 686
rect 3562 643 3569 646
rect 3566 596 3569 643
rect 3562 593 3569 596
rect 3538 536 3541 556
rect 3534 533 3541 536
rect 3410 333 3421 336
rect 3402 276 3405 326
rect 3418 286 3421 333
rect 3466 333 3473 336
rect 3498 333 3509 336
rect 3394 273 3405 276
rect 3410 283 3421 286
rect 3442 323 3461 326
rect 3298 213 3301 226
rect 3274 203 3285 206
rect 3210 193 3229 196
rect 3210 186 3213 193
rect 3202 183 3213 186
rect 3202 123 3205 183
rect 3218 133 3221 186
rect 3274 173 3277 203
rect 3266 123 3269 136
rect 3290 133 3293 206
rect 3306 203 3309 256
rect 3314 123 3317 226
rect 3322 213 3325 236
rect 3394 226 3397 273
rect 3410 263 3413 283
rect 3394 223 3405 226
rect 3322 173 3325 206
rect 3338 186 3341 206
rect 3330 133 3333 186
rect 3338 183 3349 186
rect 3338 163 3341 183
rect 3354 123 3357 206
rect 3362 203 3365 216
rect 3370 213 3381 216
rect 3370 173 3373 206
rect 3378 183 3381 206
rect 3402 203 3405 223
rect 3410 213 3429 216
rect 3418 193 3421 206
rect 3426 123 3429 206
rect 3442 203 3445 323
rect 3466 313 3469 333
rect 3482 323 3493 326
rect 3458 213 3461 296
rect 3474 243 3477 306
rect 3482 213 3485 316
rect 3490 233 3493 323
rect 3498 213 3501 326
rect 3482 203 3493 206
rect 3458 133 3461 156
rect 3498 143 3501 206
rect 3506 193 3509 333
rect 3514 313 3517 516
rect 3534 486 3537 533
rect 3562 513 3565 593
rect 3570 523 3573 536
rect 3578 513 3581 683
rect 3586 593 3589 616
rect 3594 516 3597 566
rect 3590 513 3597 516
rect 3610 513 3613 526
rect 3534 483 3541 486
rect 3522 413 3533 416
rect 3538 333 3541 483
rect 3554 393 3557 416
rect 3578 396 3581 416
rect 3570 393 3581 396
rect 3590 396 3593 513
rect 3590 393 3597 396
rect 3562 336 3565 376
rect 3554 333 3565 336
rect 3570 333 3573 393
rect 3594 373 3597 393
rect 3602 363 3605 506
rect 3586 336 3589 356
rect 3578 333 3589 336
rect 3610 333 3613 376
rect 3618 333 3621 703
rect 3634 696 3637 783
rect 3630 693 3637 696
rect 3630 556 3633 693
rect 3642 563 3645 923
rect 3650 813 3653 933
rect 3658 806 3661 926
rect 3674 913 3677 926
rect 3682 876 3685 946
rect 3690 883 3693 973
rect 3702 956 3705 1073
rect 3698 953 3705 956
rect 3698 923 3701 953
rect 3714 946 3717 1036
rect 3722 953 3725 1016
rect 3730 1013 3733 1026
rect 3738 1013 3749 1016
rect 3762 1013 3765 1036
rect 3730 1003 3749 1006
rect 3714 943 3725 946
rect 3674 873 3685 876
rect 3674 813 3677 873
rect 3650 803 3661 806
rect 3650 566 3653 803
rect 3666 773 3669 806
rect 3682 793 3685 806
rect 3658 733 3661 766
rect 3658 713 3661 726
rect 3658 613 3661 626
rect 3666 613 3669 756
rect 3674 733 3677 746
rect 3682 713 3685 786
rect 3690 753 3693 816
rect 3698 803 3701 906
rect 3706 783 3709 936
rect 3714 776 3717 926
rect 3682 613 3685 626
rect 3658 576 3661 606
rect 3674 593 3677 606
rect 3658 573 3677 576
rect 3650 563 3669 566
rect 3630 553 3637 556
rect 3626 513 3629 536
rect 3634 426 3637 553
rect 3642 456 3645 536
rect 3650 523 3653 536
rect 3642 453 3653 456
rect 3634 423 3645 426
rect 3538 323 3549 326
rect 3530 283 3533 306
rect 3546 303 3549 316
rect 3554 293 3557 326
rect 3514 203 3517 266
rect 3562 263 3565 333
rect 3626 326 3629 396
rect 3634 373 3637 416
rect 3642 383 3645 423
rect 3650 326 3653 453
rect 3658 423 3661 536
rect 3666 533 3669 563
rect 3674 523 3677 573
rect 3682 516 3685 606
rect 3690 583 3693 736
rect 3698 733 3701 776
rect 3706 773 3717 776
rect 3698 603 3701 726
rect 3706 613 3709 773
rect 3714 733 3717 766
rect 3714 636 3717 726
rect 3722 723 3725 943
rect 3730 833 3733 926
rect 3730 733 3733 746
rect 3738 723 3741 936
rect 3746 706 3749 1003
rect 3754 993 3757 1006
rect 3754 823 3757 986
rect 3770 933 3773 1133
rect 3786 1053 3789 1166
rect 3794 1123 3797 1146
rect 3810 1096 3813 1286
rect 3818 1166 3821 1306
rect 3846 1303 3853 1306
rect 3846 1246 3849 1303
rect 3862 1296 3865 1353
rect 3834 1243 3849 1246
rect 3858 1293 3865 1296
rect 3818 1163 3825 1166
rect 3822 1106 3825 1163
rect 3834 1133 3837 1243
rect 3834 1113 3837 1126
rect 3842 1123 3845 1236
rect 3858 1226 3861 1293
rect 3854 1223 3861 1226
rect 3854 1166 3857 1223
rect 3866 1213 3869 1226
rect 3882 1213 3885 1536
rect 3890 1443 3893 1616
rect 3890 1403 3893 1436
rect 3898 1413 3901 1806
rect 3906 1796 3909 1813
rect 3922 1803 3925 1846
rect 3938 1813 3941 1826
rect 3906 1793 3913 1796
rect 3910 1716 3913 1793
rect 3930 1756 3933 1806
rect 3930 1753 3941 1756
rect 3922 1733 3933 1736
rect 3910 1713 3917 1716
rect 3914 1636 3917 1713
rect 3906 1633 3917 1636
rect 3906 1613 3909 1633
rect 3914 1613 3925 1616
rect 3930 1603 3933 1726
rect 3938 1613 3941 1753
rect 3946 1743 3949 1883
rect 3946 1723 3949 1736
rect 3922 1533 3925 1576
rect 3938 1533 3941 1606
rect 3946 1563 3949 1716
rect 3946 1533 3949 1556
rect 3938 1486 3941 1526
rect 3954 1523 3957 1976
rect 3966 1946 3969 2013
rect 3962 1943 3969 1946
rect 3962 1706 3965 1943
rect 3970 1803 3973 1926
rect 3978 1756 3981 2126
rect 3986 2106 3989 2206
rect 3994 2123 3997 2216
rect 4002 2193 4005 2206
rect 4010 2173 4013 2216
rect 3986 2103 3993 2106
rect 3990 2036 3993 2103
rect 3986 2033 3993 2036
rect 4002 2033 4005 2136
rect 3986 1946 3989 2033
rect 3994 1983 3997 2016
rect 4002 2013 4005 2026
rect 4018 2016 4021 2206
rect 4034 2183 4037 2206
rect 4058 2193 4061 2216
rect 4026 2133 4029 2146
rect 4042 2133 4045 2166
rect 4010 2013 4021 2016
rect 4002 1963 4005 2006
rect 4010 1983 4013 2013
rect 4018 1993 4021 2006
rect 3986 1943 3997 1946
rect 3986 1853 3989 1936
rect 3994 1916 3997 1943
rect 4002 1933 4005 1946
rect 3994 1913 4001 1916
rect 3998 1836 4001 1913
rect 4010 1843 4013 1926
rect 4018 1906 4021 1936
rect 4026 1923 4029 2016
rect 4034 2013 4037 2126
rect 4066 2076 4069 2186
rect 4130 2173 4133 2216
rect 4146 2146 4149 2293
rect 4090 2123 4093 2146
rect 4146 2143 4157 2146
rect 4146 2106 4149 2126
rect 4050 2073 4069 2076
rect 4138 2103 4149 2106
rect 4034 1933 4037 2006
rect 4050 1976 4053 2073
rect 4138 2056 4141 2103
rect 4138 2053 4149 2056
rect 4074 1993 4077 2016
rect 4050 1973 4069 1976
rect 4042 1906 4045 1966
rect 4050 1933 4053 1956
rect 4066 1906 4069 1973
rect 4130 1953 4133 2016
rect 4138 2013 4141 2036
rect 4146 2003 4149 2053
rect 4090 1923 4093 1946
rect 4018 1903 4025 1906
rect 3994 1833 4001 1836
rect 3986 1793 3989 1806
rect 3970 1753 3981 1756
rect 3970 1723 3973 1753
rect 3978 1733 3981 1746
rect 3986 1713 3989 1726
rect 3962 1703 3973 1706
rect 3930 1483 3941 1486
rect 3914 1413 3917 1476
rect 3890 1253 3893 1396
rect 3898 1296 3901 1376
rect 3906 1303 3909 1406
rect 3930 1386 3933 1483
rect 3914 1383 3933 1386
rect 3914 1336 3917 1383
rect 3914 1333 3925 1336
rect 3914 1313 3917 1326
rect 3930 1323 3933 1336
rect 3938 1323 3941 1466
rect 3954 1413 3957 1496
rect 3946 1403 3957 1406
rect 3962 1373 3965 1636
rect 3970 1533 3973 1703
rect 3994 1633 3997 1833
rect 4022 1826 4025 1903
rect 4018 1823 4025 1826
rect 4034 1903 4045 1906
rect 4050 1903 4069 1906
rect 4002 1813 4013 1816
rect 4002 1803 4013 1806
rect 4018 1733 4021 1823
rect 4034 1763 4037 1903
rect 4034 1733 4037 1756
rect 4050 1753 4053 1903
rect 4074 1803 4077 1816
rect 4074 1776 4077 1796
rect 4070 1773 4077 1776
rect 4058 1723 4061 1746
rect 4070 1686 4073 1773
rect 4070 1683 4077 1686
rect 4074 1663 4077 1683
rect 4082 1676 4085 1766
rect 4114 1723 4117 1736
rect 4122 1723 4125 1816
rect 4130 1733 4133 1816
rect 4138 1813 4141 1846
rect 4146 1803 4149 1926
rect 4154 1793 4157 2143
rect 4082 1673 4093 1676
rect 3978 1546 3981 1616
rect 3986 1593 3989 1606
rect 3994 1553 3997 1626
rect 4002 1583 4005 1606
rect 3978 1543 3997 1546
rect 3970 1356 3973 1526
rect 3978 1496 3981 1536
rect 3986 1513 3989 1526
rect 3978 1493 3985 1496
rect 3982 1416 3985 1493
rect 3982 1413 3989 1416
rect 3978 1393 3981 1406
rect 3954 1353 3973 1356
rect 3898 1293 3917 1296
rect 3914 1236 3917 1293
rect 3906 1233 3917 1236
rect 3854 1163 3861 1166
rect 3850 1133 3853 1146
rect 3858 1123 3861 1163
rect 3866 1133 3869 1186
rect 3882 1173 3885 1206
rect 3898 1156 3901 1176
rect 3894 1153 3901 1156
rect 3874 1113 3877 1136
rect 3882 1123 3885 1136
rect 3822 1103 3837 1106
rect 3810 1093 3821 1096
rect 3786 946 3789 1046
rect 3810 993 3813 1016
rect 3778 943 3789 946
rect 3762 863 3765 926
rect 3770 883 3773 916
rect 3778 846 3781 943
rect 3786 873 3789 936
rect 3778 843 3789 846
rect 3762 756 3765 836
rect 3770 813 3773 826
rect 3778 823 3781 836
rect 3730 703 3749 706
rect 3754 753 3765 756
rect 3714 633 3725 636
rect 3714 603 3717 626
rect 3690 533 3693 546
rect 3698 523 3701 556
rect 3674 513 3685 516
rect 3674 446 3677 513
rect 3706 496 3709 596
rect 3666 443 3677 446
rect 3690 493 3709 496
rect 3658 373 3661 406
rect 3658 333 3661 366
rect 3578 323 3597 326
rect 3562 236 3565 246
rect 3522 233 3565 236
rect 3522 213 3525 233
rect 3530 213 3533 226
rect 3530 173 3533 206
rect 3506 123 3509 136
rect 3538 133 3541 206
rect 3546 196 3549 216
rect 3554 203 3557 216
rect 3562 213 3565 233
rect 3578 213 3581 306
rect 3594 213 3597 256
rect 3562 196 3565 206
rect 3602 203 3605 326
rect 3618 323 3629 326
rect 3610 213 3613 226
rect 3618 206 3621 323
rect 3626 313 3637 316
rect 3642 313 3645 326
rect 3650 323 3661 326
rect 3634 303 3637 313
rect 3650 303 3653 316
rect 3634 213 3653 216
rect 3658 213 3661 323
rect 3666 293 3669 443
rect 3682 413 3685 426
rect 3674 393 3677 406
rect 3674 333 3677 346
rect 3682 316 3685 336
rect 3690 333 3693 493
rect 3722 456 3725 633
rect 3730 593 3733 703
rect 3754 673 3757 753
rect 3770 733 3773 756
rect 3786 753 3789 843
rect 3794 826 3797 976
rect 3818 973 3821 1093
rect 3834 1056 3837 1103
rect 3830 1053 3837 1056
rect 3830 976 3833 1053
rect 3830 973 3837 976
rect 3802 833 3805 936
rect 3818 933 3821 966
rect 3826 926 3829 936
rect 3810 923 3829 926
rect 3826 913 3829 923
rect 3794 823 3801 826
rect 3798 766 3801 823
rect 3798 763 3805 766
rect 3738 613 3749 616
rect 3754 613 3757 656
rect 3746 553 3749 606
rect 3762 563 3765 636
rect 3770 623 3773 726
rect 3794 723 3797 746
rect 3802 723 3805 763
rect 3810 756 3813 906
rect 3834 903 3837 973
rect 3858 936 3861 1056
rect 3874 1026 3877 1106
rect 3894 1096 3897 1153
rect 3906 1103 3909 1233
rect 3914 1133 3917 1186
rect 3922 1176 3925 1216
rect 3930 1193 3933 1216
rect 3922 1173 3929 1176
rect 3926 1126 3929 1173
rect 3922 1123 3929 1126
rect 3894 1093 3901 1096
rect 3870 1023 3877 1026
rect 3870 966 3873 1023
rect 3870 963 3877 966
rect 3874 946 3877 963
rect 3882 953 3885 1016
rect 3898 1003 3901 1093
rect 3922 1046 3925 1123
rect 3922 1043 3929 1046
rect 3926 996 3929 1043
rect 3922 993 3929 996
rect 3874 943 3885 946
rect 3850 933 3861 936
rect 3850 886 3853 933
rect 3866 893 3869 926
rect 3850 883 3869 886
rect 3826 813 3829 826
rect 3818 773 3821 806
rect 3810 753 3817 756
rect 3778 573 3781 636
rect 3786 613 3789 626
rect 3794 613 3797 626
rect 3738 543 3749 546
rect 3746 523 3749 543
rect 3802 456 3805 716
rect 3814 636 3817 753
rect 3834 733 3837 866
rect 3842 786 3845 846
rect 3850 803 3853 816
rect 3858 793 3861 806
rect 3866 786 3869 883
rect 3882 843 3885 943
rect 3890 913 3893 926
rect 3914 913 3917 936
rect 3842 783 3849 786
rect 3846 726 3849 783
rect 3810 633 3817 636
rect 3842 723 3849 726
rect 3858 783 3869 786
rect 3810 613 3813 633
rect 3826 613 3829 626
rect 3818 583 3821 606
rect 3834 603 3837 616
rect 3842 576 3845 723
rect 3858 713 3861 783
rect 3866 753 3869 766
rect 3874 746 3877 806
rect 3882 763 3885 786
rect 3890 753 3893 816
rect 3914 813 3917 836
rect 3866 743 3877 746
rect 3866 723 3869 743
rect 3874 723 3877 736
rect 3890 733 3893 746
rect 3882 676 3885 726
rect 3898 723 3901 776
rect 3914 766 3917 806
rect 3906 763 3917 766
rect 3906 716 3909 763
rect 3898 713 3909 716
rect 3882 673 3893 676
rect 3850 583 3853 616
rect 3858 593 3861 606
rect 3842 573 3853 576
rect 3818 523 3821 556
rect 3706 453 3725 456
rect 3794 453 3805 456
rect 3674 313 3685 316
rect 3666 213 3669 256
rect 3610 203 3621 206
rect 3546 193 3565 196
rect 3554 123 3557 193
rect 3594 133 3597 156
rect 3618 103 3621 203
rect 3626 123 3629 206
rect 3634 203 3645 206
rect 3666 156 3669 206
rect 3674 203 3677 313
rect 3682 213 3685 306
rect 3690 203 3693 256
rect 3698 213 3701 386
rect 3706 376 3709 453
rect 3730 393 3733 416
rect 3706 373 3717 376
rect 3714 333 3717 373
rect 3794 366 3797 453
rect 3810 413 3813 426
rect 3730 343 3741 346
rect 3738 323 3741 343
rect 3698 196 3701 206
rect 3706 203 3709 256
rect 3714 196 3717 226
rect 3722 213 3733 216
rect 3738 213 3741 226
rect 3746 206 3749 366
rect 3794 363 3805 366
rect 3802 343 3805 363
rect 3818 353 3821 446
rect 3810 323 3813 336
rect 3762 213 3765 246
rect 3778 213 3781 316
rect 3698 193 3717 196
rect 3666 153 3677 156
rect 3674 123 3677 153
rect 3698 133 3701 146
rect 3722 123 3725 206
rect 3738 203 3749 206
rect 3762 126 3765 206
rect 3770 193 3773 206
rect 3786 203 3789 226
rect 3802 213 3805 306
rect 3810 203 3813 316
rect 3818 213 3821 236
rect 3826 223 3829 526
rect 3842 456 3845 536
rect 3850 533 3853 573
rect 3866 546 3869 606
rect 3874 583 3877 616
rect 3882 603 3885 626
rect 3866 543 3877 546
rect 3858 533 3869 536
rect 3858 523 3869 526
rect 3842 453 3853 456
rect 3842 413 3845 436
rect 3850 413 3853 453
rect 3858 406 3861 516
rect 3874 506 3877 543
rect 3834 393 3837 406
rect 3842 303 3845 406
rect 3850 403 3861 406
rect 3870 503 3877 506
rect 3850 363 3853 403
rect 3870 356 3873 503
rect 3870 353 3877 356
rect 3858 333 3869 336
rect 3858 323 3869 326
rect 3874 263 3877 353
rect 3826 203 3829 216
rect 3834 213 3837 256
rect 3882 253 3885 576
rect 3890 553 3893 673
rect 3898 583 3901 713
rect 3914 696 3917 736
rect 3910 693 3917 696
rect 3910 636 3913 693
rect 3910 633 3917 636
rect 3906 593 3909 616
rect 3890 526 3893 536
rect 3898 533 3901 566
rect 3914 563 3917 633
rect 3922 573 3925 993
rect 3938 956 3941 1156
rect 3946 1103 3949 1336
rect 3954 1333 3957 1353
rect 3954 1073 3957 1306
rect 3962 1183 3965 1336
rect 3962 1066 3965 1136
rect 3970 1123 3973 1326
rect 3978 1263 3981 1376
rect 3978 1213 3981 1256
rect 3978 1133 3981 1206
rect 3946 1063 3965 1066
rect 3946 1013 3949 1063
rect 3978 1056 3981 1126
rect 3986 1113 3989 1413
rect 3994 1323 3997 1543
rect 4002 1533 4005 1546
rect 4010 1433 4013 1526
rect 4018 1496 4021 1586
rect 4034 1533 4037 1576
rect 4050 1573 4053 1606
rect 4074 1593 4077 1616
rect 4090 1586 4093 1673
rect 4146 1613 4149 1626
rect 4082 1583 4093 1586
rect 4058 1523 4061 1546
rect 4018 1493 4029 1496
rect 4026 1436 4029 1493
rect 4074 1486 4077 1506
rect 4018 1433 4029 1436
rect 4066 1483 4077 1486
rect 4018 1413 4021 1433
rect 4066 1426 4069 1483
rect 4082 1436 4085 1583
rect 4082 1433 4093 1436
rect 4066 1423 4077 1426
rect 4026 1413 4045 1416
rect 4002 1363 4005 1406
rect 4018 1343 4021 1406
rect 4026 1403 4029 1413
rect 4050 1403 4053 1416
rect 4002 1333 4013 1336
rect 4002 1323 4013 1326
rect 4018 1313 4021 1336
rect 4034 1293 4037 1386
rect 4058 1323 4061 1346
rect 4066 1313 4069 1406
rect 3994 1213 3997 1236
rect 4002 1153 4005 1206
rect 4010 1203 4013 1256
rect 4026 1213 4029 1226
rect 4018 1193 4021 1206
rect 4010 1146 4013 1166
rect 4002 1143 4013 1146
rect 3994 1123 3997 1136
rect 3978 1053 3989 1056
rect 3938 953 3949 956
rect 3930 733 3933 946
rect 3946 866 3949 953
rect 3938 863 3949 866
rect 3938 763 3941 863
rect 3962 803 3965 1016
rect 3986 1006 3989 1053
rect 3994 1013 3997 1076
rect 4002 1013 4005 1143
rect 4010 1106 4013 1136
rect 4018 1133 4021 1146
rect 4026 1113 4029 1126
rect 4010 1103 4017 1106
rect 4014 1036 4017 1103
rect 4010 1033 4017 1036
rect 4010 1013 4013 1033
rect 4026 1013 4029 1106
rect 3986 1003 3993 1006
rect 3970 906 3973 926
rect 3978 923 3981 936
rect 3970 903 3981 906
rect 3978 836 3981 903
rect 3970 833 3981 836
rect 3970 813 3973 833
rect 3990 826 3993 1003
rect 4002 933 4005 1006
rect 4018 993 4021 1006
rect 4034 1003 4037 1206
rect 4066 1203 4069 1296
rect 4074 1253 4077 1423
rect 4090 1386 4093 1433
rect 4106 1406 4109 1566
rect 4130 1513 4133 1526
rect 4082 1383 4093 1386
rect 4102 1403 4109 1406
rect 4082 1246 4085 1383
rect 4102 1356 4105 1403
rect 4102 1353 4109 1356
rect 4082 1243 4093 1246
rect 4050 1003 4053 1176
rect 4074 1123 4077 1146
rect 4074 993 4077 1016
rect 3990 823 3997 826
rect 3978 773 3981 816
rect 3946 633 3949 756
rect 3970 723 3973 746
rect 3978 656 3981 766
rect 3986 733 3989 806
rect 3994 783 3997 823
rect 4002 776 4005 926
rect 4018 823 4021 936
rect 4026 913 4029 926
rect 4034 846 4037 936
rect 4042 913 4045 926
rect 4090 856 4093 1243
rect 4098 1213 4101 1336
rect 4106 1296 4109 1353
rect 4114 1323 4117 1396
rect 4122 1316 4125 1326
rect 4114 1313 4125 1316
rect 4106 1293 4113 1296
rect 4110 1186 4113 1293
rect 4146 1213 4149 1336
rect 4106 1183 4113 1186
rect 4106 1163 4109 1183
rect 4122 1123 4133 1126
rect 4146 1013 4149 1026
rect 4026 843 4037 846
rect 3994 773 4005 776
rect 3994 686 3997 773
rect 4010 743 4013 806
rect 4018 793 4021 816
rect 4026 746 4029 843
rect 4042 783 4045 856
rect 4082 853 4093 856
rect 4066 813 4069 826
rect 4026 743 4037 746
rect 4026 723 4029 736
rect 3994 683 4013 686
rect 3954 653 3981 656
rect 3938 613 3941 626
rect 3954 606 3957 653
rect 3946 603 3957 606
rect 3914 553 3925 556
rect 3914 533 3917 546
rect 3890 523 3909 526
rect 3906 393 3909 416
rect 3850 213 3853 226
rect 3866 213 3885 216
rect 3890 213 3893 386
rect 3898 323 3901 336
rect 3906 303 3909 346
rect 3914 323 3917 436
rect 3922 383 3925 553
rect 3930 373 3933 556
rect 3946 513 3949 603
rect 3962 436 3965 636
rect 3986 603 3989 636
rect 4002 583 4005 606
rect 4010 566 4013 683
rect 4018 613 4029 616
rect 4018 593 4021 606
rect 4002 563 4013 566
rect 3986 523 3989 546
rect 4002 456 4005 563
rect 4026 486 4029 536
rect 4018 483 4029 486
rect 4002 453 4013 456
rect 3962 433 3985 436
rect 3922 333 3925 346
rect 3938 333 3941 356
rect 3954 333 3957 406
rect 3970 373 3973 406
rect 3982 366 3985 433
rect 3994 396 3997 436
rect 4010 433 4013 453
rect 4018 413 4021 483
rect 4034 476 4037 743
rect 4066 656 4069 786
rect 4082 776 4085 853
rect 4122 813 4125 926
rect 4130 793 4133 816
rect 4082 773 4093 776
rect 4090 756 4093 773
rect 4090 753 4101 756
rect 4090 723 4093 746
rect 4098 656 4101 753
rect 4146 723 4149 806
rect 4050 653 4069 656
rect 4090 653 4101 656
rect 4050 536 4053 653
rect 4074 593 4077 616
rect 4090 576 4093 653
rect 4146 613 4149 626
rect 4090 573 4101 576
rect 4098 553 4101 573
rect 4026 473 4037 476
rect 4042 533 4053 536
rect 3994 393 4001 396
rect 4010 393 4013 406
rect 3982 363 3989 366
rect 3842 203 3853 206
rect 3810 133 3813 146
rect 3762 123 3781 126
rect 3858 123 3861 206
rect 3866 193 3869 213
rect 3874 203 3885 206
rect 3890 123 3893 206
rect 3898 193 3901 276
rect 3906 203 3909 266
rect 3922 213 3925 326
rect 3930 313 3933 326
rect 3978 323 3981 346
rect 3938 213 3949 216
rect 3962 213 3965 236
rect 3970 213 3973 226
rect 3978 206 3981 306
rect 3914 153 3917 206
rect 3922 203 3933 206
rect 3922 133 3925 146
rect 3946 123 3949 156
rect 3954 133 3957 206
rect 3970 203 3981 206
rect 3970 183 3973 203
rect 3986 143 3989 363
rect 3998 236 4001 393
rect 4026 326 4029 473
rect 4042 383 4045 533
rect 4050 523 4061 526
rect 4066 523 4069 536
rect 4146 506 4149 526
rect 4138 503 4149 506
rect 4138 436 4141 503
rect 4138 433 4149 436
rect 4058 376 4061 406
rect 4082 393 4085 416
rect 4146 413 4149 433
rect 4058 373 4069 376
rect 3994 233 4001 236
rect 4018 323 4029 326
rect 3994 213 3997 233
rect 4002 123 4005 206
rect 4010 193 4013 206
rect 4018 203 4021 323
rect 4026 203 4029 316
rect 4034 296 4037 336
rect 4066 333 4069 373
rect 4042 323 4053 326
rect 4090 313 4093 326
rect 4034 293 4045 296
rect 4042 246 4045 293
rect 4034 243 4045 246
rect 4034 213 4037 243
rect 4042 213 4053 216
rect 4082 213 4085 226
rect 4146 213 4149 326
rect 4034 203 4045 206
rect 4034 133 4037 146
rect 4058 123 4061 136
rect 4082 133 4085 206
rect 4114 123 4117 136
rect 4167 37 4187 4103
rect 4191 13 4211 4127
rect 4218 2603 4221 2796
<< metal3 >>
rect 3305 4062 3334 4067
rect 2001 4052 2030 4057
rect 2017 4042 2166 4047
rect 1969 4032 2022 4037
rect 249 4022 294 4027
rect 393 4022 438 4027
rect 513 4022 558 4027
rect 849 4022 894 4027
rect 1177 4022 1222 4027
rect 1289 4022 1334 4027
rect 1545 4022 1590 4027
rect 1657 4022 1702 4027
rect 2289 4022 2446 4027
rect 2689 4022 2726 4027
rect 2817 4022 2854 4027
rect 2945 4022 2982 4027
rect 3097 4022 3182 4027
rect 3281 4022 3342 4027
rect 3353 4022 3462 4027
rect 3777 4022 3902 4027
rect 1857 4012 1894 4017
rect 2097 4012 2142 4017
rect 129 4002 174 4007
rect 233 4002 342 4007
rect 913 4002 958 4007
rect 2201 4002 2246 4007
rect 241 3992 302 3997
rect 529 3992 638 3997
rect 809 3992 1046 3997
rect 1169 3992 1222 3997
rect 1377 3992 1478 3997
rect 1497 3992 1774 3997
rect 1857 3992 2190 3997
rect 321 3987 414 3992
rect 2185 3987 2190 3992
rect 2289 3987 2294 4022
rect 2441 4007 2446 4022
rect 3097 4017 3102 4022
rect 2657 4012 3102 4017
rect 3177 4017 3182 4022
rect 3177 4012 3254 4017
rect 3513 4012 3758 4017
rect 2441 4002 2646 4007
rect 2641 3997 2646 4002
rect 2713 4002 2742 4007
rect 2841 4002 2886 4007
rect 2969 4002 3030 4007
rect 3105 4002 3166 4007
rect 3393 4002 3470 4007
rect 2713 3997 2718 4002
rect 3393 3997 3398 4002
rect 2313 3992 2342 3997
rect 2361 3992 2430 3997
rect 2641 3992 2718 3997
rect 2777 3992 2806 3997
rect 2833 3992 2854 3997
rect 3265 3992 3286 3997
rect 3297 3992 3398 3997
rect 3465 3997 3470 4002
rect 3513 3997 3518 4012
rect 3465 3992 3518 3997
rect 3753 3997 3758 4012
rect 3753 3992 3782 3997
rect 3825 3992 3870 3997
rect 3993 3992 4038 3997
rect 161 3982 326 3987
rect 409 3982 438 3987
rect 1073 3982 1198 3987
rect 2185 3982 2294 3987
rect 2417 3982 2438 3987
rect 2873 3982 2966 3987
rect 737 3977 806 3982
rect 2873 3977 2878 3982
rect 265 3972 414 3977
rect 713 3972 742 3977
rect 801 3972 862 3977
rect 1281 3972 1326 3977
rect 1849 3972 1886 3977
rect 1913 3972 1958 3977
rect 2337 3972 2590 3977
rect 2825 3972 2878 3977
rect 2961 3977 2966 3982
rect 3113 3982 3222 3987
rect 3249 3982 3286 3987
rect 3425 3982 3454 3987
rect 3489 3982 4014 3987
rect 3113 3977 3118 3982
rect 2961 3972 2990 3977
rect 3057 3972 3118 3977
rect 3217 3977 3222 3982
rect 3281 3977 3430 3982
rect 3217 3972 3262 3977
rect 3545 3972 3894 3977
rect 3057 3967 3062 3972
rect 345 3962 430 3967
rect 625 3962 790 3967
rect 1089 3962 1342 3967
rect 1833 3962 1886 3967
rect 1969 3962 2078 3967
rect 2193 3962 2238 3967
rect 2785 3962 3062 3967
rect 3073 3962 3302 3967
rect 3361 3962 3742 3967
rect 3873 3962 3934 3967
rect 3953 3962 4022 3967
rect 625 3957 630 3962
rect 1881 3957 1974 3962
rect 3361 3957 3366 3962
rect 3737 3957 3878 3962
rect 3953 3957 3958 3962
rect 385 3952 494 3957
rect 553 3952 630 3957
rect 641 3952 718 3957
rect 825 3952 854 3957
rect 881 3952 982 3957
rect 1241 3952 1278 3957
rect 1577 3952 1670 3957
rect 1705 3952 1766 3957
rect 2737 3952 2870 3957
rect 2985 3952 3030 3957
rect 1785 3947 1862 3952
rect 3025 3947 3030 3952
rect 3097 3952 3294 3957
rect 3337 3952 3366 3957
rect 3513 3952 3558 3957
rect 3585 3952 3718 3957
rect 3897 3952 3958 3957
rect 4017 3957 4022 3962
rect 4017 3952 4070 3957
rect 3097 3947 3102 3952
rect 81 3942 198 3947
rect 289 3942 358 3947
rect 497 3942 822 3947
rect 1033 3942 1206 3947
rect 1273 3942 1302 3947
rect 1313 3942 1390 3947
rect 1537 3942 1590 3947
rect 1745 3942 1790 3947
rect 1857 3942 1942 3947
rect 2001 3942 2070 3947
rect 2081 3942 2134 3947
rect 2313 3942 2374 3947
rect 2393 3942 2558 3947
rect 2673 3942 2766 3947
rect 2777 3942 3006 3947
rect 3025 3942 3102 3947
rect 3169 3942 3342 3947
rect 3369 3942 3550 3947
rect 3569 3942 3598 3947
rect 3729 3942 3766 3947
rect 3857 3942 3886 3947
rect 3921 3942 4006 3947
rect 3921 3937 3926 3942
rect 417 3932 950 3937
rect 961 3932 998 3937
rect 1169 3932 1254 3937
rect 1265 3932 1470 3937
rect 1553 3932 1846 3937
rect 2209 3932 2918 3937
rect 3521 3932 3638 3937
rect 3705 3932 3926 3937
rect 3985 3932 4014 3937
rect 2961 3927 3030 3932
rect 3265 3927 3382 3932
rect 4009 3927 4014 3932
rect 4081 3932 4118 3937
rect 4081 3927 4086 3932
rect 361 3922 470 3927
rect 505 3922 606 3927
rect 617 3922 694 3927
rect 737 3922 902 3927
rect 1049 3922 1150 3927
rect 1193 3922 1406 3927
rect 1697 3922 1814 3927
rect 2353 3922 2838 3927
rect 2929 3922 2966 3927
rect 3025 3922 3270 3927
rect 3377 3922 3750 3927
rect 1529 3917 1646 3922
rect 1697 3917 1702 3922
rect 273 3912 398 3917
rect 417 3912 894 3917
rect 1017 3912 1182 3917
rect 1193 3912 1270 3917
rect 1337 3912 1430 3917
rect 1505 3912 1534 3917
rect 1641 3912 1702 3917
rect 1721 3912 1766 3917
rect 2113 3912 2294 3917
rect 2561 3912 2566 3922
rect 2833 3917 2934 3922
rect 3745 3917 3750 3922
rect 3857 3922 3926 3927
rect 4009 3922 4086 3927
rect 3857 3917 3862 3922
rect 2585 3912 2702 3917
rect 2769 3912 2814 3917
rect 2977 3912 3014 3917
rect 3281 3912 3390 3917
rect 3401 3912 3446 3917
rect 3553 3912 3598 3917
rect 3689 3912 3726 3917
rect 3745 3912 3862 3917
rect 3889 3912 3974 3917
rect 321 3902 390 3907
rect 401 3902 870 3907
rect 937 3902 1030 3907
rect 1065 3902 1238 3907
rect 1297 3902 1526 3907
rect 1537 3902 1606 3907
rect 1617 3902 1646 3907
rect 1777 3902 1838 3907
rect 2249 3902 2294 3907
rect 1641 3897 1782 3902
rect 2289 3897 2294 3902
rect 2393 3902 2446 3907
rect 2593 3902 2630 3907
rect 2705 3902 2790 3907
rect 2873 3902 2958 3907
rect 3393 3902 3422 3907
rect 2393 3897 2398 3902
rect 2873 3897 2878 3902
rect 553 3892 630 3897
rect 697 3892 734 3897
rect 753 3892 934 3897
rect 1001 3892 1566 3897
rect 2193 3892 2270 3897
rect 2289 3892 2398 3897
rect 2417 3892 2878 3897
rect 2953 3897 2958 3902
rect 3441 3897 3558 3902
rect 2953 3892 3118 3897
rect 3137 3892 3262 3897
rect 3337 3892 3446 3897
rect 3553 3892 3750 3897
rect 3761 3892 3854 3897
rect 3137 3887 3142 3892
rect 449 3882 1286 3887
rect 1361 3882 1470 3887
rect 1513 3882 1550 3887
rect 1601 3882 2182 3887
rect 2889 3882 3038 3887
rect 3057 3882 3142 3887
rect 3257 3887 3262 3892
rect 3257 3882 3374 3887
rect 3385 3882 3542 3887
rect 3657 3882 3822 3887
rect 305 3872 430 3877
rect 601 3872 662 3877
rect 705 3872 982 3877
rect 1025 3872 1222 3877
rect 1249 3872 1534 3877
rect 305 3867 310 3872
rect 281 3862 310 3867
rect 425 3867 430 3872
rect 1217 3867 1222 3872
rect 1601 3867 1606 3882
rect 2577 3877 2870 3882
rect 3057 3877 3062 3882
rect 3537 3877 3662 3882
rect 2553 3872 2582 3877
rect 2865 3872 3062 3877
rect 3161 3872 3230 3877
rect 3241 3872 3518 3877
rect 3513 3867 3518 3872
rect 3689 3872 3790 3877
rect 3689 3867 3694 3872
rect 425 3862 942 3867
rect 1217 3862 1606 3867
rect 2185 3862 2254 3867
rect 2297 3862 2438 3867
rect 969 3857 1126 3862
rect 2297 3857 2302 3862
rect 825 3852 974 3857
rect 1121 3852 1622 3857
rect 1641 3852 1902 3857
rect 2273 3852 2302 3857
rect 2433 3857 2438 3862
rect 2609 3862 3190 3867
rect 2609 3857 2614 3862
rect 3185 3857 3190 3862
rect 3345 3862 3494 3867
rect 3513 3862 3694 3867
rect 3345 3857 3350 3862
rect 2433 3852 2614 3857
rect 2625 3852 3078 3857
rect 3185 3852 3350 3857
rect 3713 3852 3774 3857
rect 345 3847 502 3852
rect 1641 3847 1646 3852
rect 185 3842 262 3847
rect 321 3842 350 3847
rect 497 3842 790 3847
rect 985 3842 1110 3847
rect 1289 3842 1462 3847
rect 1521 3842 1646 3847
rect 1897 3847 1902 3852
rect 1897 3842 1926 3847
rect 1969 3842 2054 3847
rect 2297 3842 2422 3847
rect 2649 3842 2742 3847
rect 3097 3842 3166 3847
rect 3577 3842 3694 3847
rect 3937 3842 4062 3847
rect 185 3837 190 3842
rect 129 3832 190 3837
rect 257 3837 262 3842
rect 785 3837 990 3842
rect 1521 3837 1526 3842
rect 1969 3837 1974 3842
rect 2761 3837 2926 3842
rect 2969 3837 3046 3842
rect 3097 3837 3102 3842
rect 257 3832 486 3837
rect 1009 3832 1054 3837
rect 1089 3832 1134 3837
rect 1329 3832 1526 3837
rect 1537 3832 1654 3837
rect 1665 3832 1886 3837
rect 1945 3832 1974 3837
rect 1993 3832 2046 3837
rect 2241 3832 2662 3837
rect 2673 3832 2766 3837
rect 2921 3832 2974 3837
rect 3041 3832 3102 3837
rect 3161 3837 3166 3842
rect 3937 3837 3942 3842
rect 3161 3832 3390 3837
rect 3505 3832 3574 3837
rect 3593 3832 3758 3837
rect 3817 3832 3902 3837
rect 1329 3827 1334 3832
rect 1665 3827 1670 3832
rect 1881 3827 1950 3832
rect 2657 3827 2662 3832
rect 3817 3827 3822 3832
rect 137 3822 166 3827
rect 201 3822 326 3827
rect 377 3822 422 3827
rect 433 3822 494 3827
rect 625 3822 670 3827
rect 753 3822 798 3827
rect 865 3822 974 3827
rect 1057 3822 1110 3827
rect 1201 3822 1334 3827
rect 1401 3822 1446 3827
rect 1465 3822 1494 3827
rect 1585 3822 1670 3827
rect 1681 3822 1726 3827
rect 1793 3822 1838 3827
rect 2009 3822 2038 3827
rect 2121 3822 2142 3827
rect 2265 3822 2406 3827
rect 2657 3822 2774 3827
rect 2833 3822 2910 3827
rect 2985 3822 3030 3827
rect 3113 3822 3150 3827
rect 3273 3822 3302 3827
rect 3409 3822 3438 3827
rect 3561 3822 3614 3827
rect 3633 3822 3678 3827
rect 3689 3822 3742 3827
rect 3793 3822 3822 3827
rect 3897 3827 3902 3832
rect 3921 3832 3942 3837
rect 4057 3837 4062 3842
rect 4057 3832 4086 3837
rect 3921 3827 3926 3832
rect 3897 3822 3926 3827
rect 3937 3822 4062 3827
rect 1489 3817 1590 3822
rect 193 3812 294 3817
rect 353 3812 462 3817
rect 801 3812 830 3817
rect 929 3812 1246 3817
rect 1609 3812 1702 3817
rect 1817 3812 1878 3817
rect 2257 3812 2318 3817
rect 2393 3812 2438 3817
rect 2449 3812 2678 3817
rect 2689 3812 2758 3817
rect 3033 3812 3174 3817
rect 3289 3812 3502 3817
rect 825 3807 934 3812
rect 1265 3807 1374 3812
rect 2449 3807 2454 3812
rect 473 3802 510 3807
rect 761 3802 798 3807
rect 953 3802 1270 3807
rect 1369 3802 1590 3807
rect 2337 3802 2454 3807
rect 2673 3807 2678 3812
rect 2673 3802 3366 3807
rect 3393 3802 3430 3807
rect 2337 3797 2342 3802
rect 3361 3797 3366 3802
rect 3449 3797 3566 3802
rect 3585 3797 3590 3817
rect 3601 3812 3646 3817
rect 3705 3812 3734 3817
rect 3745 3812 3774 3817
rect 3833 3812 4014 3817
rect 3729 3807 3734 3812
rect 3769 3807 3838 3812
rect 3617 3802 3662 3807
rect 3713 3802 3734 3807
rect 3969 3802 3998 3807
rect 3969 3797 3974 3802
rect 121 3792 318 3797
rect 529 3792 646 3797
rect 841 3792 942 3797
rect 993 3792 1158 3797
rect 1169 3792 1358 3797
rect 1521 3792 1542 3797
rect 1577 3792 1790 3797
rect 2137 3792 2238 3797
rect 2249 3792 2342 3797
rect 2353 3792 2398 3797
rect 2505 3792 2590 3797
rect 2673 3792 2742 3797
rect 3001 3792 3030 3797
rect 3113 3792 3342 3797
rect 3361 3792 3454 3797
rect 3561 3792 3590 3797
rect 3649 3792 3694 3797
rect 3753 3792 3830 3797
rect 3873 3792 3918 3797
rect 3929 3792 3974 3797
rect 4009 3792 4110 3797
rect 3025 3787 3118 3792
rect 497 3782 526 3787
rect 521 3777 526 3782
rect 657 3782 830 3787
rect 657 3777 662 3782
rect 289 3772 366 3777
rect 521 3772 662 3777
rect 825 3777 830 3782
rect 929 3782 958 3787
rect 1009 3782 1142 3787
rect 1201 3782 1414 3787
rect 1513 3782 1622 3787
rect 1817 3782 1870 3787
rect 2217 3782 2342 3787
rect 2361 3782 2406 3787
rect 2417 3782 2670 3787
rect 2721 3782 2766 3787
rect 2793 3782 2878 3787
rect 2977 3782 3006 3787
rect 929 3777 934 3782
rect 825 3772 934 3777
rect 1137 3777 1142 3782
rect 2337 3777 2342 3782
rect 2417 3777 2422 3782
rect 2793 3777 2798 3782
rect 1137 3772 1278 3777
rect 1449 3772 1550 3777
rect 289 3767 294 3772
rect 105 3762 182 3767
rect 217 3762 294 3767
rect 361 3767 366 3772
rect 1545 3767 1550 3772
rect 1633 3772 2094 3777
rect 2337 3772 2422 3777
rect 2553 3772 2574 3777
rect 2649 3772 2686 3777
rect 2753 3772 2798 3777
rect 2873 3777 2878 3782
rect 3001 3777 3006 3782
rect 3161 3782 3326 3787
rect 3337 3782 3638 3787
rect 3681 3782 3726 3787
rect 3889 3782 4038 3787
rect 3161 3777 3166 3782
rect 3745 3777 3894 3782
rect 2873 3772 2902 3777
rect 3001 3772 3166 3777
rect 3409 3772 3454 3777
rect 3513 3772 3750 3777
rect 3913 3772 3974 3777
rect 4001 3772 4030 3777
rect 1633 3767 1638 3772
rect 3241 3767 3390 3772
rect 361 3762 390 3767
rect 737 3762 806 3767
rect 985 3762 1078 3767
rect 1161 3762 1206 3767
rect 1545 3762 1638 3767
rect 1809 3762 1838 3767
rect 2457 3762 2518 3767
rect 2537 3762 2814 3767
rect 2841 3762 2894 3767
rect 3217 3762 3246 3767
rect 3385 3762 3558 3767
rect 3673 3762 3758 3767
rect 3841 3762 3966 3767
rect 4033 3762 4078 3767
rect 1225 3757 1310 3762
rect 161 3752 478 3757
rect 737 3752 926 3757
rect 969 3752 1046 3757
rect 1057 3752 1110 3757
rect 1193 3752 1230 3757
rect 1305 3752 1526 3757
rect 1777 3752 1854 3757
rect 2049 3752 2142 3757
rect 2329 3752 2382 3757
rect 2393 3752 2454 3757
rect 2577 3752 2646 3757
rect 2785 3752 2886 3757
rect 2897 3752 3518 3757
rect 3673 3752 3710 3757
rect 3753 3752 3814 3757
rect 3833 3752 3894 3757
rect 3913 3752 4094 3757
rect 3809 3747 3814 3752
rect 153 3742 238 3747
rect 345 3742 374 3747
rect 369 3737 374 3742
rect 465 3742 510 3747
rect 537 3742 590 3747
rect 617 3742 726 3747
rect 785 3742 846 3747
rect 977 3742 1014 3747
rect 1081 3742 1110 3747
rect 1153 3742 1294 3747
rect 1617 3742 1774 3747
rect 1873 3742 1926 3747
rect 1937 3742 2038 3747
rect 2105 3742 2206 3747
rect 2225 3742 2406 3747
rect 2505 3742 2550 3747
rect 2561 3742 2606 3747
rect 2649 3742 2758 3747
rect 2825 3742 2886 3747
rect 2897 3742 2934 3747
rect 2945 3742 3006 3747
rect 3129 3742 3174 3747
rect 3265 3742 3294 3747
rect 3313 3742 3398 3747
rect 3465 3742 3542 3747
rect 3553 3742 3590 3747
rect 3633 3742 3710 3747
rect 465 3737 470 3742
rect 369 3732 470 3737
rect 529 3732 822 3737
rect 169 3722 222 3727
rect 289 3722 350 3727
rect 489 3722 646 3727
rect 737 3722 926 3727
rect 1105 3722 1110 3742
rect 1137 3732 1174 3737
rect 1241 3732 1302 3737
rect 2209 3732 2246 3737
rect 2369 3732 2390 3737
rect 2409 3732 2598 3737
rect 2617 3732 2814 3737
rect 2881 3732 3014 3737
rect 3241 3732 3286 3737
rect 1169 3722 1174 3732
rect 1209 3722 1422 3727
rect 641 3717 742 3722
rect 129 3712 174 3717
rect 193 3712 246 3717
rect 257 3712 310 3717
rect 321 3712 342 3717
rect 369 3712 414 3717
rect 513 3712 550 3717
rect 569 3712 622 3717
rect 761 3712 830 3717
rect 1017 3712 1070 3717
rect 1161 3712 1198 3717
rect 1249 3712 1286 3717
rect 1401 3712 1446 3717
rect 1793 3712 1838 3717
rect 2209 3712 2214 3732
rect 2385 3727 2390 3732
rect 2593 3727 2598 3732
rect 2809 3727 2886 3732
rect 3553 3727 3558 3742
rect 3721 3737 3726 3747
rect 3745 3742 3782 3747
rect 3809 3742 3870 3747
rect 3881 3742 3942 3747
rect 4017 3742 4078 3747
rect 3657 3732 3726 3737
rect 3737 3732 3814 3737
rect 3865 3732 3910 3737
rect 3953 3732 3990 3737
rect 3953 3727 3958 3732
rect 2385 3722 2502 3727
rect 2593 3722 2758 3727
rect 2905 3722 2942 3727
rect 3081 3722 3182 3727
rect 3321 3722 3422 3727
rect 3537 3722 3558 3727
rect 3721 3722 3798 3727
rect 3873 3722 3958 3727
rect 2753 3717 2758 3722
rect 2441 3712 2614 3717
rect 2633 3712 2694 3717
rect 2753 3712 2918 3717
rect 2929 3712 3070 3717
rect 3289 3712 3390 3717
rect 3513 3712 3686 3717
rect 3697 3712 3742 3717
rect 3777 3712 3886 3717
rect 3897 3712 3926 3717
rect 3945 3712 3990 3717
rect 4001 3712 4142 3717
rect 2609 3707 2614 3712
rect 2913 3707 2918 3712
rect 3777 3707 3782 3712
rect 201 3702 342 3707
rect 337 3697 342 3702
rect 425 3702 478 3707
rect 425 3697 430 3702
rect 337 3692 430 3697
rect 473 3697 478 3702
rect 561 3702 678 3707
rect 809 3702 886 3707
rect 961 3702 1190 3707
rect 1265 3702 1334 3707
rect 2193 3702 2462 3707
rect 2521 3702 2598 3707
rect 2609 3702 2878 3707
rect 2913 3702 2950 3707
rect 3313 3702 3782 3707
rect 3801 3702 3998 3707
rect 561 3697 566 3702
rect 673 3697 678 3702
rect 2593 3697 2598 3702
rect 473 3692 566 3697
rect 617 3692 654 3697
rect 673 3692 950 3697
rect 945 3687 950 3692
rect 1033 3692 1310 3697
rect 1513 3692 1550 3697
rect 2385 3692 2414 3697
rect 1033 3687 1038 3692
rect 2409 3687 2414 3692
rect 2513 3692 2542 3697
rect 2593 3692 2614 3697
rect 2513 3687 2518 3692
rect 2609 3687 2614 3692
rect 2721 3692 2750 3697
rect 2761 3692 3086 3697
rect 3385 3692 3414 3697
rect 3545 3692 3574 3697
rect 3809 3692 3966 3697
rect 2721 3687 2726 3692
rect 3409 3687 3550 3692
rect 817 3682 854 3687
rect 945 3682 1038 3687
rect 1057 3682 1110 3687
rect 849 3667 854 3682
rect 1057 3667 1062 3682
rect 409 3662 534 3667
rect 553 3662 662 3667
rect 849 3662 1062 3667
rect 1105 3667 1110 3682
rect 1249 3682 1278 3687
rect 1521 3682 1550 3687
rect 2409 3682 2518 3687
rect 2537 3682 2574 3687
rect 2609 3682 2726 3687
rect 2825 3682 2982 3687
rect 3793 3682 3854 3687
rect 3897 3682 3974 3687
rect 1249 3667 1254 3682
rect 3001 3677 3134 3682
rect 2873 3672 3006 3677
rect 3129 3672 3158 3677
rect 3177 3672 3254 3677
rect 3177 3667 3182 3672
rect 1105 3662 1254 3667
rect 1273 3662 1814 3667
rect 2145 3662 2230 3667
rect 2665 3662 2750 3667
rect 2809 3662 3182 3667
rect 3249 3667 3254 3672
rect 3393 3672 3494 3677
rect 3561 3672 4014 3677
rect 3393 3667 3398 3672
rect 3249 3662 3398 3667
rect 3489 3667 3494 3672
rect 3489 3662 3614 3667
rect 3825 3662 3950 3667
rect 553 3657 558 3662
rect 481 3652 558 3657
rect 657 3657 662 3662
rect 2665 3657 2670 3662
rect 657 3652 726 3657
rect 1777 3652 1798 3657
rect 2529 3652 2670 3657
rect 2745 3657 2750 3662
rect 2745 3652 2774 3657
rect 2793 3652 3294 3657
rect 3329 3652 3366 3657
rect 3417 3652 3478 3657
rect 3633 3652 3806 3657
rect 3633 3647 3638 3652
rect 3801 3647 3982 3652
rect 529 3642 638 3647
rect 777 3642 830 3647
rect 1089 3642 1350 3647
rect 1369 3642 1454 3647
rect 1369 3637 1374 3642
rect 601 3632 694 3637
rect 705 3632 798 3637
rect 945 3632 1150 3637
rect 1305 3632 1374 3637
rect 1449 3637 1454 3642
rect 1577 3642 1726 3647
rect 1745 3642 1886 3647
rect 1897 3642 1926 3647
rect 2409 3642 2502 3647
rect 2521 3642 2662 3647
rect 2777 3642 2838 3647
rect 2921 3642 3038 3647
rect 3049 3642 3126 3647
rect 3185 3642 3342 3647
rect 3441 3642 3638 3647
rect 3977 3642 4070 3647
rect 1577 3637 1582 3642
rect 1449 3632 1486 3637
rect 1553 3632 1582 3637
rect 1721 3637 1726 3642
rect 2497 3637 2502 3642
rect 2833 3637 2926 3642
rect 3673 3637 3742 3642
rect 1721 3632 1958 3637
rect 1985 3632 2006 3637
rect 2177 3632 2238 3637
rect 2377 3632 2478 3637
rect 2497 3632 2534 3637
rect 2545 3632 2814 3637
rect 2945 3632 3318 3637
rect 3649 3632 3678 3637
rect 3737 3632 3966 3637
rect 689 3627 694 3632
rect 241 3622 286 3627
rect 441 3622 502 3627
rect 577 3622 678 3627
rect 689 3622 790 3627
rect 801 3622 846 3627
rect 1025 3622 1070 3627
rect 785 3617 790 3622
rect 1089 3617 1094 3627
rect 1321 3622 1382 3627
rect 1393 3622 1438 3627
rect 1561 3622 1782 3627
rect 1801 3622 1846 3627
rect 1889 3622 1934 3627
rect 1945 3622 1990 3627
rect 2177 3622 2214 3627
rect 265 3612 398 3617
rect 641 3612 718 3617
rect 785 3612 1094 3617
rect 1113 3612 1158 3617
rect 1217 3612 1414 3617
rect 1537 3612 1582 3617
rect 1593 3612 1630 3617
rect 417 3607 550 3612
rect 1857 3607 1862 3617
rect 1881 3612 1910 3617
rect 2009 3612 2038 3617
rect 2169 3612 2206 3617
rect 2321 3612 2390 3617
rect 1905 3607 2014 3612
rect 129 3602 174 3607
rect 289 3602 422 3607
rect 545 3602 622 3607
rect 697 3602 742 3607
rect 961 3602 1222 3607
rect 1737 3602 1830 3607
rect 1857 3602 1878 3607
rect 2153 3602 2230 3607
rect 2337 3602 2446 3607
rect 2481 3602 2486 3627
rect 2577 3622 2606 3627
rect 2697 3622 2822 3627
rect 2977 3622 2998 3627
rect 3057 3617 3062 3627
rect 3153 3622 3190 3627
rect 3233 3622 3262 3627
rect 3345 3622 3454 3627
rect 3497 3622 3726 3627
rect 3937 3622 4054 3627
rect 2505 3612 2694 3617
rect 2729 3612 2766 3617
rect 2777 3612 2854 3617
rect 3057 3612 3126 3617
rect 3137 3612 3182 3617
rect 2873 3607 2990 3612
rect 2673 3602 2878 3607
rect 2985 3602 3014 3607
rect 3233 3602 3238 3622
rect 3721 3617 3726 3622
rect 3833 3617 3942 3622
rect 3257 3612 3302 3617
rect 3425 3612 3526 3617
rect 3673 3612 3702 3617
rect 3721 3612 3838 3617
rect 3961 3612 4014 3617
rect 3521 3607 3678 3612
rect 3449 3602 3502 3607
rect 3857 3602 3934 3607
rect 1217 3597 1518 3602
rect 2225 3597 2230 3602
rect 2673 3597 2678 3602
rect 81 3592 150 3597
rect 273 3592 358 3597
rect 377 3592 478 3597
rect 497 3592 534 3597
rect 761 3592 814 3597
rect 1057 3592 1134 3597
rect 1177 3592 1198 3597
rect 1513 3592 1542 3597
rect 1809 3592 1966 3597
rect 2113 3592 2206 3597
rect 2225 3592 2254 3597
rect 2369 3592 2398 3597
rect 2473 3592 2502 3597
rect 2569 3592 2598 3597
rect 2657 3592 2678 3597
rect 2689 3592 2734 3597
rect 2769 3592 2870 3597
rect 2921 3592 2966 3597
rect 3057 3592 3086 3597
rect 3105 3592 3150 3597
rect 3225 3592 3270 3597
rect 3369 3592 3446 3597
rect 3473 3592 3590 3597
rect 3633 3592 3718 3597
rect 3777 3592 3806 3597
rect 3865 3592 3894 3597
rect 4033 3592 4094 3597
rect 353 3587 358 3592
rect 2865 3587 2870 3592
rect 353 3582 470 3587
rect 553 3582 670 3587
rect 689 3582 910 3587
rect 921 3582 1582 3587
rect 1873 3582 1942 3587
rect 2185 3582 2270 3587
rect 2329 3582 2390 3587
rect 2441 3582 2646 3587
rect 2657 3582 2686 3587
rect 2737 3582 2846 3587
rect 2865 3582 3150 3587
rect 3465 3582 3734 3587
rect 3793 3582 3822 3587
rect 553 3577 558 3582
rect 377 3572 414 3577
rect 449 3572 558 3577
rect 665 3577 670 3582
rect 3817 3577 3822 3582
rect 3905 3582 4014 3587
rect 3905 3577 3910 3582
rect 665 3572 878 3577
rect 897 3572 934 3577
rect 945 3572 982 3577
rect 1153 3572 1190 3577
rect 1217 3572 1326 3577
rect 1449 3572 1486 3577
rect 1617 3572 1734 3577
rect 1753 3572 1942 3577
rect 2065 3572 2126 3577
rect 2193 3572 2334 3577
rect 2449 3572 2718 3577
rect 2777 3572 2934 3577
rect 2953 3572 3022 3577
rect 3065 3572 3142 3577
rect 3457 3572 3526 3577
rect 3713 3572 3758 3577
rect 3817 3572 3910 3577
rect 4001 3572 4142 3577
rect 977 3567 1158 3572
rect 1617 3567 1622 3572
rect 177 3562 294 3567
rect 393 3562 846 3567
rect 889 3562 958 3567
rect 1177 3562 1342 3567
rect 1353 3562 1622 3567
rect 1729 3567 1734 3572
rect 1729 3562 1790 3567
rect 2073 3562 2134 3567
rect 2169 3562 2214 3567
rect 2273 3562 2558 3567
rect 2641 3562 2758 3567
rect 2769 3562 2894 3567
rect 2905 3562 2958 3567
rect 2969 3562 3006 3567
rect 3041 3562 3198 3567
rect 3521 3562 3558 3567
rect 4049 3562 4086 3567
rect 2769 3557 2774 3562
rect 3737 3557 3830 3562
rect 81 3552 198 3557
rect 401 3552 702 3557
rect 729 3552 910 3557
rect 1081 3552 1190 3557
rect 1233 3552 1294 3557
rect 1321 3552 1422 3557
rect 1497 3552 1534 3557
rect 1545 3552 2022 3557
rect 2065 3552 2110 3557
rect 2137 3552 2190 3557
rect 2217 3552 2262 3557
rect 2329 3552 2358 3557
rect 2425 3552 2494 3557
rect 2505 3552 2774 3557
rect 2785 3552 2886 3557
rect 2977 3552 3110 3557
rect 3177 3552 3206 3557
rect 3217 3552 3278 3557
rect 3297 3552 3438 3557
rect 3577 3552 3742 3557
rect 3825 3552 3870 3557
rect 3945 3552 3990 3557
rect 4041 3552 4118 3557
rect 2257 3547 2262 3552
rect 3297 3547 3302 3552
rect 161 3542 422 3547
rect 449 3542 582 3547
rect 889 3542 1486 3547
rect 1545 3542 1574 3547
rect 1609 3542 1654 3547
rect 1777 3542 1814 3547
rect 2033 3542 2102 3547
rect 2169 3542 2246 3547
rect 2257 3542 2494 3547
rect 577 3537 806 3542
rect 1481 3537 1550 3542
rect 2489 3537 2494 3542
rect 2585 3542 2734 3547
rect 2833 3542 3302 3547
rect 3433 3547 3438 3552
rect 3433 3542 3470 3547
rect 3489 3542 3534 3547
rect 3753 3542 3782 3547
rect 3841 3542 3878 3547
rect 3937 3542 3966 3547
rect 3977 3542 4022 3547
rect 4033 3542 4150 3547
rect 2585 3537 2590 3542
rect 2729 3537 2838 3542
rect 385 3532 462 3537
rect 513 3532 558 3537
rect 801 3532 942 3537
rect 1033 3532 1094 3537
rect 1105 3532 1222 3537
rect 1241 3532 1286 3537
rect 1393 3532 1438 3537
rect 1625 3532 1662 3537
rect 2417 3532 2438 3537
rect 2449 3532 2470 3537
rect 2489 3532 2590 3537
rect 2609 3532 2630 3537
rect 2665 3532 2710 3537
rect 2857 3532 3022 3537
rect 3033 3532 3078 3537
rect 3105 3532 3374 3537
rect 3401 3532 3422 3537
rect 3745 3532 3790 3537
rect 2417 3527 2422 3532
rect 193 3522 238 3527
rect 249 3522 366 3527
rect 425 3522 454 3527
rect 641 3522 790 3527
rect 1121 3522 1166 3527
rect 1177 3522 1238 3527
rect 1553 3522 1614 3527
rect 1673 3522 1830 3527
rect 1897 3522 1926 3527
rect 1945 3522 1966 3527
rect 2121 3522 2158 3527
rect 2417 3522 2446 3527
rect 2465 3522 2470 3532
rect 489 3517 622 3522
rect 1257 3517 1502 3522
rect 1609 3517 1678 3522
rect 2609 3517 2614 3532
rect 3953 3527 3958 3537
rect 3993 3532 4014 3537
rect 2673 3522 2774 3527
rect 2817 3522 3142 3527
rect 3217 3522 3246 3527
rect 3265 3522 3294 3527
rect 3409 3522 3494 3527
rect 3505 3522 3606 3527
rect 3769 3522 3878 3527
rect 3953 3522 3982 3527
rect 4049 3522 4094 3527
rect 2769 3517 2774 3522
rect 3137 3517 3142 3522
rect 145 3512 206 3517
rect 217 3512 262 3517
rect 273 3512 318 3517
rect 433 3512 494 3517
rect 617 3512 782 3517
rect 993 3512 1102 3517
rect 1145 3512 1190 3517
rect 1217 3512 1262 3517
rect 1497 3512 1526 3517
rect 1769 3512 1798 3517
rect 1809 3512 1862 3517
rect 1953 3512 1982 3517
rect 2009 3512 2054 3517
rect 2217 3512 2310 3517
rect 2353 3512 2382 3517
rect 2449 3512 2614 3517
rect 2625 3512 2678 3517
rect 2689 3512 2718 3517
rect 2737 3512 2758 3517
rect 2769 3512 2918 3517
rect 2937 3512 2966 3517
rect 3137 3512 3422 3517
rect 3441 3512 3574 3517
rect 3761 3512 3974 3517
rect 993 3507 998 3512
rect 2625 3507 2630 3512
rect 161 3502 414 3507
rect 505 3502 558 3507
rect 617 3502 678 3507
rect 673 3497 678 3502
rect 777 3502 998 3507
rect 1225 3502 1406 3507
rect 1417 3502 1638 3507
rect 1729 3502 1774 3507
rect 1929 3502 1982 3507
rect 2001 3502 2054 3507
rect 2321 3502 2390 3507
rect 2433 3502 2630 3507
rect 2641 3502 3038 3507
rect 3193 3502 3558 3507
rect 3569 3502 3574 3512
rect 3745 3502 3838 3507
rect 777 3497 782 3502
rect 1633 3497 1638 3502
rect 3553 3497 3558 3502
rect 3833 3497 3838 3502
rect 3897 3502 3942 3507
rect 4041 3502 4078 3507
rect 3897 3497 3902 3502
rect 225 3492 366 3497
rect 257 3482 302 3487
rect 361 3477 366 3492
rect 545 3492 606 3497
rect 673 3492 782 3497
rect 1153 3492 1614 3497
rect 1633 3492 1950 3497
rect 2249 3492 2326 3497
rect 2401 3492 2550 3497
rect 2657 3492 3046 3497
rect 3185 3492 3398 3497
rect 3417 3492 3502 3497
rect 3553 3492 3638 3497
rect 3649 3492 3814 3497
rect 3833 3492 3902 3497
rect 545 3477 550 3492
rect 2545 3487 2662 3492
rect 3393 3487 3398 3492
rect 569 3482 654 3487
rect 1017 3482 1134 3487
rect 1193 3482 1278 3487
rect 1345 3482 1382 3487
rect 1473 3482 1502 3487
rect 1993 3482 2046 3487
rect 2401 3482 2526 3487
rect 2681 3482 2862 3487
rect 2929 3482 3270 3487
rect 3393 3482 3582 3487
rect 1017 3477 1022 3482
rect 361 3472 550 3477
rect 817 3472 966 3477
rect 985 3472 1022 3477
rect 1129 3477 1134 3482
rect 1129 3472 1518 3477
rect 2281 3472 2430 3477
rect 2529 3472 2606 3477
rect 2625 3472 2662 3477
rect 2793 3472 2982 3477
rect 3025 3472 3438 3477
rect 817 3467 822 3472
rect 793 3462 822 3467
rect 961 3467 966 3472
rect 3505 3467 3622 3472
rect 961 3462 1158 3467
rect 1201 3462 1510 3467
rect 1809 3462 1870 3467
rect 2289 3462 2614 3467
rect 2721 3462 3238 3467
rect 3377 3462 3406 3467
rect 3481 3462 3510 3467
rect 3617 3462 3646 3467
rect 3233 3457 3382 3462
rect 137 3452 342 3457
rect 817 3452 974 3457
rect 1001 3452 1254 3457
rect 1273 3452 1582 3457
rect 2153 3452 2278 3457
rect 2273 3447 2278 3452
rect 2337 3452 2886 3457
rect 2913 3452 3214 3457
rect 3409 3452 3750 3457
rect 2337 3447 2342 3452
rect 297 3442 398 3447
rect 417 3442 510 3447
rect 561 3442 710 3447
rect 841 3442 878 3447
rect 961 3442 1310 3447
rect 1345 3442 1390 3447
rect 1465 3442 1486 3447
rect 2273 3442 2342 3447
rect 2361 3442 2454 3447
rect 2505 3442 2622 3447
rect 2649 3442 2822 3447
rect 2937 3442 3782 3447
rect 3833 3442 3950 3447
rect 417 3437 422 3442
rect 265 3432 302 3437
rect 329 3432 422 3437
rect 505 3437 510 3442
rect 3833 3437 3838 3442
rect 505 3432 798 3437
rect 1089 3432 1238 3437
rect 1401 3432 1574 3437
rect 1617 3432 1654 3437
rect 2393 3432 2414 3437
rect 1233 3427 1406 3432
rect 1617 3427 1622 3432
rect 2433 3427 2438 3437
rect 2489 3432 2726 3437
rect 2801 3432 3030 3437
rect 3097 3432 3190 3437
rect 3185 3427 3190 3432
rect 3473 3432 3678 3437
rect 3689 3432 3838 3437
rect 3945 3437 3950 3442
rect 3945 3432 3990 3437
rect 3473 3427 3478 3432
rect 145 3422 174 3427
rect 185 3422 230 3427
rect 385 3422 494 3427
rect 641 3422 750 3427
rect 761 3422 854 3427
rect 865 3422 918 3427
rect 1065 3422 1094 3427
rect 1185 3422 1214 3427
rect 1441 3422 1486 3427
rect 1545 3422 1622 3427
rect 1633 3422 1662 3427
rect 1681 3422 1726 3427
rect 1745 3422 1790 3427
rect 2001 3422 2038 3427
rect 2217 3422 2254 3427
rect 2313 3422 2438 3427
rect 2497 3422 2566 3427
rect 2945 3422 3094 3427
rect 3185 3422 3478 3427
rect 3497 3422 3590 3427
rect 289 3412 414 3417
rect 545 3412 598 3417
rect 737 3412 774 3417
rect 849 3407 854 3422
rect 1089 3417 1190 3422
rect 3585 3417 3590 3422
rect 3689 3422 4014 3427
rect 4033 3422 4086 3427
rect 3689 3417 3694 3422
rect 977 3412 1054 3417
rect 1265 3412 1342 3417
rect 1505 3412 1606 3417
rect 1801 3412 1894 3417
rect 2209 3412 2294 3417
rect 2305 3412 2358 3417
rect 2433 3412 2510 3417
rect 2553 3412 2726 3417
rect 2857 3412 2942 3417
rect 3001 3412 3054 3417
rect 3121 3412 3166 3417
rect 1361 3407 1486 3412
rect 3537 3407 3542 3417
rect 3585 3412 3694 3417
rect 3721 3412 3766 3417
rect 3793 3407 3798 3417
rect 4057 3412 4102 3417
rect 185 3402 270 3407
rect 297 3402 342 3407
rect 849 3402 878 3407
rect 929 3402 1142 3407
rect 1329 3402 1366 3407
rect 1481 3402 1542 3407
rect 2265 3402 2318 3407
rect 2425 3402 2846 3407
rect 2913 3402 3046 3407
rect 3209 3402 3414 3407
rect 3537 3402 3566 3407
rect 3777 3402 3798 3407
rect 3881 3402 4054 3407
rect 185 3397 190 3402
rect 161 3392 190 3397
rect 265 3397 270 3402
rect 2841 3397 2918 3402
rect 265 3392 502 3397
rect 521 3392 718 3397
rect 745 3392 830 3397
rect 1129 3392 1286 3397
rect 1393 3392 1422 3397
rect 1473 3392 1526 3397
rect 1585 3392 1702 3397
rect 1873 3392 1942 3397
rect 2369 3392 2446 3397
rect 2521 3392 2558 3397
rect 2577 3392 2670 3397
rect 2705 3392 2734 3397
rect 2937 3392 2966 3397
rect 3121 3392 3190 3397
rect 3393 3392 3422 3397
rect 3489 3392 3550 3397
rect 3585 3392 3614 3397
rect 3729 3392 3798 3397
rect 4057 3392 4078 3397
rect 745 3387 750 3392
rect 825 3387 1006 3392
rect 121 3382 182 3387
rect 233 3382 374 3387
rect 521 3382 542 3387
rect 721 3382 750 3387
rect 1001 3382 1094 3387
rect 1617 3382 1806 3387
rect 185 3372 254 3377
rect 377 3372 414 3377
rect 513 3372 990 3377
rect 1329 3372 1350 3377
rect 137 3362 182 3367
rect 217 3362 334 3367
rect 361 3362 534 3367
rect 945 3362 982 3367
rect 1233 3362 1310 3367
rect 1665 3362 1670 3382
rect 809 3357 886 3362
rect 1233 3357 1238 3362
rect 145 3352 206 3357
rect 697 3352 814 3357
rect 881 3352 910 3357
rect 953 3352 1014 3357
rect 1209 3352 1238 3357
rect 1305 3357 1310 3362
rect 1305 3352 1374 3357
rect 1553 3352 1774 3357
rect 1921 3347 1926 3392
rect 3121 3387 3126 3392
rect 3185 3387 3374 3392
rect 2305 3382 2398 3387
rect 2465 3382 2494 3387
rect 2585 3382 2742 3387
rect 2761 3382 2902 3387
rect 2921 3382 2990 3387
rect 3097 3382 3126 3387
rect 3369 3382 3574 3387
rect 3625 3382 3918 3387
rect 2489 3377 2590 3382
rect 2761 3377 2766 3382
rect 1945 3372 2022 3377
rect 2609 3372 2766 3377
rect 2897 3377 2902 3382
rect 2897 3372 3454 3377
rect 2305 3367 2414 3372
rect 3449 3367 3454 3372
rect 3577 3372 3654 3377
rect 3921 3372 3958 3377
rect 3577 3367 3582 3372
rect 3753 3367 3862 3372
rect 2241 3362 2310 3367
rect 2409 3362 2438 3367
rect 2489 3362 2646 3367
rect 2657 3362 2758 3367
rect 2809 3362 3214 3367
rect 3449 3362 3582 3367
rect 3729 3362 3758 3367
rect 3857 3362 3910 3367
rect 3993 3362 4070 3367
rect 4089 3362 4226 3367
rect 2641 3357 2646 3362
rect 3233 3357 3406 3362
rect 3905 3357 3998 3362
rect 2017 3352 2118 3357
rect 2321 3352 2526 3357
rect 2569 3352 2630 3357
rect 2641 3352 3238 3357
rect 3401 3352 3430 3357
rect 3601 3352 3646 3357
rect 3745 3352 3846 3357
rect 4041 3352 4062 3357
rect 2017 3347 2022 3352
rect 273 3342 446 3347
rect 497 3342 622 3347
rect 825 3342 918 3347
rect 1129 3342 1230 3347
rect 1265 3342 1302 3347
rect 1449 3342 1534 3347
rect 1785 3342 1830 3347
rect 1921 3342 2022 3347
rect 1449 3337 1454 3342
rect 721 3332 750 3337
rect 921 3332 966 3337
rect 1113 3332 1206 3337
rect 1217 3332 1454 3337
rect 1529 3337 1534 3342
rect 2033 3337 2038 3347
rect 2113 3342 2166 3347
rect 2209 3342 2286 3347
rect 2449 3342 2510 3347
rect 2561 3342 2806 3347
rect 2841 3342 2902 3347
rect 2921 3342 2982 3347
rect 3049 3342 3118 3347
rect 3161 3342 3230 3347
rect 3273 3342 3326 3347
rect 3369 3342 3446 3347
rect 3457 3342 3510 3347
rect 3529 3342 3566 3347
rect 3689 3342 3718 3347
rect 3753 3342 3830 3347
rect 3849 3342 3926 3347
rect 2337 3337 2430 3342
rect 2561 3337 2566 3342
rect 1529 3332 2038 3337
rect 2313 3332 2342 3337
rect 2425 3332 2566 3337
rect 2577 3332 3550 3337
rect 3721 3332 3742 3337
rect 233 3322 254 3327
rect 473 3322 550 3327
rect 601 3322 702 3327
rect 921 3322 1198 3327
rect 601 3317 606 3322
rect 129 3312 174 3317
rect 305 3312 350 3317
rect 481 3312 526 3317
rect 577 3312 606 3317
rect 697 3317 702 3322
rect 1217 3317 1222 3332
rect 2577 3327 2582 3332
rect 3569 3327 3638 3332
rect 1305 3322 1398 3327
rect 1761 3322 1782 3327
rect 2265 3322 2470 3327
rect 2521 3322 2582 3327
rect 2593 3322 2774 3327
rect 2897 3322 2926 3327
rect 2465 3317 2470 3322
rect 2921 3317 2926 3322
rect 2993 3322 3574 3327
rect 3633 3322 3734 3327
rect 3937 3322 3942 3347
rect 4025 3342 4094 3347
rect 4153 3332 4226 3337
rect 4065 3322 4110 3327
rect 2993 3317 2998 3322
rect 697 3312 766 3317
rect 785 3312 814 3317
rect 841 3312 870 3317
rect 897 3312 942 3317
rect 1113 3312 1222 3317
rect 1313 3312 1358 3317
rect 1465 3312 1534 3317
rect 1681 3312 1734 3317
rect 1769 3312 1822 3317
rect 2161 3312 2270 3317
rect 2265 3307 2270 3312
rect 2377 3312 2406 3317
rect 2465 3312 2494 3317
rect 2577 3312 2782 3317
rect 2849 3312 2878 3317
rect 2921 3312 2998 3317
rect 3097 3312 3142 3317
rect 3177 3312 3206 3317
rect 3233 3312 3454 3317
rect 3481 3312 3518 3317
rect 3529 3312 3622 3317
rect 3841 3312 3894 3317
rect 3913 3312 3990 3317
rect 4129 3312 4226 3317
rect 2377 3307 2382 3312
rect 161 3302 198 3307
rect 441 3302 774 3307
rect 801 3302 878 3307
rect 1305 3302 1366 3307
rect 1497 3302 1566 3307
rect 1713 3302 1926 3307
rect 2265 3302 2382 3307
rect 2657 3302 2806 3307
rect 3017 3302 3118 3307
rect 3425 3302 3742 3307
rect 3761 3302 4102 3307
rect 3273 3297 3406 3302
rect 457 3292 486 3297
rect 745 3292 790 3297
rect 961 3292 1094 3297
rect 1745 3292 1790 3297
rect 2193 3292 2246 3297
rect 2513 3292 2646 3297
rect 481 3287 750 3292
rect 961 3287 966 3292
rect 817 3282 966 3287
rect 1089 3287 1094 3292
rect 1809 3287 1878 3292
rect 1089 3282 1118 3287
rect 1137 3282 1286 3287
rect 1137 3277 1142 3282
rect 553 3272 718 3277
rect 737 3272 846 3277
rect 977 3272 1142 3277
rect 1281 3277 1286 3282
rect 1401 3282 1470 3287
rect 1489 3282 1534 3287
rect 1585 3282 1678 3287
rect 1777 3282 1814 3287
rect 1873 3282 2174 3287
rect 2545 3282 2606 3287
rect 1401 3277 1406 3282
rect 1281 3272 1406 3277
rect 1465 3277 1470 3282
rect 1585 3277 1590 3282
rect 1465 3272 1590 3277
rect 1673 3277 1678 3282
rect 2641 3277 2646 3292
rect 2817 3292 2918 3297
rect 3073 3292 3158 3297
rect 3249 3292 3278 3297
rect 3401 3292 3630 3297
rect 3705 3292 3750 3297
rect 4009 3292 4038 3297
rect 2817 3277 2822 3292
rect 3745 3287 3750 3292
rect 3865 3287 4014 3292
rect 3049 3282 3078 3287
rect 1673 3272 1766 3277
rect 1833 3272 1862 3277
rect 2641 3272 2822 3277
rect 3073 3277 3078 3282
rect 3169 3282 3238 3287
rect 3169 3277 3174 3282
rect 3073 3272 3174 3277
rect 3233 3277 3238 3282
rect 3297 3282 3350 3287
rect 3401 3282 3430 3287
rect 3297 3277 3302 3282
rect 3233 3272 3302 3277
rect 3425 3277 3430 3282
rect 3497 3282 3526 3287
rect 3745 3282 3870 3287
rect 3497 3277 3502 3282
rect 3425 3272 3502 3277
rect 3537 3272 3726 3277
rect 3889 3272 3982 3277
rect 4001 3272 4062 3277
rect 553 3267 558 3272
rect 281 3262 382 3267
rect 529 3262 558 3267
rect 713 3267 718 3272
rect 841 3267 982 3272
rect 1761 3267 1838 3272
rect 3889 3267 3894 3272
rect 713 3262 822 3267
rect 1097 3262 1198 3267
rect 1417 3262 1494 3267
rect 1545 3262 1662 3267
rect 2225 3262 2374 3267
rect 577 3257 694 3262
rect 1329 3257 1398 3262
rect 2225 3257 2230 3262
rect 433 3252 582 3257
rect 689 3252 1086 3257
rect 1169 3252 1334 3257
rect 1393 3252 1486 3257
rect 1681 3252 1758 3257
rect 241 3247 342 3252
rect 433 3247 438 3252
rect 1681 3247 1686 3252
rect 217 3242 246 3247
rect 337 3242 438 3247
rect 449 3242 734 3247
rect 729 3237 734 3242
rect 889 3242 918 3247
rect 1153 3242 1190 3247
rect 1345 3242 1406 3247
rect 1593 3242 1686 3247
rect 1753 3247 1758 3252
rect 1801 3252 2062 3257
rect 2185 3252 2230 3257
rect 2369 3257 2374 3262
rect 3745 3262 3846 3267
rect 3865 3262 3894 3267
rect 3977 3267 3982 3272
rect 3977 3262 4158 3267
rect 3745 3257 3750 3262
rect 2369 3252 2398 3257
rect 3257 3252 3350 3257
rect 1801 3247 1806 3252
rect 1753 3242 1806 3247
rect 2057 3247 2062 3252
rect 3257 3247 3262 3252
rect 2057 3242 2086 3247
rect 2241 3242 2782 3247
rect 3145 3242 3262 3247
rect 3345 3247 3350 3252
rect 3513 3252 3750 3257
rect 3841 3257 3846 3262
rect 3841 3252 4094 3257
rect 3513 3247 3518 3252
rect 3345 3242 3518 3247
rect 3761 3242 3830 3247
rect 3889 3242 4110 3247
rect 889 3237 894 3242
rect 1209 3237 1302 3242
rect 3825 3237 3894 3242
rect 161 3232 470 3237
rect 585 3232 678 3237
rect 729 3232 894 3237
rect 1185 3232 1214 3237
rect 1297 3232 1326 3237
rect 1361 3232 1390 3237
rect 1481 3232 1550 3237
rect 1577 3232 1742 3237
rect 1817 3232 1942 3237
rect 1961 3232 2038 3237
rect 2257 3232 2390 3237
rect 2769 3232 2790 3237
rect 3497 3232 3710 3237
rect 3745 3232 3782 3237
rect 3921 3232 4006 3237
rect 2057 3227 2134 3232
rect 129 3222 174 3227
rect 185 3222 230 3227
rect 353 3222 390 3227
rect 633 3222 678 3227
rect 689 3222 710 3227
rect 961 3222 998 3227
rect 1065 3222 1094 3227
rect 1241 3222 1286 3227
rect 1377 3222 1422 3227
rect 1529 3222 1598 3227
rect 1673 3222 1718 3227
rect 1833 3222 1878 3227
rect 1897 3222 1950 3227
rect 1969 3222 2062 3227
rect 2129 3222 2198 3227
rect 2777 3222 2838 3227
rect 2849 3222 2886 3227
rect 2937 3222 3126 3227
rect 3273 3222 3334 3227
rect 3905 3222 3950 3227
rect 689 3217 694 3222
rect 2937 3217 2942 3222
rect 273 3212 326 3217
rect 409 3212 486 3217
rect 609 3212 694 3217
rect 713 3212 830 3217
rect 969 3212 1230 3217
rect 1297 3212 1366 3217
rect 1433 3212 1542 3217
rect 1561 3212 1830 3217
rect 1921 3212 1998 3217
rect 409 3207 414 3212
rect 257 3202 414 3207
rect 481 3207 486 3212
rect 1225 3207 1302 3212
rect 1361 3207 1438 3212
rect 1825 3207 1926 3212
rect 2065 3207 2070 3217
rect 2089 3212 2118 3217
rect 2217 3212 2254 3217
rect 2785 3212 2942 3217
rect 3121 3217 3126 3222
rect 3425 3217 3662 3222
rect 3705 3217 3782 3222
rect 3121 3212 3150 3217
rect 3209 3212 3238 3217
rect 3321 3212 3430 3217
rect 3657 3212 3710 3217
rect 3777 3212 3894 3217
rect 3905 3212 3926 3217
rect 2113 3207 2118 3212
rect 3233 3207 3326 3212
rect 481 3202 510 3207
rect 777 3202 878 3207
rect 1025 3202 1158 3207
rect 1577 3202 1806 3207
rect 1953 3202 1982 3207
rect 2017 3202 2070 3207
rect 2097 3202 2118 3207
rect 2241 3202 2286 3207
rect 2633 3202 2678 3207
rect 3089 3202 3142 3207
rect 3345 3202 3374 3207
rect 161 3192 278 3197
rect 273 3187 278 3192
rect 425 3192 470 3197
rect 521 3192 542 3197
rect 665 3192 734 3197
rect 1001 3192 1590 3197
rect 1609 3192 1782 3197
rect 1793 3192 1822 3197
rect 425 3187 430 3192
rect 753 3187 918 3192
rect 1817 3187 1822 3192
rect 1937 3192 1966 3197
rect 1937 3187 1942 3192
rect 2097 3187 2102 3202
rect 3369 3197 3374 3202
rect 3441 3202 3502 3207
rect 3553 3202 3646 3207
rect 3729 3202 3766 3207
rect 3881 3202 3902 3207
rect 3441 3197 3446 3202
rect 3641 3197 3734 3202
rect 2113 3192 2134 3197
rect 2177 3192 2254 3197
rect 2465 3192 2526 3197
rect 2545 3192 2622 3197
rect 2681 3192 3046 3197
rect 3185 3192 3262 3197
rect 3369 3192 3446 3197
rect 3465 3192 3486 3197
rect 3577 3192 3622 3197
rect 3753 3192 3822 3197
rect 3865 3192 3982 3197
rect 2545 3187 2550 3192
rect 2617 3187 2686 3192
rect 185 3182 246 3187
rect 273 3182 430 3187
rect 449 3182 478 3187
rect 473 3177 478 3182
rect 553 3182 654 3187
rect 553 3177 558 3182
rect 209 3172 254 3177
rect 473 3172 558 3177
rect 649 3177 654 3182
rect 721 3182 758 3187
rect 913 3182 942 3187
rect 1057 3182 1142 3187
rect 1337 3182 1366 3187
rect 1577 3182 1606 3187
rect 1617 3182 1686 3187
rect 1817 3182 1942 3187
rect 2001 3182 2070 3187
rect 2097 3182 2118 3187
rect 2129 3182 2198 3187
rect 721 3177 726 3182
rect 1361 3177 1494 3182
rect 1577 3177 1582 3182
rect 2193 3177 2198 3182
rect 2273 3182 2550 3187
rect 2705 3182 2750 3187
rect 3217 3182 3326 3187
rect 3537 3182 3606 3187
rect 3729 3182 3926 3187
rect 2273 3177 2278 3182
rect 649 3172 726 3177
rect 745 3172 894 3177
rect 1153 3172 1238 3177
rect 1489 3172 1582 3177
rect 2033 3172 2062 3177
rect 2073 3172 2110 3177
rect 2193 3172 2278 3177
rect 2521 3172 2630 3177
rect 3017 3172 3406 3177
rect 3425 3172 3518 3177
rect 3425 3167 3430 3172
rect 3513 3167 3662 3172
rect 769 3162 982 3167
rect 1081 3162 1142 3167
rect 1201 3162 1342 3167
rect 1433 3162 1470 3167
rect 2017 3162 2070 3167
rect 2865 3162 2894 3167
rect 3161 3162 3430 3167
rect 3657 3162 3686 3167
rect 3785 3162 3894 3167
rect 1137 3157 1206 3162
rect 3785 3157 3790 3162
rect 353 3152 390 3157
rect 441 3152 582 3157
rect 601 3152 694 3157
rect 713 3152 918 3157
rect 1065 3152 1094 3157
rect 1225 3152 1470 3157
rect 1617 3152 1694 3157
rect 2097 3152 2174 3157
rect 2369 3152 2414 3157
rect 2713 3152 2790 3157
rect 3225 3152 3350 3157
rect 3401 3152 3790 3157
rect 3889 3157 3894 3162
rect 3889 3152 4070 3157
rect 353 3147 358 3152
rect 601 3147 606 3152
rect 65 3142 86 3147
rect 193 3142 358 3147
rect 377 3142 430 3147
rect 553 3142 606 3147
rect 689 3147 694 3152
rect 2713 3147 2718 3152
rect 689 3142 742 3147
rect 841 3142 886 3147
rect 945 3142 1182 3147
rect 1209 3142 1390 3147
rect 1633 3142 1654 3147
rect 1889 3142 1926 3147
rect 1993 3142 2030 3147
rect 2201 3142 2238 3147
rect 2353 3142 2382 3147
rect 2625 3142 2718 3147
rect 2785 3147 2790 3152
rect 2785 3142 3014 3147
rect 3121 3142 3254 3147
rect 65 3117 70 3142
rect 1033 3132 1110 3137
rect 1585 3132 1798 3137
rect 1841 3132 1870 3137
rect 2273 3132 2326 3137
rect 2441 3132 2582 3137
rect 2729 3132 2774 3137
rect 2785 3132 2830 3137
rect 2985 3132 3006 3137
rect 3137 3132 3166 3137
rect 1313 3127 1438 3132
rect 3161 3127 3166 3132
rect 3225 3132 3270 3137
rect 3225 3127 3230 3132
rect 81 3122 238 3127
rect 537 3122 686 3127
rect 913 3122 1318 3127
rect 1433 3122 1750 3127
rect 1745 3117 1750 3122
rect 1937 3122 1982 3127
rect 1937 3117 1942 3122
rect 65 3112 86 3117
rect 129 3112 174 3117
rect 193 3112 214 3117
rect 321 3112 358 3117
rect 401 3112 478 3117
rect 521 3112 558 3117
rect 625 3112 670 3117
rect 705 3112 742 3117
rect 777 3112 902 3117
rect 1001 3112 1062 3117
rect 1081 3112 1110 3117
rect 1329 3112 1358 3117
rect 1377 3112 1422 3117
rect 1553 3112 1582 3117
rect 1681 3112 1726 3117
rect 1745 3112 1942 3117
rect 1977 3117 1982 3122
rect 2041 3122 2446 3127
rect 3161 3122 3230 3127
rect 3265 3122 3270 3132
rect 3297 3132 3326 3137
rect 2041 3117 2046 3122
rect 1977 3112 2046 3117
rect 2209 3112 2238 3117
rect 2233 3107 2238 3112
rect 2353 3112 2382 3117
rect 2849 3112 2966 3117
rect 3009 3112 3094 3117
rect 3249 3112 3286 3117
rect 2353 3107 2358 3112
rect 225 3102 262 3107
rect 489 3102 534 3107
rect 625 3102 678 3107
rect 721 3102 774 3107
rect 993 3102 1222 3107
rect 1433 3102 1486 3107
rect 2233 3102 2358 3107
rect 2385 3102 2430 3107
rect 3185 3102 3262 3107
rect 3297 3102 3302 3132
rect 3313 3102 3318 3127
rect 3345 3102 3350 3152
rect 3497 3142 3878 3147
rect 3377 3127 3382 3137
rect 3641 3132 3702 3137
rect 3849 3132 3998 3137
rect 3377 3122 3406 3127
rect 3633 3122 3782 3127
rect 3881 3117 3966 3122
rect 3385 3112 3550 3117
rect 3737 3112 3798 3117
rect 3817 3112 3846 3117
rect 3857 3112 3886 3117
rect 3961 3112 4094 3117
rect 3905 3102 3950 3107
rect 3713 3097 3870 3102
rect 217 3092 246 3097
rect 241 3087 246 3092
rect 313 3092 614 3097
rect 689 3092 886 3097
rect 1337 3092 1830 3097
rect 3273 3092 3326 3097
rect 3593 3092 3670 3097
rect 3689 3092 3718 3097
rect 3865 3092 3894 3097
rect 313 3087 318 3092
rect 241 3082 318 3087
rect 609 3087 614 3092
rect 905 3087 1070 3092
rect 3593 3087 3598 3092
rect 609 3082 910 3087
rect 1065 3082 1342 3087
rect 1457 3082 1526 3087
rect 2937 3082 2982 3087
rect 3001 3082 3254 3087
rect 3369 3082 3550 3087
rect 3569 3082 3598 3087
rect 3665 3087 3670 3092
rect 3665 3082 3886 3087
rect 4025 3082 4142 3087
rect 3001 3077 3006 3082
rect 3249 3077 3374 3082
rect 3545 3077 3550 3082
rect 737 3072 862 3077
rect 873 3072 910 3077
rect 929 3072 1062 3077
rect 1521 3072 1606 3077
rect 1625 3072 1742 3077
rect 553 3067 718 3072
rect 1625 3067 1630 3072
rect 409 3062 558 3067
rect 713 3062 1006 3067
rect 1081 3062 1310 3067
rect 1417 3062 1494 3067
rect 1585 3062 1630 3067
rect 1737 3067 1742 3072
rect 1849 3072 2038 3077
rect 2057 3072 2086 3077
rect 2129 3072 2246 3077
rect 2969 3072 3006 3077
rect 3545 3072 3686 3077
rect 1849 3067 1854 3072
rect 1737 3062 1854 3067
rect 2033 3067 2038 3072
rect 2129 3067 2134 3072
rect 2033 3062 2134 3067
rect 2241 3067 2246 3072
rect 3681 3067 3686 3072
rect 3777 3072 3806 3077
rect 3777 3067 3782 3072
rect 2241 3062 2270 3067
rect 2761 3062 2958 3067
rect 1081 3057 1086 3062
rect 569 3052 902 3057
rect 1017 3052 1086 3057
rect 1305 3057 1310 3062
rect 2953 3057 2958 3062
rect 3017 3062 3310 3067
rect 3017 3057 3022 3062
rect 3305 3057 3310 3062
rect 3385 3062 3462 3067
rect 3385 3057 3390 3062
rect 1305 3052 1598 3057
rect 1609 3052 1726 3057
rect 1833 3052 1910 3057
rect 2089 3052 2118 3057
rect 2281 3052 2462 3057
rect 2953 3052 3022 3057
rect 3257 3052 3278 3057
rect 3305 3052 3390 3057
rect 3457 3057 3462 3062
rect 3633 3062 3662 3067
rect 3681 3062 3782 3067
rect 3633 3057 3638 3062
rect 3457 3052 3638 3057
rect 1721 3047 1838 3052
rect 2113 3047 2118 3052
rect 2217 3047 2286 3052
rect 441 3042 550 3047
rect 609 3042 662 3047
rect 777 3042 1086 3047
rect 1129 3042 1190 3047
rect 1241 3042 1294 3047
rect 1449 3042 1470 3047
rect 1593 3042 1630 3047
rect 1857 3042 2062 3047
rect 2113 3042 2222 3047
rect 2601 3042 2742 3047
rect 3089 3042 3286 3047
rect 441 3037 446 3042
rect 249 3032 446 3037
rect 545 3037 550 3042
rect 657 3037 782 3042
rect 1329 3037 1430 3042
rect 2601 3037 2606 3042
rect 545 3032 574 3037
rect 617 3032 638 3037
rect 801 3032 870 3037
rect 897 3032 1118 3037
rect 1161 3032 1262 3037
rect 1305 3032 1334 3037
rect 1425 3032 1606 3037
rect 1617 3032 1654 3037
rect 1721 3032 1774 3037
rect 1905 3032 1942 3037
rect 2241 3032 2294 3037
rect 2577 3032 2606 3037
rect 2737 3037 2742 3042
rect 3281 3037 3286 3042
rect 2737 3032 2798 3037
rect 2921 3032 3262 3037
rect 3281 3032 3438 3037
rect 3721 3032 3774 3037
rect 3793 3032 3902 3037
rect 1617 3027 1622 3032
rect 3793 3027 3798 3032
rect 233 3022 270 3027
rect 457 3022 502 3027
rect 545 3022 646 3027
rect 745 3022 814 3027
rect 857 3022 1174 3027
rect 1233 3022 1294 3027
rect 1313 3022 1374 3027
rect 1385 3022 1438 3027
rect 1561 3022 1622 3027
rect 1633 3022 1678 3027
rect 1737 3022 1862 3027
rect 1921 3022 1982 3027
rect 2257 3022 2310 3027
rect 2385 3022 2414 3027
rect 2441 3022 2518 3027
rect 2657 3022 2742 3027
rect 2785 3022 2886 3027
rect 2945 3022 2974 3027
rect 3065 3022 3102 3027
rect 3201 3022 3374 3027
rect 3465 3022 3510 3027
rect 3649 3022 3798 3027
rect 3897 3027 3902 3032
rect 3897 3022 3926 3027
rect 4025 3022 4054 3027
rect 2441 3017 2446 3022
rect 409 3012 446 3017
rect 521 3012 622 3017
rect 289 3002 358 3007
rect 657 2997 662 3017
rect 985 3012 1014 3017
rect 1025 3012 1094 3017
rect 1113 3012 1166 3017
rect 1249 3012 1310 3017
rect 1329 3012 1414 3017
rect 1577 3012 1654 3017
rect 1761 3012 1966 3017
rect 2209 3012 2350 3017
rect 2417 3012 2446 3017
rect 2513 3017 2518 3022
rect 3121 3017 3206 3022
rect 2513 3012 2542 3017
rect 2609 3012 2638 3017
rect 2745 3012 2814 3017
rect 2833 3012 2902 3017
rect 2977 3012 3126 3017
rect 3217 3012 3254 3017
rect 3265 3012 3494 3017
rect 3521 3012 3582 3017
rect 3769 3012 3862 3017
rect 4033 3012 4070 3017
rect 705 3002 790 3007
rect 841 3002 950 3007
rect 273 2992 382 2997
rect 489 2992 542 2997
rect 641 2992 750 2997
rect 761 2992 838 2997
rect 857 2992 910 2997
rect 945 2987 950 3002
rect 969 2992 990 2997
rect 1009 2987 1014 3012
rect 1161 3007 1254 3012
rect 1097 3002 1142 3007
rect 1273 3002 1326 3007
rect 1505 3002 1550 3007
rect 2209 3002 2214 3012
rect 2417 3007 2422 3012
rect 3265 3007 3270 3012
rect 2225 3002 2294 3007
rect 2305 3002 2334 3007
rect 2345 3002 2422 3007
rect 2481 3002 2718 3007
rect 2825 3002 2854 3007
rect 2953 3002 3030 3007
rect 2305 2997 2310 3002
rect 3025 2997 3030 3002
rect 3113 3002 3198 3007
rect 3217 3002 3270 3007
rect 3353 3002 3454 3007
rect 3513 3002 3638 3007
rect 3673 3002 3774 3007
rect 3113 2997 3118 3002
rect 3785 2997 3790 3007
rect 3873 3002 4022 3007
rect 4081 3002 4142 3007
rect 4017 2997 4086 3002
rect 1225 2992 1302 2997
rect 1505 2992 1934 2997
rect 2129 2992 2166 2997
rect 2177 2992 2254 2997
rect 2273 2992 2310 2997
rect 2369 2992 2518 2997
rect 2513 2987 2518 2992
rect 2601 2992 2638 2997
rect 2777 2992 2846 2997
rect 2945 2992 2998 2997
rect 3025 2992 3118 2997
rect 3177 2992 3366 2997
rect 3521 2992 3574 2997
rect 3585 2992 3718 2997
rect 3785 2992 3806 2997
rect 3905 2992 3942 2997
rect 2601 2987 2606 2992
rect 257 2982 350 2987
rect 657 2982 726 2987
rect 825 2982 894 2987
rect 945 2982 974 2987
rect 985 2982 1014 2987
rect 1081 2982 1446 2987
rect 1457 2982 1502 2987
rect 1537 2982 1590 2987
rect 1793 2982 1870 2987
rect 2081 2982 2126 2987
rect 2209 2982 2342 2987
rect 2353 2982 2430 2987
rect 2513 2982 2606 2987
rect 2625 2982 2670 2987
rect 3137 2982 3350 2987
rect 3537 2982 3598 2987
rect 3977 2982 4022 2987
rect 4065 2982 4110 2987
rect 1441 2977 1446 2982
rect 3617 2977 3734 2982
rect 441 2972 590 2977
rect 753 2972 798 2977
rect 865 2972 1014 2977
rect 1441 2972 1518 2977
rect 2081 2972 2222 2977
rect 2393 2972 2494 2977
rect 2721 2972 2902 2977
rect 3049 2972 3206 2977
rect 3273 2972 3318 2977
rect 3353 2972 3374 2977
rect 3393 2972 3478 2977
rect 3489 2972 3622 2977
rect 3729 2972 3814 2977
rect 441 2967 446 2972
rect 201 2962 254 2967
rect 273 2962 398 2967
rect 417 2962 446 2967
rect 585 2967 590 2972
rect 585 2962 614 2967
rect 729 2962 782 2967
rect 849 2962 894 2967
rect 273 2957 278 2962
rect 161 2952 278 2957
rect 393 2957 398 2962
rect 393 2952 470 2957
rect 481 2952 630 2957
rect 705 2952 862 2957
rect 145 2942 262 2947
rect 297 2942 382 2947
rect 473 2942 502 2947
rect 593 2942 646 2947
rect 377 2937 478 2942
rect 705 2937 710 2952
rect 961 2947 966 2967
rect 977 2962 1022 2967
rect 1089 2962 1126 2967
rect 1609 2962 1758 2967
rect 2193 2962 2286 2967
rect 2329 2962 2390 2967
rect 2441 2962 2486 2967
rect 2593 2962 2662 2967
rect 3113 2962 3182 2967
rect 3233 2962 3302 2967
rect 3345 2962 3878 2967
rect 1609 2957 1614 2962
rect 1281 2952 1390 2957
rect 1553 2952 1614 2957
rect 1753 2957 1758 2962
rect 1753 2952 1982 2957
rect 2009 2952 2046 2957
rect 2169 2952 2222 2957
rect 2273 2952 2374 2957
rect 2401 2952 2430 2957
rect 3097 2952 3190 2957
rect 3233 2952 3238 2962
rect 3257 2952 3294 2957
rect 3377 2952 3534 2957
rect 3625 2952 3686 2957
rect 3697 2952 3750 2957
rect 3809 2952 4038 2957
rect 3681 2947 3686 2952
rect 4033 2947 4038 2952
rect 785 2942 830 2947
rect 905 2942 1014 2947
rect 1033 2942 1174 2947
rect 1193 2942 1214 2947
rect 1273 2942 1342 2947
rect 1425 2942 1526 2947
rect 1545 2942 1742 2947
rect 1817 2942 1902 2947
rect 1993 2942 2038 2947
rect 2161 2942 2190 2947
rect 2289 2942 2350 2947
rect 2361 2942 2406 2947
rect 2521 2942 2758 2947
rect 2809 2942 2846 2947
rect 3001 2942 3086 2947
rect 3153 2942 3174 2947
rect 3225 2942 3302 2947
rect 3361 2942 3614 2947
rect 3681 2942 3710 2947
rect 3817 2942 3926 2947
rect 4033 2942 4054 2947
rect 1033 2937 1038 2942
rect 137 2932 198 2937
rect 673 2932 710 2937
rect 729 2932 1038 2937
rect 1169 2937 1174 2942
rect 1425 2937 1430 2942
rect 1169 2932 1302 2937
rect 1345 2932 1382 2937
rect 1401 2932 1430 2937
rect 1521 2937 1526 2942
rect 1521 2932 1574 2937
rect 1825 2932 1854 2937
rect 2137 2932 2166 2937
rect 193 2927 198 2932
rect 1057 2927 1150 2932
rect 193 2922 222 2927
rect 337 2922 454 2927
rect 545 2922 606 2927
rect 633 2922 1062 2927
rect 1145 2922 1526 2927
rect 1537 2922 1582 2927
rect 1609 2922 1654 2927
rect 545 2917 550 2922
rect 1825 2917 1830 2932
rect 2161 2927 2166 2932
rect 2249 2932 2310 2937
rect 2417 2932 2446 2937
rect 2249 2927 2254 2932
rect 2481 2927 2694 2932
rect 2753 2927 2758 2942
rect 3705 2937 3822 2942
rect 2825 2932 2870 2937
rect 3049 2932 3070 2937
rect 3105 2932 3174 2937
rect 3193 2927 3286 2932
rect 1857 2922 1878 2927
rect 2161 2922 2254 2927
rect 2313 2922 2374 2927
rect 2385 2922 2414 2927
rect 2457 2922 2486 2927
rect 2689 2922 2718 2927
rect 2753 2922 2814 2927
rect 2873 2922 2926 2927
rect 3017 2922 3198 2927
rect 3281 2922 3310 2927
rect 3337 2922 3366 2927
rect 145 2912 174 2917
rect 361 2912 406 2917
rect 497 2912 550 2917
rect 601 2912 654 2917
rect 689 2912 766 2917
rect 881 2912 958 2917
rect 993 2912 1086 2917
rect 1137 2912 1294 2917
rect 1313 2912 1334 2917
rect 1377 2912 1422 2917
rect 1513 2912 1622 2917
rect 1633 2912 1678 2917
rect 1697 2912 1806 2917
rect 1825 2912 1862 2917
rect 1881 2912 1926 2917
rect 1945 2912 2070 2917
rect 2273 2912 2334 2917
rect 2385 2912 2390 2922
rect 3441 2917 3446 2937
rect 3657 2932 3678 2937
rect 3905 2932 4046 2937
rect 4073 2932 4142 2937
rect 3529 2922 3830 2927
rect 3841 2922 3894 2927
rect 3825 2917 3830 2922
rect 2497 2912 2838 2917
rect 3049 2912 3102 2917
rect 3193 2912 3254 2917
rect 3281 2912 3382 2917
rect 3401 2912 3422 2917
rect 3441 2912 3470 2917
rect 3505 2912 3558 2917
rect 3633 2912 3654 2917
rect 3785 2912 3806 2917
rect 3825 2912 3854 2917
rect 1617 2907 1622 2912
rect 1697 2907 1702 2912
rect 457 2902 510 2907
rect 721 2902 830 2907
rect 937 2902 998 2907
rect 1081 2902 1254 2907
rect 1321 2902 1550 2907
rect 1617 2902 1702 2907
rect 1801 2907 1806 2912
rect 3281 2907 3286 2912
rect 3849 2907 3854 2912
rect 3945 2912 4030 2917
rect 3945 2907 3950 2912
rect 1801 2902 1934 2907
rect 2289 2902 2374 2907
rect 2393 2902 2422 2907
rect 2417 2897 2422 2902
rect 2545 2902 2574 2907
rect 2689 2902 2766 2907
rect 2937 2902 3038 2907
rect 3121 2902 3286 2907
rect 3465 2902 3510 2907
rect 2545 2897 2550 2902
rect 3505 2897 3510 2902
rect 3569 2902 3782 2907
rect 3793 2902 3830 2907
rect 3849 2902 3950 2907
rect 3569 2897 3574 2902
rect 3777 2897 3782 2902
rect 601 2892 702 2897
rect 873 2892 1566 2897
rect 1577 2892 1606 2897
rect 1689 2892 2118 2897
rect 2233 2892 2342 2897
rect 2417 2892 2550 2897
rect 2865 2892 2926 2897
rect 3169 2892 3486 2897
rect 3505 2892 3574 2897
rect 3617 2892 3718 2897
rect 3777 2892 3798 2897
rect 601 2887 606 2892
rect 441 2882 526 2887
rect 553 2882 606 2887
rect 697 2887 702 2892
rect 1601 2887 1694 2892
rect 2921 2887 2926 2892
rect 3057 2887 3174 2892
rect 697 2882 806 2887
rect 905 2882 974 2887
rect 1089 2882 1150 2887
rect 1177 2882 1230 2887
rect 1257 2882 1574 2887
rect 1713 2882 1982 2887
rect 1977 2877 1982 2882
rect 2073 2882 2102 2887
rect 2121 2882 2158 2887
rect 2209 2882 2246 2887
rect 2921 2882 3062 2887
rect 3193 2882 3222 2887
rect 2073 2877 2078 2882
rect 3481 2877 3486 2892
rect 3617 2877 3622 2892
rect 209 2872 294 2877
rect 617 2872 686 2877
rect 777 2872 958 2877
rect 1033 2872 1278 2877
rect 1305 2872 1446 2877
rect 1497 2872 1702 2877
rect 1745 2872 1958 2877
rect 1977 2872 2078 2877
rect 3081 2872 3206 2877
rect 3481 2872 3622 2877
rect 209 2867 214 2872
rect 185 2862 214 2867
rect 289 2867 294 2872
rect 681 2867 782 2872
rect 289 2862 558 2867
rect 609 2862 646 2867
rect 801 2862 1110 2867
rect 1161 2862 1190 2867
rect 1273 2862 1302 2867
rect 1337 2862 1366 2867
rect 1537 2862 1838 2867
rect 1857 2862 1886 2867
rect 3249 2862 3438 2867
rect 1185 2857 1278 2862
rect 1361 2857 1542 2862
rect 3065 2857 3142 2862
rect 3249 2857 3254 2862
rect 217 2852 334 2857
rect 585 2852 630 2857
rect 761 2852 1038 2857
rect 1057 2852 1166 2857
rect 1561 2852 1734 2857
rect 2569 2852 2686 2857
rect 3041 2852 3070 2857
rect 3137 2852 3254 2857
rect 3433 2857 3438 2862
rect 3761 2862 3918 2867
rect 3433 2852 3462 2857
rect 3641 2852 3718 2857
rect 3641 2847 3646 2852
rect 489 2842 854 2847
rect 961 2842 1046 2847
rect 1129 2842 1270 2847
rect 1417 2842 1494 2847
rect 1545 2842 1630 2847
rect 2969 2842 3022 2847
rect 3033 2842 3126 2847
rect 3305 2842 3646 2847
rect 3713 2847 3718 2852
rect 3761 2847 3766 2862
rect 3913 2847 3918 2862
rect 3937 2852 4030 2857
rect 3713 2842 3766 2847
rect 3793 2842 3862 2847
rect 3913 2842 4070 2847
rect 1041 2837 1134 2842
rect 3793 2837 3798 2842
rect 313 2832 430 2837
rect 513 2832 550 2837
rect 569 2832 654 2837
rect 729 2832 854 2837
rect 945 2832 1022 2837
rect 1153 2832 1198 2837
rect 1209 2832 1254 2837
rect 1305 2832 1398 2837
rect 1577 2832 1638 2837
rect 1665 2832 1806 2837
rect 1937 2832 2038 2837
rect 2345 2832 2390 2837
rect 2505 2832 2574 2837
rect 1305 2827 1310 2832
rect 129 2822 174 2827
rect 281 2822 326 2827
rect 353 2807 358 2827
rect 369 2822 614 2827
rect 625 2822 662 2827
rect 673 2822 766 2827
rect 833 2822 870 2827
rect 1025 2822 1078 2827
rect 609 2817 614 2822
rect 673 2817 678 2822
rect 889 2817 990 2822
rect 1089 2817 1094 2827
rect 1121 2822 1174 2827
rect 1193 2822 1238 2827
rect 1281 2822 1310 2827
rect 1393 2827 1398 2832
rect 2569 2827 2574 2832
rect 2649 2832 2774 2837
rect 3025 2832 3070 2837
rect 3265 2832 3294 2837
rect 2649 2827 2654 2832
rect 1393 2822 1566 2827
rect 1585 2822 1614 2827
rect 1737 2822 1782 2827
rect 1793 2822 1870 2827
rect 2057 2822 2134 2827
rect 2217 2822 2310 2827
rect 2401 2822 2438 2827
rect 2449 2822 2550 2827
rect 2569 2822 2654 2827
rect 2953 2822 2998 2827
rect 3225 2822 3246 2827
rect 609 2812 678 2817
rect 753 2812 790 2817
rect 857 2812 894 2817
rect 985 2812 1014 2817
rect 1089 2812 1134 2817
rect 1281 2812 1302 2817
rect 1321 2812 1398 2817
rect 1521 2812 1606 2817
rect 473 2807 590 2812
rect 1153 2807 1262 2812
rect 1649 2807 1654 2817
rect 1761 2812 1822 2817
rect 1857 2812 1878 2817
rect 1969 2812 2222 2817
rect 2401 2812 2422 2817
rect 169 2802 206 2807
rect 321 2802 358 2807
rect 449 2802 478 2807
rect 585 2802 814 2807
rect 833 2802 966 2807
rect 1025 2802 1158 2807
rect 1257 2802 1566 2807
rect 1593 2802 1654 2807
rect 2289 2802 2398 2807
rect 2433 2802 2438 2822
rect 3017 2812 3054 2817
rect 3081 2812 3126 2817
rect 3265 2812 3270 2832
rect 3313 2817 3318 2837
rect 3345 2832 3390 2837
rect 3433 2832 3470 2837
rect 3665 2832 3798 2837
rect 3857 2837 3862 2842
rect 3857 2832 3974 2837
rect 3985 2832 4014 2837
rect 4057 2832 4094 2837
rect 3353 2822 3382 2827
rect 3393 2822 3478 2827
rect 3505 2822 3566 2827
rect 3601 2822 3678 2827
rect 3809 2822 3846 2827
rect 3921 2822 3958 2827
rect 4001 2822 4078 2827
rect 3313 2812 3358 2817
rect 3369 2812 3398 2817
rect 3481 2812 3598 2817
rect 3961 2812 4014 2817
rect 2889 2802 2974 2807
rect 3009 2802 3038 2807
rect 961 2797 1030 2802
rect 1953 2797 2102 2802
rect 3033 2797 3038 2802
rect 3129 2802 3254 2807
rect 3129 2797 3134 2802
rect 3249 2797 3254 2802
rect 3409 2802 3630 2807
rect 3409 2797 3414 2802
rect 161 2792 478 2797
rect 505 2792 590 2797
rect 601 2792 670 2797
rect 857 2792 942 2797
rect 1137 2792 1206 2797
rect 1241 2792 1270 2797
rect 1321 2792 1502 2797
rect 1585 2792 1622 2797
rect 1641 2792 1686 2797
rect 1737 2792 1838 2797
rect 1929 2792 1958 2797
rect 2097 2792 2150 2797
rect 2217 2792 2278 2797
rect 2449 2792 2798 2797
rect 2833 2792 2854 2797
rect 2905 2792 2990 2797
rect 3033 2792 3134 2797
rect 3153 2792 3230 2797
rect 3249 2792 3414 2797
rect 3537 2792 3582 2797
rect 3753 2792 3782 2797
rect 4041 2792 4222 2797
rect 705 2787 838 2792
rect 2273 2787 2454 2792
rect 81 2782 238 2787
rect 257 2782 542 2787
rect 561 2782 614 2787
rect 681 2782 710 2787
rect 833 2782 918 2787
rect 961 2782 1054 2787
rect 1073 2782 1398 2787
rect 1497 2782 1670 2787
rect 1689 2782 1774 2787
rect 1833 2782 2206 2787
rect 3529 2782 3606 2787
rect 3665 2782 3766 2787
rect 961 2777 966 2782
rect 225 2772 278 2777
rect 289 2772 422 2777
rect 433 2772 694 2777
rect 745 2772 830 2777
rect 921 2772 966 2777
rect 1049 2777 1054 2782
rect 1393 2777 1478 2782
rect 1049 2772 1078 2777
rect 1089 2772 1302 2777
rect 1313 2772 1374 2777
rect 1473 2772 2358 2777
rect 2377 2772 2494 2777
rect 3369 2772 3542 2777
rect 3649 2772 3678 2777
rect 4009 2772 4102 2777
rect 825 2767 926 2772
rect 1089 2767 1094 2772
rect 2377 2767 2382 2772
rect 265 2762 374 2767
rect 401 2762 806 2767
rect 945 2762 1094 2767
rect 1137 2762 1318 2767
rect 1329 2762 1414 2767
rect 1433 2762 1750 2767
rect 1793 2762 1934 2767
rect 2073 2762 2142 2767
rect 2249 2762 2382 2767
rect 2489 2767 2494 2772
rect 3537 2767 3654 2772
rect 2489 2762 2758 2767
rect 3329 2762 3350 2767
rect 3489 2762 3518 2767
rect 3785 2762 3894 2767
rect 193 2752 262 2757
rect 329 2752 422 2757
rect 441 2752 950 2757
rect 1129 2752 1174 2757
rect 1249 2752 1278 2757
rect 1289 2752 1342 2757
rect 1377 2752 1462 2757
rect 1553 2752 1606 2757
rect 1625 2752 1686 2757
rect 1745 2747 1750 2762
rect 1953 2757 2046 2762
rect 3785 2757 3790 2762
rect 1825 2752 1958 2757
rect 2041 2752 2070 2757
rect 2081 2752 2478 2757
rect 2689 2752 2750 2757
rect 3185 2752 3214 2757
rect 3233 2752 3310 2757
rect 3641 2752 3790 2757
rect 3889 2757 3894 2762
rect 3889 2752 3918 2757
rect 4017 2752 4054 2757
rect 241 2742 390 2747
rect 473 2742 526 2747
rect 641 2742 862 2747
rect 961 2742 982 2747
rect 1025 2742 1238 2747
rect 1305 2742 1654 2747
rect 1665 2742 1726 2747
rect 1745 2742 1950 2747
rect 1985 2742 2174 2747
rect 2193 2742 2230 2747
rect 2337 2742 2486 2747
rect 2633 2742 2670 2747
rect 3273 2742 3486 2747
rect 3609 2742 3662 2747
rect 3809 2742 3910 2747
rect 1233 2737 1310 2742
rect 2481 2737 2486 2742
rect 161 2732 206 2737
rect 281 2732 310 2737
rect 377 2732 414 2737
rect 793 2732 1038 2737
rect 1057 2732 1142 2737
rect 1329 2732 1366 2737
rect 1393 2732 1422 2737
rect 1057 2727 1062 2732
rect 1417 2727 1422 2732
rect 1553 2732 1902 2737
rect 2481 2732 2694 2737
rect 2801 2732 2870 2737
rect 3161 2732 3254 2737
rect 1553 2727 1558 2732
rect 2017 2727 2414 2732
rect 3161 2727 3166 2732
rect 297 2722 342 2727
rect 353 2722 462 2727
rect 705 2722 862 2727
rect 1025 2722 1062 2727
rect 1073 2722 1286 2727
rect 1297 2722 1342 2727
rect 1417 2722 1558 2727
rect 1577 2722 1814 2727
rect 1025 2717 1030 2722
rect 177 2712 254 2717
rect 273 2712 294 2717
rect 321 2712 382 2717
rect 393 2712 438 2717
rect 521 2712 566 2717
rect 689 2712 734 2717
rect 793 2712 1030 2717
rect 1049 2712 1398 2717
rect 1633 2712 1686 2717
rect 1697 2712 1798 2717
rect 1809 2712 1814 2722
rect 1793 2707 1798 2712
rect 265 2702 334 2707
rect 417 2702 454 2707
rect 553 2702 710 2707
rect 721 2702 774 2707
rect 1033 2702 1334 2707
rect 1345 2702 1390 2707
rect 1465 2702 1670 2707
rect 1793 2702 1886 2707
rect 1937 2702 1942 2727
rect 1993 2722 2022 2727
rect 2409 2722 2438 2727
rect 2913 2722 2966 2727
rect 3113 2722 3166 2727
rect 3249 2727 3254 2732
rect 3249 2722 3374 2727
rect 2433 2717 2438 2722
rect 2001 2712 2070 2717
rect 2097 2712 2334 2717
rect 2369 2712 2422 2717
rect 2433 2712 2534 2717
rect 2609 2712 2774 2717
rect 2817 2712 2886 2717
rect 2969 2712 3086 2717
rect 3177 2712 3238 2717
rect 3393 2707 3398 2737
rect 3689 2732 3790 2737
rect 3801 2732 3862 2737
rect 3945 2732 3998 2737
rect 3665 2722 3926 2727
rect 3457 2712 3518 2717
rect 3641 2712 4046 2717
rect 1961 2702 2254 2707
rect 2345 2702 2390 2707
rect 2425 2702 2550 2707
rect 2865 2702 2934 2707
rect 2985 2702 3126 2707
rect 3201 2702 3278 2707
rect 3345 2702 3414 2707
rect 3489 2702 3526 2707
rect 3681 2702 3926 2707
rect 705 2697 710 2702
rect 2569 2697 2718 2702
rect 3921 2697 3926 2702
rect 3993 2702 4150 2707
rect 3993 2697 3998 2702
rect 185 2692 270 2697
rect 265 2687 270 2692
rect 329 2692 358 2697
rect 593 2692 614 2697
rect 705 2692 790 2697
rect 833 2692 934 2697
rect 953 2692 1438 2697
rect 1761 2692 1926 2697
rect 2041 2692 2318 2697
rect 2337 2692 2574 2697
rect 2713 2692 3102 2697
rect 3209 2692 3262 2697
rect 3505 2692 3542 2697
rect 3921 2692 3998 2697
rect 329 2687 334 2692
rect 833 2687 838 2692
rect 153 2682 246 2687
rect 265 2682 334 2687
rect 553 2682 798 2687
rect 809 2682 838 2687
rect 929 2687 934 2692
rect 1937 2687 2046 2692
rect 3681 2687 3750 2692
rect 929 2682 1486 2687
rect 1505 2682 1590 2687
rect 1609 2682 1726 2687
rect 1785 2682 1814 2687
rect 1609 2677 1614 2682
rect 377 2672 486 2677
rect 505 2672 630 2677
rect 713 2672 774 2677
rect 809 2672 830 2677
rect 873 2672 926 2677
rect 1017 2672 1206 2677
rect 1257 2672 1286 2677
rect 1393 2672 1614 2677
rect 1721 2677 1726 2682
rect 1809 2677 1814 2682
rect 1937 2677 1942 2687
rect 2065 2682 2702 2687
rect 2865 2682 3030 2687
rect 2697 2677 2870 2682
rect 1721 2672 1750 2677
rect 1809 2672 1942 2677
rect 2017 2672 2102 2677
rect 2113 2672 2190 2677
rect 2241 2672 2270 2677
rect 2385 2672 2438 2677
rect 2481 2672 2678 2677
rect 2889 2672 2950 2677
rect 377 2667 382 2672
rect 209 2662 382 2667
rect 481 2667 486 2672
rect 1281 2667 1398 2672
rect 3025 2667 3030 2682
rect 3265 2682 3334 2687
rect 3265 2667 3270 2682
rect 3329 2677 3334 2682
rect 3425 2682 3686 2687
rect 3745 2682 3774 2687
rect 3425 2677 3430 2682
rect 3329 2672 3430 2677
rect 3497 2672 3526 2677
rect 481 2662 510 2667
rect 537 2662 870 2667
rect 945 2662 1246 2667
rect 1417 2662 1766 2667
rect 2033 2662 2206 2667
rect 2489 2662 2662 2667
rect 2753 2662 3006 2667
rect 3025 2662 3270 2667
rect 3521 2657 3526 2672
rect 3697 2672 3726 2677
rect 3697 2657 3702 2672
rect 633 2652 758 2657
rect 833 2652 974 2657
rect 1081 2652 1110 2657
rect 1137 2652 1158 2657
rect 1289 2652 1318 2657
rect 1401 2652 1782 2657
rect 1873 2652 1998 2657
rect 2105 2652 2182 2657
rect 2537 2652 2566 2657
rect 2561 2647 2566 2652
rect 2657 2652 2742 2657
rect 2953 2652 2990 2657
rect 3521 2652 3702 2657
rect 2657 2647 2662 2652
rect 2865 2647 2934 2652
rect 353 2642 558 2647
rect 673 2642 702 2647
rect 769 2642 854 2647
rect 921 2642 1014 2647
rect 1025 2642 1078 2647
rect 1161 2642 1214 2647
rect 1433 2642 1478 2647
rect 1521 2642 1638 2647
rect 1689 2642 1846 2647
rect 1857 2642 1990 2647
rect 2001 2642 2086 2647
rect 2097 2642 2158 2647
rect 2561 2642 2662 2647
rect 2681 2642 2758 2647
rect 2793 2642 2870 2647
rect 2929 2642 2974 2647
rect 3289 2642 3310 2647
rect 4001 2642 4102 2647
rect 697 2637 774 2642
rect 1233 2637 1414 2642
rect 81 2632 110 2637
rect 369 2632 422 2637
rect 825 2632 1238 2637
rect 1409 2632 1518 2637
rect 1753 2632 1790 2637
rect 1865 2632 1958 2637
rect 1993 2632 2022 2637
rect 2153 2632 2278 2637
rect 2721 2632 2782 2637
rect 2881 2632 3046 2637
rect 81 2607 86 2632
rect 1537 2627 1734 2632
rect 113 2617 118 2627
rect 153 2622 206 2627
rect 313 2622 350 2627
rect 401 2622 446 2627
rect 545 2622 614 2627
rect 649 2622 718 2627
rect 777 2622 1542 2627
rect 1729 2622 1782 2627
rect 1897 2622 2038 2627
rect 2089 2622 2166 2627
rect 2209 2622 2262 2627
rect 2353 2622 2398 2627
rect 2473 2622 2558 2627
rect 2617 2622 2670 2627
rect 2729 2622 2798 2627
rect 2833 2622 2862 2627
rect 2905 2622 2998 2627
rect 3121 2622 3158 2627
rect 3313 2617 3318 2637
rect 3401 2622 3430 2627
rect 113 2612 206 2617
rect 377 2612 542 2617
rect 577 2612 662 2617
rect 817 2612 846 2617
rect 865 2612 886 2617
rect 897 2612 942 2617
rect 969 2612 1046 2617
rect 1057 2612 1198 2617
rect 1313 2612 1582 2617
rect 1593 2612 1806 2617
rect 1953 2612 2726 2617
rect 2761 2612 2878 2617
rect 81 2602 110 2607
rect 145 2602 238 2607
rect 345 2602 622 2607
rect 817 2597 822 2612
rect 849 2602 870 2607
rect 113 2592 174 2597
rect 265 2592 422 2597
rect 521 2592 726 2597
rect 817 2592 846 2597
rect 529 2582 558 2587
rect 553 2577 558 2582
rect 673 2582 838 2587
rect 881 2582 886 2612
rect 1041 2607 1046 2612
rect 1193 2607 1318 2612
rect 1825 2607 1934 2612
rect 945 2602 990 2607
rect 1001 2602 1022 2607
rect 1041 2602 1110 2607
rect 1121 2602 1174 2607
rect 1337 2602 1830 2607
rect 1929 2602 2366 2607
rect 2737 2602 2838 2607
rect 2537 2597 2718 2602
rect 969 2592 1054 2597
rect 1137 2592 1158 2597
rect 1225 2592 1446 2597
rect 1457 2592 1598 2597
rect 1657 2592 1958 2597
rect 1969 2592 2030 2597
rect 2049 2592 2542 2597
rect 2713 2592 2766 2597
rect 2801 2592 2886 2597
rect 1457 2587 1462 2592
rect 985 2582 1046 2587
rect 1057 2582 1406 2587
rect 1433 2582 1462 2587
rect 1545 2582 1814 2587
rect 1825 2582 2062 2587
rect 2145 2582 2238 2587
rect 2337 2582 2390 2587
rect 2553 2582 2758 2587
rect 2801 2582 2894 2587
rect 2913 2582 2918 2617
rect 3177 2612 3246 2617
rect 3313 2612 3398 2617
rect 3177 2607 3182 2612
rect 3137 2602 3182 2607
rect 3241 2607 3246 2612
rect 3241 2602 3270 2607
rect 2929 2592 2958 2597
rect 2969 2592 3102 2597
rect 3217 2592 3246 2597
rect 3289 2592 3326 2597
rect 3097 2587 3222 2592
rect 2953 2582 3062 2587
rect 3345 2582 3454 2587
rect 3473 2582 3478 2637
rect 3873 2632 3894 2637
rect 3953 2632 4030 2637
rect 3529 2622 3566 2627
rect 3681 2622 3814 2627
rect 3873 2607 3878 2632
rect 3905 2622 3934 2627
rect 3897 2612 3918 2617
rect 4097 2612 4102 2642
rect 3769 2602 3790 2607
rect 3873 2602 4030 2607
rect 3497 2592 3702 2597
rect 3785 2592 3966 2597
rect 3793 2582 3862 2587
rect 673 2577 678 2582
rect 881 2577 966 2582
rect 1057 2577 1062 2582
rect 1809 2577 1814 2582
rect 2409 2577 2534 2582
rect 3345 2577 3350 2582
rect 553 2572 678 2577
rect 753 2572 782 2577
rect 809 2572 870 2577
rect 961 2572 1014 2577
rect 1041 2572 1062 2577
rect 1089 2572 1206 2577
rect 1217 2572 1254 2577
rect 1313 2572 1470 2577
rect 1729 2572 1766 2577
rect 1809 2572 1902 2577
rect 1985 2572 2062 2577
rect 2113 2572 2246 2577
rect 2289 2572 2414 2577
rect 2529 2572 2990 2577
rect 2289 2567 2294 2572
rect 2985 2567 2990 2572
rect 3073 2572 3350 2577
rect 3449 2577 3454 2582
rect 3449 2572 3710 2577
rect 3073 2567 3078 2572
rect 65 2562 142 2567
rect 833 2562 878 2567
rect 921 2562 1030 2567
rect 1105 2562 1422 2567
rect 1465 2562 1686 2567
rect 2057 2562 2294 2567
rect 2305 2562 2710 2567
rect 2769 2562 2798 2567
rect 2809 2562 2966 2567
rect 2985 2562 3078 2567
rect 3377 2562 3502 2567
rect 3513 2562 3646 2567
rect 1681 2557 1958 2562
rect 3377 2557 3382 2562
rect 481 2552 606 2557
rect 713 2552 790 2557
rect 809 2552 1238 2557
rect 1337 2552 1374 2557
rect 1953 2552 1982 2557
rect 2041 2552 2094 2557
rect 2121 2552 2654 2557
rect 2673 2552 2702 2557
rect 2785 2552 2814 2557
rect 2881 2552 2958 2557
rect 3161 2552 3190 2557
rect 3241 2552 3382 2557
rect 3393 2552 3438 2557
rect 4113 2552 4150 2557
rect 785 2547 790 2552
rect 2697 2547 2790 2552
rect 3393 2547 3398 2552
rect 3457 2547 3574 2552
rect 81 2542 206 2547
rect 593 2542 670 2547
rect 785 2542 878 2547
rect 897 2542 982 2547
rect 993 2542 1366 2547
rect 1377 2542 1406 2547
rect 1497 2542 1574 2547
rect 1593 2542 1710 2547
rect 1721 2542 1878 2547
rect 1897 2542 2030 2547
rect 2201 2542 2230 2547
rect 2241 2542 2398 2547
rect 2409 2542 2534 2547
rect 2593 2542 2678 2547
rect 2865 2542 2950 2547
rect 3081 2542 3134 2547
rect 3297 2542 3398 2547
rect 3409 2542 3462 2547
rect 3569 2542 3726 2547
rect 993 2537 998 2542
rect 1377 2537 1382 2542
rect 1497 2537 1502 2542
rect 225 2532 462 2537
rect 673 2532 718 2537
rect 921 2532 998 2537
rect 1009 2532 1094 2537
rect 1137 2532 1206 2537
rect 1353 2532 1382 2537
rect 1441 2532 1502 2537
rect 1569 2537 1574 2542
rect 2241 2537 2246 2542
rect 1569 2532 1718 2537
rect 1753 2532 1814 2537
rect 2057 2532 2150 2537
rect 2169 2532 2246 2537
rect 2257 2532 2318 2537
rect 2337 2532 2382 2537
rect 105 2522 206 2527
rect 225 2517 230 2532
rect 129 2512 230 2517
rect 457 2517 462 2532
rect 737 2527 902 2532
rect 1225 2527 1294 2532
rect 2057 2527 2062 2532
rect 601 2522 638 2527
rect 705 2522 742 2527
rect 897 2522 1046 2527
rect 1057 2522 1230 2527
rect 1289 2522 2062 2527
rect 2145 2527 2150 2532
rect 2433 2527 2438 2542
rect 3153 2537 3302 2542
rect 2449 2532 2494 2537
rect 2785 2532 3158 2537
rect 3321 2532 3398 2537
rect 3425 2532 3558 2537
rect 3737 2532 3894 2537
rect 2657 2527 2758 2532
rect 2145 2522 2438 2527
rect 2593 2522 2614 2527
rect 2633 2522 2662 2527
rect 2753 2522 2782 2527
rect 2825 2522 2934 2527
rect 3025 2522 3118 2527
rect 3129 2522 3998 2527
rect 457 2512 646 2517
rect 689 2512 926 2517
rect 945 2512 990 2517
rect 1049 2512 1118 2517
rect 1201 2512 1278 2517
rect 1409 2512 1454 2517
rect 1561 2512 1622 2517
rect 1689 2512 1766 2517
rect 1809 2512 1854 2517
rect 2073 2512 2158 2517
rect 2233 2512 2302 2517
rect 2385 2512 2606 2517
rect 2641 2512 2670 2517
rect 2689 2512 2734 2517
rect 3001 2512 3070 2517
rect 3113 2512 3158 2517
rect 3241 2512 3270 2517
rect 3393 2512 3422 2517
rect 3489 2512 3566 2517
rect 3705 2512 3750 2517
rect 3833 2512 3886 2517
rect 3937 2512 3966 2517
rect 4009 2512 4062 2517
rect 1297 2507 1390 2512
rect 185 2502 502 2507
rect 713 2502 830 2507
rect 873 2502 1062 2507
rect 1113 2502 1190 2507
rect 1265 2502 1302 2507
rect 1385 2502 1806 2507
rect 1865 2502 2574 2507
rect 2649 2502 2678 2507
rect 2873 2502 2910 2507
rect 2985 2502 3046 2507
rect 3161 2502 3830 2507
rect 1185 2497 1270 2502
rect 1801 2497 1870 2502
rect 737 2492 774 2497
rect 993 2492 1150 2497
rect 1289 2492 1310 2497
rect 1361 2492 1414 2497
rect 1753 2492 1782 2497
rect 2049 2492 2094 2497
rect 2105 2492 2142 2497
rect 2153 2492 2190 2497
rect 2329 2492 2382 2497
rect 2417 2492 2446 2497
rect 2569 2492 2662 2497
rect 2793 2492 2902 2497
rect 2953 2492 3022 2497
rect 3153 2492 3390 2497
rect 3689 2492 3766 2497
rect 3873 2492 3950 2497
rect 1625 2487 1734 2492
rect 1929 2487 2030 2492
rect 2209 2487 2310 2492
rect 3041 2487 3134 2492
rect 3873 2487 3878 2492
rect 273 2482 646 2487
rect 849 2482 1278 2487
rect 1425 2482 1630 2487
rect 1729 2482 1934 2487
rect 2025 2482 2214 2487
rect 2305 2482 2782 2487
rect 2857 2482 2886 2487
rect 2945 2482 3046 2487
rect 3129 2482 3174 2487
rect 3249 2482 3326 2487
rect 3385 2482 3878 2487
rect 3945 2487 3950 2492
rect 3945 2482 3974 2487
rect 273 2477 278 2482
rect 249 2472 278 2477
rect 641 2477 646 2482
rect 1273 2477 1430 2482
rect 2777 2477 2862 2482
rect 641 2472 670 2477
rect 697 2472 830 2477
rect 977 2472 1078 2477
rect 1089 2472 1110 2477
rect 1641 2472 1710 2477
rect 1737 2472 1782 2477
rect 1945 2472 1990 2477
rect 2001 2472 2390 2477
rect 2665 2472 2702 2477
rect 3017 2472 3166 2477
rect 3329 2472 3414 2477
rect 3817 2472 4030 2477
rect 305 2467 438 2472
rect 697 2467 702 2472
rect 825 2467 958 2472
rect 1129 2467 1238 2472
rect 2409 2467 2630 2472
rect 121 2462 214 2467
rect 289 2462 310 2467
rect 433 2462 662 2467
rect 673 2462 702 2467
rect 953 2462 1134 2467
rect 1233 2462 1438 2467
rect 1505 2462 1582 2467
rect 1681 2462 1942 2467
rect 1953 2462 2414 2467
rect 2625 2462 2654 2467
rect 209 2457 294 2462
rect 1937 2457 1942 2462
rect 2649 2457 2654 2462
rect 2713 2462 2854 2467
rect 3097 2462 3934 2467
rect 2713 2457 2718 2462
rect 3929 2457 3934 2462
rect 4017 2462 4046 2467
rect 4017 2457 4022 2462
rect 321 2452 1222 2457
rect 1473 2452 1630 2457
rect 1713 2452 1774 2457
rect 1937 2452 2006 2457
rect 2025 2452 2310 2457
rect 2425 2452 2462 2457
rect 2513 2452 2630 2457
rect 2649 2452 2718 2457
rect 2897 2452 2998 2457
rect 3041 2452 3662 2457
rect 3785 2452 3814 2457
rect 3929 2452 4022 2457
rect 1793 2447 1918 2452
rect 2897 2447 2902 2452
rect 169 2442 582 2447
rect 593 2442 622 2447
rect 649 2442 758 2447
rect 945 2442 1118 2447
rect 1241 2442 1358 2447
rect 1401 2442 1798 2447
rect 1913 2442 1942 2447
rect 1969 2442 2014 2447
rect 2137 2442 2166 2447
rect 2177 2442 2294 2447
rect 2465 2442 2542 2447
rect 2761 2442 2902 2447
rect 2993 2447 2998 2452
rect 3657 2447 3790 2452
rect 2993 2442 3542 2447
rect 777 2437 926 2442
rect 1137 2437 1246 2442
rect 1353 2437 1358 2442
rect 2337 2437 2422 2442
rect 105 2432 166 2437
rect 313 2432 782 2437
rect 921 2432 1142 2437
rect 1353 2432 1382 2437
rect 1505 2432 2342 2437
rect 2417 2432 2454 2437
rect 2577 2432 2726 2437
rect 2913 2432 3094 2437
rect 3113 2432 3206 2437
rect 1377 2427 1510 2432
rect 2449 2427 2582 2432
rect 3089 2427 3094 2432
rect 97 2422 142 2427
rect 241 2422 294 2427
rect 337 2422 382 2427
rect 401 2422 926 2427
rect 1041 2422 1110 2427
rect 1129 2422 1230 2427
rect 1281 2422 1342 2427
rect 1529 2422 1574 2427
rect 1585 2422 1622 2427
rect 1633 2422 1686 2427
rect 289 2417 294 2422
rect 401 2417 406 2422
rect 921 2417 1046 2422
rect 1713 2417 1718 2427
rect 153 2412 174 2417
rect 193 2412 254 2417
rect 289 2412 406 2417
rect 449 2412 470 2417
rect 545 2412 854 2417
rect 881 2412 902 2417
rect 1065 2412 1158 2417
rect 849 2407 854 2412
rect 1265 2407 1270 2417
rect 1377 2412 1718 2417
rect 1729 2407 1734 2427
rect 1793 2422 1838 2427
rect 1897 2422 1934 2427
rect 2217 2422 2262 2427
rect 2353 2422 2406 2427
rect 2617 2422 2710 2427
rect 2961 2422 3030 2427
rect 3049 2422 3078 2427
rect 3089 2422 3174 2427
rect 3193 2422 3230 2427
rect 1953 2417 2150 2422
rect 3169 2417 3174 2422
rect 3281 2417 3286 2437
rect 3305 2432 3350 2437
rect 3441 2432 3462 2437
rect 3345 2417 3350 2432
rect 3369 2422 3438 2427
rect 1769 2412 1798 2417
rect 1881 2412 1958 2417
rect 2145 2412 2990 2417
rect 3065 2412 3094 2417
rect 3169 2412 3254 2417
rect 3281 2412 3310 2417
rect 3345 2412 3382 2417
rect 3457 2412 3462 2432
rect 1793 2407 1886 2412
rect 377 2402 494 2407
rect 649 2402 686 2407
rect 769 2402 830 2407
rect 849 2402 886 2407
rect 961 2402 1030 2407
rect 1233 2402 1270 2407
rect 1329 2402 1358 2407
rect 1657 2402 1734 2407
rect 1905 2402 2134 2407
rect 2257 2402 2278 2407
rect 2353 2402 2382 2407
rect 2721 2402 2750 2407
rect 2889 2402 2910 2407
rect 3033 2402 3078 2407
rect 3105 2402 3366 2407
rect 3377 2402 3382 2412
rect 3473 2402 3478 2437
rect 3553 2432 3590 2437
rect 3601 2432 3710 2437
rect 3785 2432 3926 2437
rect 3945 2432 4014 2437
rect 3945 2427 3950 2432
rect 3537 2417 3542 2427
rect 3641 2422 3678 2427
rect 3881 2422 3950 2427
rect 4009 2427 4014 2432
rect 4009 2422 4062 2427
rect 3521 2412 3542 2417
rect 3553 2412 3614 2417
rect 3873 2407 3878 2417
rect 3785 2402 3830 2407
rect 3873 2402 3894 2407
rect 3913 2402 3998 2407
rect 1489 2397 1558 2402
rect 2401 2397 2702 2402
rect 2769 2397 2870 2402
rect 3513 2397 3614 2402
rect 145 2392 278 2397
rect 385 2392 406 2397
rect 425 2392 462 2397
rect 553 2392 1222 2397
rect 1369 2392 1494 2397
rect 1553 2392 1854 2397
rect 1873 2392 1926 2397
rect 2097 2392 2406 2397
rect 2697 2392 2774 2397
rect 2865 2392 3246 2397
rect 3393 2392 3518 2397
rect 3609 2392 3742 2397
rect 3753 2392 3798 2397
rect 3825 2392 3886 2397
rect 1217 2387 1374 2392
rect 2009 2387 2078 2392
rect 3241 2387 3398 2392
rect 457 2382 646 2387
rect 665 2382 726 2387
rect 737 2382 830 2387
rect 881 2382 902 2387
rect 1505 2382 1542 2387
rect 1641 2382 1702 2387
rect 1745 2382 2014 2387
rect 2073 2382 2958 2387
rect 3065 2382 3102 2387
rect 3161 2382 3222 2387
rect 3529 2382 3598 2387
rect 3873 2382 3902 2387
rect 921 2377 1014 2382
rect 337 2372 758 2377
rect 769 2372 798 2377
rect 809 2372 926 2377
rect 1009 2372 1038 2377
rect 1065 2372 1126 2377
rect 1145 2372 1406 2377
rect 1425 2372 1510 2377
rect 1721 2372 1870 2377
rect 1881 2372 1918 2377
rect 2025 2372 2134 2377
rect 2329 2372 2398 2377
rect 2441 2372 2942 2377
rect 3009 2372 3070 2377
rect 3289 2372 3462 2377
rect 3729 2372 4094 2377
rect 1145 2367 1150 2372
rect 137 2362 190 2367
rect 305 2362 398 2367
rect 617 2362 926 2367
rect 961 2362 1062 2367
rect 1073 2362 1150 2367
rect 1401 2367 1406 2372
rect 1529 2367 1702 2372
rect 2153 2367 2310 2372
rect 3289 2367 3294 2372
rect 1401 2362 1534 2367
rect 1697 2362 2158 2367
rect 2305 2362 3294 2367
rect 3457 2367 3462 2372
rect 3457 2362 3486 2367
rect 393 2357 398 2362
rect 497 2357 622 2362
rect 1273 2357 1350 2362
rect 393 2352 502 2357
rect 641 2352 670 2357
rect 689 2352 870 2357
rect 897 2352 1278 2357
rect 1345 2352 1438 2357
rect 1521 2352 2670 2357
rect 2841 2352 2878 2357
rect 2937 2352 3054 2357
rect 3305 2352 3510 2357
rect 3553 2352 3662 2357
rect 3737 2352 3838 2357
rect 689 2347 694 2352
rect 2689 2347 2822 2352
rect 3553 2347 3558 2352
rect 161 2342 278 2347
rect 321 2342 374 2347
rect 521 2342 590 2347
rect 609 2342 694 2347
rect 713 2342 950 2347
rect 1057 2342 1094 2347
rect 1289 2342 1366 2347
rect 1425 2342 1462 2347
rect 1513 2342 1558 2347
rect 1633 2342 1742 2347
rect 1841 2342 1934 2347
rect 1961 2342 2694 2347
rect 2817 2342 2974 2347
rect 2985 2342 3414 2347
rect 521 2337 526 2342
rect 153 2332 342 2337
rect 497 2332 526 2337
rect 585 2337 590 2342
rect 3409 2337 3414 2342
rect 3537 2342 3558 2347
rect 3641 2342 3726 2347
rect 3537 2337 3542 2342
rect 585 2332 902 2337
rect 921 2332 1190 2337
rect 1417 2332 1446 2337
rect 1569 2332 3110 2337
rect 3265 2332 3326 2337
rect 3409 2332 3542 2337
rect 3721 2337 3726 2342
rect 3825 2342 3854 2347
rect 4041 2342 4142 2347
rect 3825 2337 3830 2342
rect 3721 2332 3830 2337
rect 361 2327 478 2332
rect 1209 2327 1318 2332
rect 1441 2327 1574 2332
rect 0 2322 366 2327
rect 473 2322 1214 2327
rect 1313 2322 1382 2327
rect 1601 2322 1638 2327
rect 1697 2322 1742 2327
rect 1849 2322 1934 2327
rect 2049 2322 2446 2327
rect 2553 2322 2598 2327
rect 2753 2322 3254 2327
rect 3361 2322 3390 2327
rect 2593 2317 2758 2322
rect 3249 2317 3366 2322
rect 3569 2317 3574 2327
rect 3873 2322 4014 2327
rect 3873 2317 3878 2322
rect 193 2312 254 2317
rect 353 2312 462 2317
rect 577 2312 630 2317
rect 649 2312 686 2317
rect 697 2312 758 2317
rect 769 2312 830 2317
rect 977 2312 1110 2317
rect 1217 2312 1302 2317
rect 1401 2312 1582 2317
rect 1777 2312 1830 2317
rect 2201 2312 2254 2317
rect 2393 2312 2454 2317
rect 2489 2312 2574 2317
rect 2777 2312 2822 2317
rect 2849 2312 2894 2317
rect 2969 2312 3062 2317
rect 3409 2312 3526 2317
rect 3545 2312 3574 2317
rect 3593 2312 3686 2317
rect 3705 2312 3774 2317
rect 3841 2312 3878 2317
rect 4009 2317 4014 2322
rect 4009 2312 4062 2317
rect 753 2307 758 2312
rect 849 2307 950 2312
rect 1321 2307 1406 2312
rect 1577 2307 1582 2312
rect 1849 2307 2182 2312
rect 2273 2307 2374 2312
rect 3409 2307 3414 2312
rect 241 2302 406 2307
rect 673 2302 718 2307
rect 753 2302 854 2307
rect 945 2302 974 2307
rect 1001 2302 1326 2307
rect 1577 2302 1854 2307
rect 2177 2302 2278 2307
rect 2369 2302 2958 2307
rect 401 2297 406 2302
rect 489 2297 654 2302
rect 2953 2297 2958 2302
rect 3073 2302 3414 2307
rect 3521 2307 3526 2312
rect 3593 2307 3598 2312
rect 3521 2302 3598 2307
rect 3681 2307 3686 2312
rect 3681 2302 3758 2307
rect 3073 2297 3078 2302
rect 401 2292 494 2297
rect 649 2292 710 2297
rect 745 2292 798 2297
rect 817 2292 854 2297
rect 865 2292 982 2297
rect 1153 2292 1566 2297
rect 1817 2292 1902 2297
rect 1929 2292 2430 2297
rect 2537 2292 2582 2297
rect 2745 2292 2862 2297
rect 2953 2292 3078 2297
rect 3169 2292 3198 2297
rect 1001 2287 1158 2292
rect 1561 2287 1702 2292
rect 3193 2287 3198 2292
rect 3425 2292 3670 2297
rect 3425 2287 3430 2292
rect 3665 2287 3670 2292
rect 3769 2292 3998 2297
rect 3769 2287 3774 2292
rect 505 2282 1006 2287
rect 1169 2282 1214 2287
rect 1265 2282 1358 2287
rect 1697 2282 1870 2287
rect 1953 2282 2158 2287
rect 2385 2282 2478 2287
rect 2657 2282 2718 2287
rect 3193 2282 3430 2287
rect 3449 2282 3478 2287
rect 3505 2282 3638 2287
rect 3665 2282 3774 2287
rect 4009 2282 4046 2287
rect 1865 2277 1958 2282
rect 2153 2277 2390 2282
rect 2497 2277 2598 2282
rect 313 2272 454 2277
rect 449 2267 454 2272
rect 737 2272 1214 2277
rect 1369 2272 1526 2277
rect 1577 2272 1678 2277
rect 1809 2272 1846 2277
rect 2409 2272 2502 2277
rect 2593 2272 2622 2277
rect 2737 2272 2846 2277
rect 2881 2272 3006 2277
rect 3025 2272 3070 2277
rect 737 2267 742 2272
rect 1209 2267 1374 2272
rect 1577 2267 1582 2272
rect 393 2262 430 2267
rect 449 2262 742 2267
rect 761 2262 1134 2267
rect 1145 2262 1190 2267
rect 1185 2257 1190 2262
rect 1537 2262 1582 2267
rect 1673 2267 1678 2272
rect 1977 2267 2134 2272
rect 2881 2267 2886 2272
rect 1673 2262 1798 2267
rect 1857 2262 1982 2267
rect 2129 2262 2886 2267
rect 3001 2267 3006 2272
rect 3633 2267 3638 2282
rect 4009 2267 4014 2282
rect 3001 2262 3438 2267
rect 1537 2257 1542 2262
rect 1793 2257 1862 2262
rect 3433 2257 3438 2262
rect 3521 2262 3614 2267
rect 3633 2262 4014 2267
rect 3521 2257 3526 2262
rect 225 2252 302 2257
rect 769 2252 1054 2257
rect 1185 2252 1542 2257
rect 1593 2252 1662 2257
rect 1993 2252 2054 2257
rect 2081 2252 2118 2257
rect 2585 2252 2790 2257
rect 2897 2252 3054 2257
rect 3433 2252 3526 2257
rect 2409 2247 2566 2252
rect 641 2242 710 2247
rect 857 2242 886 2247
rect 961 2242 1054 2247
rect 1073 2242 1166 2247
rect 1657 2242 1774 2247
rect 1793 2242 1974 2247
rect 2057 2242 2118 2247
rect 2201 2242 2414 2247
rect 2561 2242 2590 2247
rect 2609 2242 3358 2247
rect 1073 2237 1078 2242
rect 169 2232 206 2237
rect 409 2232 446 2237
rect 473 2232 558 2237
rect 865 2232 950 2237
rect 1009 2232 1078 2237
rect 1161 2237 1166 2242
rect 1793 2237 1798 2242
rect 1161 2232 1798 2237
rect 1969 2237 1974 2242
rect 2609 2237 2614 2242
rect 1969 2232 2190 2237
rect 2345 2232 2614 2237
rect 2665 2232 2766 2237
rect 2785 2232 2814 2237
rect 2961 2232 3030 2237
rect 3545 2232 3638 2237
rect 945 2227 1014 2232
rect 2185 2227 2350 2232
rect 409 2222 526 2227
rect 641 2222 678 2227
rect 1033 2222 1086 2227
rect 1105 2222 1150 2227
rect 1617 2222 2158 2227
rect 2369 2222 2422 2227
rect 2457 2222 2502 2227
rect 2729 2222 2758 2227
rect 2769 2222 2814 2227
rect 1105 2217 1110 2222
rect 289 2212 390 2217
rect 505 2212 1110 2217
rect 1137 2212 1254 2217
rect 1649 2212 1686 2217
rect 1713 2212 1758 2217
rect 1769 2212 1846 2217
rect 1929 2212 1974 2217
rect 2049 2212 2078 2217
rect 2105 2212 2294 2217
rect 2361 2212 2566 2217
rect 2585 2212 2710 2217
rect 2841 2212 2942 2217
rect 289 2207 294 2212
rect 265 2202 294 2207
rect 385 2207 390 2212
rect 385 2202 558 2207
rect 993 2202 1110 2207
rect 649 2197 718 2202
rect 81 2192 182 2197
rect 193 2192 222 2197
rect 289 2192 350 2197
rect 457 2192 486 2197
rect 545 2192 654 2197
rect 713 2192 742 2197
rect 833 2192 870 2197
rect 1033 2192 1102 2197
rect 345 2187 462 2192
rect 665 2182 702 2187
rect 833 2182 878 2187
rect 1137 2182 1142 2212
rect 2585 2207 2590 2212
rect 2705 2207 2774 2212
rect 2841 2207 2846 2212
rect 1337 2202 2190 2207
rect 2185 2197 2190 2202
rect 2289 2202 2590 2207
rect 2769 2202 2846 2207
rect 2937 2207 2942 2212
rect 3049 2212 3246 2217
rect 3049 2207 3054 2212
rect 2937 2202 3054 2207
rect 3241 2207 3246 2212
rect 3369 2212 3622 2217
rect 3369 2207 3374 2212
rect 3241 2202 3374 2207
rect 3617 2207 3622 2212
rect 3617 2202 3646 2207
rect 3833 2202 3870 2207
rect 3889 2202 3966 2207
rect 2289 2197 2294 2202
rect 3889 2197 3894 2202
rect 1161 2192 1254 2197
rect 1361 2192 1406 2197
rect 1593 2192 1630 2197
rect 1665 2192 1966 2197
rect 1961 2187 1966 2192
rect 2081 2192 2110 2197
rect 2185 2192 2294 2197
rect 2393 2192 2510 2197
rect 2585 2192 2678 2197
rect 2697 2192 2758 2197
rect 2857 2192 3118 2197
rect 3169 2192 3230 2197
rect 3433 2192 3510 2197
rect 3521 2192 3790 2197
rect 3809 2192 3894 2197
rect 3961 2197 3966 2202
rect 3961 2192 3990 2197
rect 4001 2192 4062 2197
rect 2081 2187 2086 2192
rect 3169 2187 3174 2192
rect 3521 2187 3526 2192
rect 3809 2187 3814 2192
rect 1225 2182 1254 2187
rect 1409 2182 1670 2187
rect 1777 2182 1846 2187
rect 1961 2182 2086 2187
rect 2353 2182 2414 2187
rect 2425 2182 2502 2187
rect 2665 2182 2782 2187
rect 2977 2182 3174 2187
rect 3385 2182 3526 2187
rect 3649 2182 3694 2187
rect 3713 2182 3814 2187
rect 3897 2182 4070 2187
rect 489 2177 590 2182
rect 385 2172 494 2177
rect 585 2172 614 2177
rect 961 2172 1094 2177
rect 1649 2172 1702 2177
rect 1769 2172 1870 2177
rect 2121 2172 2166 2177
rect 2313 2172 2574 2177
rect 2609 2172 2678 2177
rect 2713 2172 2734 2177
rect 2913 2172 2998 2177
rect 3137 2172 3774 2177
rect 3809 2172 4134 2177
rect 633 2167 782 2172
rect 3017 2167 3110 2172
rect 257 2162 374 2167
rect 505 2162 638 2167
rect 777 2162 1014 2167
rect 1425 2162 1510 2167
rect 1553 2162 1606 2167
rect 1697 2162 1742 2167
rect 1793 2162 1838 2167
rect 1961 2162 2006 2167
rect 2105 2162 2142 2167
rect 2249 2162 2494 2167
rect 2705 2162 2782 2167
rect 2801 2162 2878 2167
rect 2945 2162 3022 2167
rect 3105 2162 3134 2167
rect 3569 2162 4046 2167
rect 369 2157 510 2162
rect 1009 2157 1118 2162
rect 529 2152 766 2157
rect 1113 2152 1950 2157
rect 2017 2152 2518 2157
rect 2609 2152 2630 2157
rect 2657 2152 2726 2157
rect 1945 2147 2022 2152
rect 2801 2147 2806 2162
rect 2873 2157 2878 2162
rect 3153 2157 3406 2162
rect 3441 2157 3550 2162
rect 2873 2152 2934 2157
rect 2993 2152 3158 2157
rect 3401 2152 3446 2157
rect 3545 2152 3606 2157
rect 3681 2152 3718 2157
rect 3785 2152 3902 2157
rect 2929 2147 2998 2152
rect 161 2142 222 2147
rect 265 2142 366 2147
rect 409 2142 518 2147
rect 561 2142 606 2147
rect 633 2142 702 2147
rect 977 2142 1102 2147
rect 1489 2142 1518 2147
rect 1713 2142 1846 2147
rect 1889 2142 1918 2147
rect 2137 2142 2198 2147
rect 2305 2142 2326 2147
rect 2385 2142 2422 2147
rect 2481 2142 2622 2147
rect 1513 2137 1614 2142
rect 1713 2137 1718 2142
rect 2321 2137 2326 2142
rect 2617 2137 2622 2142
rect 2737 2142 2806 2147
rect 2825 2142 2862 2147
rect 3017 2142 3286 2147
rect 3297 2142 3390 2147
rect 3457 2142 3718 2147
rect 3817 2142 3942 2147
rect 4025 2142 4094 2147
rect 2737 2137 2742 2142
rect 3281 2137 3286 2142
rect 3457 2137 3462 2142
rect 137 2132 206 2137
rect 241 2132 310 2137
rect 457 2132 630 2137
rect 713 2132 878 2137
rect 937 2132 1022 2137
rect 1265 2132 1342 2137
rect 1609 2132 1718 2137
rect 1873 2132 1910 2137
rect 2041 2132 2118 2137
rect 2233 2132 2294 2137
rect 2321 2132 2398 2137
rect 2465 2132 2550 2137
rect 2617 2132 2742 2137
rect 2929 2132 2950 2137
rect 2969 2132 3158 2137
rect 3201 2132 3262 2137
rect 3281 2132 3486 2137
rect 3497 2132 3566 2137
rect 3609 2132 3790 2137
rect 3857 2132 3926 2137
rect 305 2127 462 2132
rect 625 2127 718 2132
rect 1265 2127 1270 2132
rect 105 2122 222 2127
rect 249 2122 286 2127
rect 481 2122 510 2127
rect 505 2117 510 2122
rect 569 2122 606 2127
rect 809 2122 902 2127
rect 953 2122 1182 2127
rect 1241 2122 1270 2127
rect 1337 2127 1342 2132
rect 1873 2127 1878 2132
rect 2041 2127 2046 2132
rect 2113 2127 2214 2132
rect 2465 2127 2470 2132
rect 1337 2122 1366 2127
rect 1553 2122 1590 2127
rect 1857 2122 1878 2127
rect 1889 2122 2046 2127
rect 2209 2122 2470 2127
rect 2481 2122 2598 2127
rect 2889 2122 3006 2127
rect 3033 2122 3062 2127
rect 3121 2122 3334 2127
rect 3617 2122 3638 2127
rect 3713 2122 3886 2127
rect 569 2117 574 2122
rect 1889 2117 1894 2122
rect 145 2112 174 2117
rect 193 2112 262 2117
rect 345 2112 406 2117
rect 505 2112 574 2117
rect 593 2112 638 2117
rect 689 2112 766 2117
rect 889 2112 910 2117
rect 1257 2112 1374 2117
rect 1465 2112 1510 2117
rect 1577 2112 1622 2117
rect 1737 2112 1774 2117
rect 1841 2112 1894 2117
rect 1905 2112 1950 2117
rect 2041 2112 2102 2117
rect 2129 2112 2158 2117
rect 2185 2112 2230 2117
rect 2329 2112 2558 2117
rect 2569 2112 2630 2117
rect 2649 2112 2798 2117
rect 2817 2112 2846 2117
rect 2865 2112 3030 2117
rect 3089 2112 3214 2117
rect 3225 2112 3286 2117
rect 689 2107 694 2112
rect 201 2102 230 2107
rect 241 2102 318 2107
rect 377 2102 462 2107
rect 665 2102 694 2107
rect 761 2107 766 2112
rect 1153 2107 1238 2112
rect 2649 2107 2654 2112
rect 761 2102 1158 2107
rect 1233 2102 1318 2107
rect 1385 2102 1454 2107
rect 1521 2102 1566 2107
rect 1633 2102 1830 2107
rect 1961 2102 2654 2107
rect 2793 2107 2798 2112
rect 3281 2107 3286 2112
rect 3345 2112 3686 2117
rect 3705 2112 3782 2117
rect 3833 2112 3878 2117
rect 3913 2112 3982 2117
rect 3345 2107 3350 2112
rect 2793 2102 3198 2107
rect 3281 2102 3350 2107
rect 3665 2102 3830 2107
rect 1313 2097 1390 2102
rect 1449 2097 1526 2102
rect 1561 2097 1638 2102
rect 1825 2097 1966 2102
rect 705 2092 750 2097
rect 1169 2092 1206 2097
rect 1217 2092 1294 2097
rect 1721 2092 1798 2097
rect 1993 2092 2070 2097
rect 2113 2092 2166 2097
rect 2345 2092 2430 2097
rect 2521 2092 2742 2097
rect 2929 2092 3022 2097
rect 3073 2092 3190 2097
rect 3545 2092 3894 2097
rect 985 2087 1150 2092
rect 2425 2087 2526 2092
rect 2769 2087 2910 2092
rect 289 2082 318 2087
rect 313 2077 318 2082
rect 393 2082 486 2087
rect 537 2082 654 2087
rect 393 2077 398 2082
rect 313 2072 398 2077
rect 649 2077 654 2082
rect 961 2082 990 2087
rect 1145 2082 1318 2087
rect 1337 2082 1574 2087
rect 1593 2082 1638 2087
rect 1697 2082 1734 2087
rect 1817 2082 1926 2087
rect 2313 2082 2406 2087
rect 2545 2082 2726 2087
rect 2745 2082 2774 2087
rect 2905 2082 3558 2087
rect 961 2077 966 2082
rect 1337 2077 1342 2082
rect 649 2072 966 2077
rect 985 2072 1342 2077
rect 1569 2077 1574 2082
rect 1817 2077 1822 2082
rect 1569 2072 1822 2077
rect 1921 2077 1926 2082
rect 2721 2077 2726 2082
rect 3553 2077 3558 2082
rect 3633 2082 3662 2087
rect 3681 2082 3750 2087
rect 3769 2082 3846 2087
rect 3633 2077 3638 2082
rect 1921 2072 2694 2077
rect 2721 2072 2934 2077
rect 2977 2072 3222 2077
rect 3553 2072 3638 2077
rect 3745 2077 3750 2082
rect 3745 2072 3854 2077
rect 1465 2067 1550 2072
rect 2689 2067 2694 2072
rect 1065 2062 1206 2067
rect 1353 2062 1470 2067
rect 1545 2062 1910 2067
rect 2377 2062 2422 2067
rect 2569 2062 2670 2067
rect 2689 2062 3038 2067
rect 3129 2062 3302 2067
rect 3353 2062 3422 2067
rect 3441 2062 3534 2067
rect 3745 2062 3766 2067
rect 1201 2057 1358 2062
rect 3353 2057 3358 2062
rect 1481 2052 1542 2057
rect 2105 2052 2254 2057
rect 2473 2052 2494 2057
rect 2577 2052 2614 2057
rect 2625 2052 3358 2057
rect 3417 2057 3422 2062
rect 3417 2052 3486 2057
rect 1065 2047 1182 2052
rect 1561 2047 1694 2052
rect 1777 2047 1918 2052
rect 2105 2047 2110 2052
rect 785 2042 1070 2047
rect 1177 2042 1350 2047
rect 1345 2037 1350 2042
rect 1449 2042 1566 2047
rect 1689 2042 1782 2047
rect 1913 2042 2110 2047
rect 2249 2047 2254 2052
rect 3481 2047 3486 2052
rect 3545 2052 3766 2057
rect 3545 2047 3550 2052
rect 2249 2042 2766 2047
rect 3153 2042 3270 2047
rect 3369 2042 3438 2047
rect 1449 2037 1454 2042
rect 2889 2037 2974 2042
rect 3457 2037 3462 2047
rect 3481 2042 3550 2047
rect 3705 2042 3806 2047
rect 3857 2042 3942 2047
rect 3857 2037 3862 2042
rect 193 2032 390 2037
rect 457 2032 526 2037
rect 1081 2032 1166 2037
rect 1345 2032 1454 2037
rect 1529 2032 1582 2037
rect 1641 2032 1678 2037
rect 1793 2032 1902 2037
rect 2121 2032 2238 2037
rect 2561 2032 2894 2037
rect 2969 2032 3462 2037
rect 3833 2032 3862 2037
rect 3937 2037 3942 2042
rect 3937 2032 4006 2037
rect 4033 2032 4142 2037
rect 1921 2027 2014 2032
rect 113 2022 174 2027
rect 185 2022 214 2027
rect 513 2022 558 2027
rect 713 2022 806 2027
rect 1289 2022 1318 2027
rect 1625 2022 1694 2027
rect 1873 2022 1926 2027
rect 2009 2022 2038 2027
rect 2105 2022 2142 2027
rect 2153 2022 2182 2027
rect 1153 2017 1246 2022
rect 1713 2017 1854 2022
rect 577 2012 694 2017
rect 897 2012 1022 2017
rect 1129 2012 1158 2017
rect 1241 2012 1326 2017
rect 1473 2012 1718 2017
rect 1849 2012 2126 2017
rect 577 2007 582 2012
rect 433 2002 582 2007
rect 689 2007 694 2012
rect 689 2002 774 2007
rect 1121 2002 1230 2007
rect 1305 2002 1414 2007
rect 1561 2002 1582 2007
rect 1641 2002 1710 2007
rect 1753 2002 1942 2007
rect 2033 2002 2230 2007
rect 2241 2002 2246 2027
rect 2257 2022 2326 2027
rect 2393 2022 2478 2027
rect 2497 2022 2582 2027
rect 2601 2022 2646 2027
rect 2697 2022 2726 2027
rect 2905 2022 2958 2027
rect 3145 2022 3230 2027
rect 3257 2022 3430 2027
rect 3465 2022 3518 2027
rect 3633 2022 3702 2027
rect 3769 2022 3830 2027
rect 3977 2022 4006 2027
rect 2393 2017 2398 2022
rect 2265 2012 2398 2017
rect 2473 2017 2478 2022
rect 2801 2017 2886 2022
rect 3633 2017 3638 2022
rect 2473 2012 2806 2017
rect 2881 2012 3118 2017
rect 3217 2012 3310 2017
rect 3505 2012 3638 2017
rect 3801 2012 4038 2017
rect 2409 2002 2750 2007
rect 2817 2002 2942 2007
rect 3081 2002 3142 2007
rect 3289 2002 3358 2007
rect 3393 2002 3470 2007
rect 857 1997 1046 2002
rect 161 1992 342 1997
rect 689 1992 726 1997
rect 753 1992 862 1997
rect 1041 1992 1070 1997
rect 1121 1992 1126 2002
rect 1473 1997 1542 2002
rect 1937 1997 2038 2002
rect 1201 1992 1478 1997
rect 1537 1992 1638 1997
rect 1889 1992 1918 1997
rect 2057 1992 2278 1997
rect 2361 1992 2726 1997
rect 2881 1992 2966 1997
rect 3105 1992 3142 1997
rect 3241 1992 3270 1997
rect 3297 1992 3382 1997
rect 393 1987 606 1992
rect 1633 1987 1894 1992
rect 2273 1987 2278 1992
rect 2745 1987 2862 1992
rect 3393 1987 3398 2002
rect 3553 1992 3614 1997
rect 3737 1992 3822 1997
rect 3833 1992 3854 1997
rect 3865 1992 3926 1997
rect 4017 1992 4078 1997
rect 177 1982 238 1987
rect 369 1982 398 1987
rect 601 1982 630 1987
rect 649 1982 686 1987
rect 873 1982 1270 1987
rect 1281 1982 1334 1987
rect 1489 1982 1534 1987
rect 1577 1982 1614 1987
rect 1913 1982 1966 1987
rect 2153 1982 2182 1987
rect 2233 1982 2262 1987
rect 2273 1982 2390 1987
rect 2449 1982 2510 1987
rect 2545 1982 2750 1987
rect 2857 1982 3094 1987
rect 3209 1982 3334 1987
rect 3345 1982 3398 1987
rect 3449 1982 3502 1987
rect 3841 1982 3998 1987
rect 4009 1982 4038 1987
rect 1353 1977 1454 1982
rect 385 1972 1358 1977
rect 1449 1972 1478 1977
rect 1513 1972 1814 1977
rect 1873 1972 1958 1977
rect 2001 1972 2118 1977
rect 2353 1972 2414 1977
rect 2521 1972 2574 1977
rect 2601 1972 2662 1977
rect 2721 1972 3038 1977
rect 3049 1972 3438 1977
rect 3465 1972 3510 1977
rect 3673 1972 3958 1977
rect 193 1962 262 1967
rect 497 1962 726 1967
rect 833 1962 998 1967
rect 1113 1962 1262 1967
rect 1313 1962 1374 1967
rect 1385 1962 1462 1967
rect 1529 1962 1646 1967
rect 2089 1962 2126 1967
rect 2145 1962 2286 1967
rect 2385 1962 2542 1967
rect 2561 1962 2646 1967
rect 2705 1962 2742 1967
rect 2753 1962 2894 1967
rect 3273 1962 3550 1967
rect 3833 1962 3886 1967
rect 3905 1962 4046 1967
rect 297 1957 406 1962
rect 1665 1957 1814 1962
rect 1889 1957 2070 1962
rect 2145 1957 2150 1962
rect 81 1952 238 1957
rect 273 1952 302 1957
rect 401 1952 486 1957
rect 505 1952 1518 1957
rect 1569 1952 1670 1957
rect 1809 1952 1894 1957
rect 2065 1952 2150 1957
rect 2281 1957 2286 1962
rect 2753 1957 2758 1962
rect 2281 1952 2758 1957
rect 2865 1952 2958 1957
rect 3065 1952 3094 1957
rect 3321 1952 3366 1957
rect 3401 1952 3574 1957
rect 3825 1952 4030 1957
rect 4049 1952 4134 1957
rect 481 1947 486 1952
rect 3089 1947 3094 1952
rect 145 1942 190 1947
rect 209 1942 462 1947
rect 481 1942 582 1947
rect 609 1942 702 1947
rect 833 1942 878 1947
rect 969 1942 1014 1947
rect 1057 1942 1094 1947
rect 1113 1942 1174 1947
rect 1185 1942 1310 1947
rect 1369 1942 1446 1947
rect 1537 1942 1566 1947
rect 1601 1942 1726 1947
rect 1745 1942 1798 1947
rect 1905 1942 1958 1947
rect 1977 1942 2086 1947
rect 2113 1942 2270 1947
rect 2425 1942 2534 1947
rect 2609 1942 2902 1947
rect 2913 1942 2942 1947
rect 2953 1942 3070 1947
rect 3089 1942 3222 1947
rect 3265 1942 3366 1947
rect 3425 1942 3510 1947
rect 3537 1942 3574 1947
rect 3713 1942 3854 1947
rect 3873 1942 3910 1947
rect 4001 1942 4094 1947
rect 313 1932 414 1937
rect 513 1932 622 1937
rect 657 1932 726 1937
rect 889 1932 958 1937
rect 953 1927 958 1932
rect 1041 1932 1678 1937
rect 1697 1932 1718 1937
rect 1041 1927 1046 1932
rect 1745 1927 1750 1942
rect 1953 1937 1958 1942
rect 2289 1937 2406 1942
rect 1953 1932 2142 1937
rect 2241 1932 2294 1937
rect 2401 1932 2566 1937
rect 2137 1927 2246 1932
rect 2609 1927 2614 1942
rect 3505 1937 3510 1942
rect 2633 1932 2766 1937
rect 2801 1932 2838 1937
rect 3025 1932 3422 1937
rect 3505 1932 3534 1937
rect 3561 1932 3638 1937
rect 2857 1927 3006 1932
rect 3761 1927 3870 1932
rect 145 1922 198 1927
rect 417 1922 502 1927
rect 577 1922 646 1927
rect 953 1922 1046 1927
rect 1065 1922 1086 1927
rect 1153 1922 1494 1927
rect 1633 1922 1750 1927
rect 1993 1922 2062 1927
rect 2097 1922 2118 1927
rect 2265 1922 2614 1927
rect 2625 1922 2686 1927
rect 2777 1922 2862 1927
rect 3001 1922 3638 1927
rect 3665 1922 3766 1927
rect 3865 1922 3894 1927
rect 641 1917 646 1922
rect 1513 1917 1614 1922
rect 121 1912 174 1917
rect 185 1912 278 1917
rect 409 1912 454 1917
rect 585 1912 630 1917
rect 641 1912 662 1917
rect 705 1912 774 1917
rect 889 1912 918 1917
rect 1081 1912 1118 1917
rect 1185 1912 1230 1917
rect 1265 1912 1518 1917
rect 1609 1912 1982 1917
rect 2081 1912 2630 1917
rect 2673 1912 2750 1917
rect 2857 1912 3030 1917
rect 3073 1912 3454 1917
rect 3481 1912 3542 1917
rect 3553 1912 3614 1917
rect 3777 1912 3846 1917
rect 3865 1912 3918 1917
rect 1977 1907 2086 1912
rect 161 1902 214 1907
rect 489 1902 574 1907
rect 649 1902 1070 1907
rect 1129 1902 1222 1907
rect 1313 1902 1638 1907
rect 1657 1902 1686 1907
rect 1761 1902 1806 1907
rect 2105 1902 2142 1907
rect 2241 1902 2358 1907
rect 2377 1902 2422 1907
rect 2473 1902 2550 1907
rect 2625 1902 2630 1912
rect 2945 1902 2974 1907
rect 3049 1902 3142 1907
rect 3313 1902 3414 1907
rect 3641 1902 3806 1907
rect 569 1897 654 1902
rect 1065 1897 1134 1902
rect 1217 1897 1318 1902
rect 1825 1897 1958 1902
rect 2625 1897 2838 1902
rect 3161 1897 3278 1902
rect 481 1892 534 1897
rect 801 1892 830 1897
rect 873 1892 902 1897
rect 1153 1892 1198 1897
rect 1457 1892 1830 1897
rect 1953 1892 1982 1897
rect 2041 1892 2070 1897
rect 2833 1892 3166 1897
rect 3273 1892 3302 1897
rect 529 1887 534 1892
rect 673 1887 806 1892
rect 1337 1887 1438 1892
rect 2193 1887 2606 1892
rect 3297 1887 3302 1892
rect 3409 1892 3486 1897
rect 3545 1892 3710 1897
rect 3409 1887 3414 1892
rect 457 1882 510 1887
rect 529 1882 678 1887
rect 969 1882 1342 1887
rect 1433 1882 1502 1887
rect 1641 1882 2198 1887
rect 2601 1882 2822 1887
rect 3009 1882 3158 1887
rect 3201 1882 3270 1887
rect 3297 1882 3414 1887
rect 3433 1882 3742 1887
rect 1497 1877 1646 1882
rect 2817 1877 3014 1882
rect 697 1872 910 1877
rect 1169 1872 1206 1877
rect 1353 1872 1406 1877
rect 1425 1872 1478 1877
rect 1665 1872 1782 1877
rect 1889 1872 1990 1877
rect 2209 1872 2798 1877
rect 3033 1872 3062 1877
rect 3145 1872 3246 1877
rect 3497 1872 3678 1877
rect 3689 1872 3766 1877
rect 2097 1867 2190 1872
rect 929 1862 1150 1867
rect 681 1857 934 1862
rect 1145 1857 1150 1862
rect 1225 1862 1334 1867
rect 1497 1862 1646 1867
rect 1673 1862 2102 1867
rect 2185 1862 3558 1867
rect 3873 1862 3966 1867
rect 1225 1857 1230 1862
rect 1329 1857 1502 1862
rect 1641 1857 1646 1862
rect 3873 1857 3878 1862
rect 321 1852 422 1857
rect 657 1852 686 1857
rect 1145 1852 1230 1857
rect 1641 1852 1742 1857
rect 1777 1852 2014 1857
rect 2113 1852 2142 1857
rect 2153 1852 2734 1857
rect 3033 1852 3118 1857
rect 3249 1852 3278 1857
rect 3465 1852 3574 1857
rect 3649 1852 3838 1857
rect 3849 1852 3878 1857
rect 3961 1857 3966 1862
rect 3961 1852 3990 1857
rect 321 1837 326 1852
rect 417 1847 422 1852
rect 2929 1847 3014 1852
rect 3137 1847 3230 1852
rect 3297 1847 3422 1852
rect 417 1842 446 1847
rect 601 1842 974 1847
rect 1033 1842 1062 1847
rect 1089 1842 1206 1847
rect 1257 1842 1398 1847
rect 1409 1842 1766 1847
rect 1793 1842 1862 1847
rect 2033 1842 2062 1847
rect 2073 1842 2542 1847
rect 2745 1842 2934 1847
rect 3009 1842 3142 1847
rect 3225 1842 3302 1847
rect 3417 1842 3686 1847
rect 3785 1842 3902 1847
rect 3921 1842 4142 1847
rect 1881 1837 2014 1842
rect 2537 1837 2750 1842
rect 161 1832 326 1837
rect 417 1832 662 1837
rect 753 1832 798 1837
rect 929 1832 1454 1837
rect 1841 1832 1886 1837
rect 2009 1832 2158 1837
rect 2201 1832 2254 1837
rect 2945 1832 2990 1837
rect 3041 1832 3102 1837
rect 3161 1832 3206 1837
rect 3249 1832 3406 1837
rect 3521 1832 3614 1837
rect 3689 1832 3774 1837
rect 3865 1832 3918 1837
rect 417 1827 422 1832
rect 817 1827 910 1832
rect 1449 1827 1846 1832
rect 2273 1827 2518 1832
rect 2841 1827 2926 1832
rect 3769 1827 3870 1832
rect 113 1822 174 1827
rect 201 1822 294 1827
rect 305 1822 334 1827
rect 345 1822 422 1827
rect 577 1822 630 1827
rect 769 1822 822 1827
rect 905 1822 1430 1827
rect 1865 1822 2278 1827
rect 2513 1822 2846 1827
rect 2921 1822 3150 1827
rect 3249 1822 3326 1827
rect 3417 1822 3718 1827
rect 3889 1822 3942 1827
rect 4025 1822 4094 1827
rect 353 1812 382 1817
rect 641 1812 678 1817
rect 801 1812 1070 1817
rect 1185 1812 1374 1817
rect 1425 1807 1430 1822
rect 3145 1817 3254 1822
rect 3321 1817 3422 1822
rect 4025 1817 4030 1822
rect 1441 1812 1646 1817
rect 1745 1812 1990 1817
rect 2129 1812 2502 1817
rect 2857 1812 3014 1817
rect 1441 1807 1446 1812
rect 345 1802 374 1807
rect 817 1802 838 1807
rect 897 1802 1246 1807
rect 1377 1802 1414 1807
rect 1425 1802 1446 1807
rect 1641 1807 1646 1812
rect 1985 1807 2134 1812
rect 2497 1807 2694 1812
rect 1641 1802 1886 1807
rect 1921 1802 1966 1807
rect 2153 1802 2478 1807
rect 657 1797 798 1802
rect 1481 1797 1606 1802
rect 2689 1797 2694 1807
rect 2857 1797 2862 1812
rect 3009 1807 3014 1812
rect 3273 1812 3302 1817
rect 3441 1812 3494 1817
rect 3273 1807 3278 1812
rect 3505 1807 3510 1817
rect 3569 1812 3598 1817
rect 3681 1812 3710 1817
rect 3793 1812 3830 1817
rect 3841 1812 4030 1817
rect 4089 1817 4094 1822
rect 4089 1812 4126 1817
rect 3593 1807 3686 1812
rect 3825 1807 3830 1812
rect 2929 1802 2990 1807
rect 3009 1802 3278 1807
rect 3353 1802 3446 1807
rect 3505 1802 3534 1807
rect 3721 1802 3806 1807
rect 3825 1802 3902 1807
rect 4009 1802 4078 1807
rect 3441 1797 3446 1802
rect 257 1792 342 1797
rect 377 1792 414 1797
rect 633 1792 662 1797
rect 793 1792 822 1797
rect 961 1792 990 1797
rect 1017 1792 1094 1797
rect 1169 1792 1230 1797
rect 1321 1792 1366 1797
rect 817 1787 966 1792
rect 1089 1787 1094 1792
rect 1361 1787 1366 1792
rect 1457 1792 1486 1797
rect 1601 1792 1630 1797
rect 1857 1792 1886 1797
rect 2089 1792 2134 1797
rect 2225 1792 2438 1797
rect 2457 1792 2542 1797
rect 2641 1792 2670 1797
rect 2689 1792 2862 1797
rect 2881 1792 2950 1797
rect 3361 1792 3430 1797
rect 3441 1792 3494 1797
rect 3521 1792 3782 1797
rect 3841 1792 3990 1797
rect 4073 1792 4158 1797
rect 1457 1787 1462 1792
rect 1721 1787 1838 1792
rect 2225 1787 2230 1792
rect 2433 1787 2438 1792
rect 201 1782 230 1787
rect 281 1782 326 1787
rect 609 1782 798 1787
rect 1089 1782 1214 1787
rect 1361 1782 1462 1787
rect 1481 1782 1526 1787
rect 1537 1782 1598 1787
rect 1697 1782 1726 1787
rect 1833 1782 1870 1787
rect 1937 1782 2070 1787
rect 2113 1782 2230 1787
rect 2249 1782 2342 1787
rect 2433 1782 2558 1787
rect 3145 1782 3214 1787
rect 3393 1782 3518 1787
rect 3561 1782 3614 1787
rect 3769 1782 3934 1787
rect 1937 1777 1942 1782
rect 689 1772 726 1777
rect 809 1772 902 1777
rect 969 1772 1342 1777
rect 1481 1772 1566 1777
rect 1601 1772 1942 1777
rect 2065 1777 2070 1782
rect 3145 1777 3150 1782
rect 2065 1772 2158 1777
rect 2233 1772 2270 1777
rect 2353 1772 2398 1777
rect 2585 1772 2662 1777
rect 3001 1772 3150 1777
rect 3209 1777 3214 1782
rect 3305 1777 3374 1782
rect 3209 1772 3310 1777
rect 3369 1772 3422 1777
rect 3465 1772 3526 1777
rect 3777 1772 3886 1777
rect 737 1767 814 1772
rect 897 1767 902 1772
rect 2433 1767 2542 1772
rect 249 1762 318 1767
rect 345 1762 430 1767
rect 505 1762 542 1767
rect 657 1762 742 1767
rect 857 1762 886 1767
rect 897 1762 958 1767
rect 345 1757 350 1762
rect 281 1752 350 1757
rect 425 1757 430 1762
rect 953 1757 958 1762
rect 1089 1762 1470 1767
rect 1529 1762 1726 1767
rect 1945 1762 2342 1767
rect 2409 1762 2438 1767
rect 2537 1762 2710 1767
rect 3321 1762 3438 1767
rect 3457 1762 3502 1767
rect 3537 1762 3566 1767
rect 3729 1762 3758 1767
rect 4033 1762 4086 1767
rect 1089 1757 1094 1762
rect 1465 1757 1534 1762
rect 2337 1757 2414 1762
rect 3457 1757 3462 1762
rect 425 1752 454 1757
rect 641 1752 822 1757
rect 865 1752 902 1757
rect 953 1752 1094 1757
rect 1113 1752 1214 1757
rect 1233 1752 1382 1757
rect 1553 1752 1582 1757
rect 1713 1752 1742 1757
rect 1753 1752 2118 1757
rect 2129 1752 2166 1757
rect 2289 1752 2318 1757
rect 2449 1752 2526 1757
rect 2593 1752 2662 1757
rect 3161 1752 3198 1757
rect 3345 1752 3462 1757
rect 3473 1752 3518 1757
rect 3617 1752 3710 1757
rect 1577 1747 1718 1752
rect 3617 1747 3622 1752
rect 361 1742 494 1747
rect 529 1742 670 1747
rect 745 1742 854 1747
rect 865 1742 894 1747
rect 1201 1742 1262 1747
rect 1281 1742 1318 1747
rect 1345 1742 1398 1747
rect 1465 1742 1494 1747
rect 1777 1742 1990 1747
rect 2001 1742 2062 1747
rect 2121 1742 2166 1747
rect 2177 1742 2302 1747
rect 2337 1742 2430 1747
rect 2497 1742 2590 1747
rect 2729 1742 2798 1747
rect 3009 1742 3126 1747
rect 3217 1742 3334 1747
rect 3369 1742 3406 1747
rect 3433 1742 3486 1747
rect 3497 1742 3622 1747
rect 3705 1747 3710 1752
rect 3825 1752 4054 1757
rect 3825 1747 3830 1752
rect 3705 1742 3830 1747
rect 3977 1742 4062 1747
rect 1281 1737 1286 1742
rect 833 1732 886 1737
rect 993 1732 1022 1737
rect 1041 1732 1174 1737
rect 1193 1732 1286 1737
rect 1313 1737 1318 1742
rect 1985 1737 1990 1742
rect 2337 1737 2342 1742
rect 1313 1732 1374 1737
rect 1385 1732 1470 1737
rect 1513 1732 1662 1737
rect 1985 1732 2342 1737
rect 2425 1737 2430 1742
rect 2609 1737 2710 1742
rect 2425 1732 2614 1737
rect 2705 1732 2870 1737
rect 3313 1732 3334 1737
rect 3409 1732 3446 1737
rect 3929 1732 4014 1737
rect 313 1727 494 1732
rect 1041 1727 1046 1732
rect 241 1722 318 1727
rect 489 1722 606 1727
rect 985 1722 1046 1727
rect 1169 1727 1174 1732
rect 1513 1727 1518 1732
rect 1169 1722 1518 1727
rect 1657 1727 1662 1732
rect 1817 1727 1894 1732
rect 3081 1727 3158 1732
rect 3505 1727 3582 1732
rect 4009 1727 4014 1732
rect 4073 1732 4118 1737
rect 4073 1727 4078 1732
rect 1657 1722 1822 1727
rect 1889 1722 2790 1727
rect 2841 1722 2878 1727
rect 3057 1722 3086 1727
rect 3153 1722 3510 1727
rect 3577 1722 3774 1727
rect 3841 1722 3950 1727
rect 4009 1722 4078 1727
rect 137 1712 190 1717
rect 329 1712 374 1717
rect 433 1712 478 1717
rect 705 1712 758 1717
rect 801 1712 838 1717
rect 961 1712 1182 1717
rect 1233 1712 1262 1717
rect 1305 1712 1334 1717
rect 1489 1712 1526 1717
rect 1577 1712 1646 1717
rect 1833 1712 1878 1717
rect 1953 1712 2014 1717
rect 2081 1712 2134 1717
rect 2153 1712 2198 1717
rect 2297 1712 2334 1717
rect 2433 1712 2478 1717
rect 2513 1712 2550 1717
rect 1353 1707 1470 1712
rect 1665 1707 1814 1712
rect 2569 1707 2734 1712
rect 2785 1707 2790 1722
rect 2897 1712 2998 1717
rect 3017 1712 3054 1717
rect 3121 1712 3142 1717
rect 3393 1712 3454 1717
rect 3529 1712 3566 1717
rect 3721 1712 3806 1717
rect 3929 1712 3990 1717
rect 2897 1707 2902 1712
rect 169 1702 246 1707
rect 313 1702 390 1707
rect 425 1702 478 1707
rect 689 1702 718 1707
rect 801 1702 926 1707
rect 1081 1702 1358 1707
rect 1465 1702 1670 1707
rect 1809 1702 2574 1707
rect 2729 1702 2758 1707
rect 2785 1702 2902 1707
rect 2993 1707 2998 1712
rect 2993 1702 3446 1707
rect 3481 1702 3526 1707
rect 713 1697 806 1702
rect 377 1692 430 1697
rect 497 1692 670 1697
rect 961 1692 1006 1697
rect 1153 1692 1198 1697
rect 1209 1692 1246 1697
rect 1265 1692 1310 1697
rect 1321 1692 1350 1697
rect 1409 1692 1814 1697
rect 1969 1692 2022 1697
rect 2041 1692 2982 1697
rect 3537 1692 3622 1697
rect 265 1682 446 1687
rect 497 1677 502 1692
rect 385 1672 502 1677
rect 665 1677 670 1692
rect 825 1687 942 1692
rect 1025 1687 1134 1692
rect 1833 1687 1950 1692
rect 2977 1687 3142 1692
rect 3313 1687 3542 1692
rect 721 1682 774 1687
rect 801 1682 830 1687
rect 937 1682 1030 1687
rect 1129 1682 1838 1687
rect 1945 1682 2230 1687
rect 2473 1682 2694 1687
rect 2809 1682 2838 1687
rect 3137 1682 3318 1687
rect 3649 1682 3870 1687
rect 2225 1677 2478 1682
rect 2689 1677 2814 1682
rect 665 1672 822 1677
rect 881 1672 1422 1677
rect 1513 1672 1598 1677
rect 1761 1672 1998 1677
rect 2057 1672 2086 1677
rect 2601 1672 2670 1677
rect 2993 1672 3118 1677
rect 3337 1672 3502 1677
rect 1417 1667 1518 1672
rect 1593 1667 1766 1672
rect 2105 1667 2206 1672
rect 2497 1667 2582 1672
rect 449 1662 542 1667
rect 585 1662 654 1667
rect 713 1662 982 1667
rect 1081 1662 1398 1667
rect 1537 1662 1574 1667
rect 1785 1662 2110 1667
rect 2201 1662 2502 1667
rect 2577 1662 2870 1667
rect 649 1657 718 1662
rect 2865 1657 2870 1662
rect 3649 1657 3654 1682
rect 3865 1667 3870 1682
rect 3713 1662 3782 1667
rect 3865 1662 4078 1667
rect 3713 1657 3718 1662
rect 209 1652 366 1657
rect 505 1652 534 1657
rect 737 1652 1350 1657
rect 1409 1652 1518 1657
rect 1681 1652 1726 1657
rect 1889 1652 2190 1657
rect 2513 1652 2566 1657
rect 2641 1652 2718 1657
rect 2865 1652 2974 1657
rect 3009 1652 3062 1657
rect 3081 1652 3158 1657
rect 3273 1652 3382 1657
rect 3433 1652 3654 1657
rect 3673 1652 3718 1657
rect 3777 1657 3782 1662
rect 3777 1652 3854 1657
rect 209 1637 214 1652
rect 185 1632 214 1637
rect 361 1637 366 1652
rect 1345 1647 1414 1652
rect 2209 1647 2310 1652
rect 2737 1647 2830 1652
rect 2969 1647 2974 1652
rect 3081 1647 3086 1652
rect 417 1642 494 1647
rect 529 1642 630 1647
rect 817 1642 974 1647
rect 529 1637 534 1642
rect 969 1637 974 1642
rect 1057 1642 1086 1647
rect 1105 1642 1150 1647
rect 1273 1642 1326 1647
rect 1497 1642 1534 1647
rect 1545 1642 1630 1647
rect 1705 1642 2214 1647
rect 2305 1642 2742 1647
rect 2825 1642 2854 1647
rect 2969 1642 3086 1647
rect 3153 1647 3158 1652
rect 3153 1642 3270 1647
rect 3729 1642 3766 1647
rect 1057 1637 1062 1642
rect 361 1632 534 1637
rect 545 1632 726 1637
rect 545 1627 550 1632
rect 721 1627 726 1632
rect 785 1632 886 1637
rect 969 1632 1062 1637
rect 1121 1632 1334 1637
rect 1545 1632 1758 1637
rect 1825 1632 1878 1637
rect 2001 1632 2070 1637
rect 2097 1632 2294 1637
rect 2537 1632 2582 1637
rect 2633 1632 2686 1637
rect 2705 1632 2750 1637
rect 2801 1632 2838 1637
rect 2857 1632 2942 1637
rect 2953 1632 3142 1637
rect 3209 1632 3246 1637
rect 3297 1632 3406 1637
rect 3465 1632 3526 1637
rect 3697 1632 3726 1637
rect 3809 1632 3878 1637
rect 3961 1632 3998 1637
rect 785 1627 790 1632
rect 113 1622 174 1627
rect 281 1622 326 1627
rect 441 1622 550 1627
rect 569 1622 614 1627
rect 721 1622 790 1627
rect 905 1622 950 1627
rect 1137 1617 1142 1627
rect 1161 1622 1238 1627
rect 1249 1622 1558 1627
rect 1817 1622 1942 1627
rect 1977 1622 2086 1627
rect 209 1597 214 1617
rect 337 1612 414 1617
rect 641 1612 670 1617
rect 1009 1612 1086 1617
rect 1105 1612 1182 1617
rect 641 1607 646 1612
rect 1009 1607 1014 1612
rect 225 1602 374 1607
rect 609 1602 646 1607
rect 809 1602 830 1607
rect 881 1602 1014 1607
rect 1081 1607 1086 1612
rect 1249 1607 1254 1622
rect 1601 1617 1710 1622
rect 2081 1617 2086 1622
rect 2217 1622 2246 1627
rect 2297 1622 2406 1627
rect 3993 1622 4150 1627
rect 2217 1617 2222 1622
rect 1313 1612 1358 1617
rect 1521 1612 1606 1617
rect 1705 1612 1734 1617
rect 1937 1612 2030 1617
rect 2081 1612 2222 1617
rect 1313 1607 1318 1612
rect 1377 1607 1502 1612
rect 2401 1607 2406 1622
rect 2889 1617 3230 1622
rect 3657 1617 3742 1622
rect 2417 1612 2502 1617
rect 2545 1612 2582 1617
rect 2793 1612 2894 1617
rect 3225 1612 3254 1617
rect 3265 1612 3294 1617
rect 3633 1612 3662 1617
rect 3737 1612 3918 1617
rect 1081 1602 1254 1607
rect 1273 1602 1318 1607
rect 1337 1602 1382 1607
rect 1497 1602 1526 1607
rect 1593 1602 1670 1607
rect 1889 1602 1982 1607
rect 1993 1602 2062 1607
rect 2345 1602 2390 1607
rect 2401 1602 2710 1607
rect 2905 1602 3078 1607
rect 3089 1602 3222 1607
rect 3281 1602 3374 1607
rect 3697 1602 3726 1607
rect 2705 1597 2710 1602
rect 185 1592 214 1597
rect 289 1592 350 1597
rect 433 1592 582 1597
rect 601 1592 686 1597
rect 801 1592 942 1597
rect 1065 1592 1166 1597
rect 1289 1592 1382 1597
rect 1393 1592 1582 1597
rect 1657 1592 1782 1597
rect 2001 1592 2030 1597
rect 2081 1592 2182 1597
rect 2201 1592 2302 1597
rect 2377 1592 2470 1597
rect 2561 1592 2694 1597
rect 2705 1592 2798 1597
rect 3009 1592 3038 1597
rect 289 1587 294 1592
rect 433 1587 438 1592
rect 161 1582 294 1587
rect 361 1582 438 1587
rect 577 1587 582 1592
rect 2081 1587 2086 1592
rect 577 1582 710 1587
rect 1025 1582 1054 1587
rect 729 1577 830 1582
rect 1049 1577 1054 1582
rect 1177 1582 2086 1587
rect 2177 1587 2182 1592
rect 3033 1587 3038 1592
rect 3097 1592 3150 1597
rect 3201 1592 3238 1597
rect 3305 1592 3366 1597
rect 3401 1592 3510 1597
rect 3665 1592 3726 1597
rect 3769 1592 3838 1597
rect 3985 1592 4078 1597
rect 3097 1587 3102 1592
rect 3769 1587 3774 1592
rect 2177 1582 2470 1587
rect 2609 1582 2638 1587
rect 3033 1582 3102 1587
rect 3249 1582 3390 1587
rect 3705 1582 3774 1587
rect 3833 1587 3838 1592
rect 3833 1582 4022 1587
rect 1177 1577 1182 1582
rect 193 1572 262 1577
rect 401 1572 734 1577
rect 825 1572 886 1577
rect 905 1572 926 1577
rect 993 1572 1014 1577
rect 1049 1572 1182 1577
rect 1265 1572 1518 1577
rect 1529 1572 1638 1577
rect 1809 1572 1886 1577
rect 2217 1572 2238 1577
rect 2265 1572 2310 1577
rect 2329 1572 2382 1577
rect 2753 1572 2886 1577
rect 3121 1572 3182 1577
rect 3193 1572 3294 1577
rect 3609 1572 3710 1577
rect 3785 1572 3846 1577
rect 3921 1572 4054 1577
rect 1657 1567 1790 1572
rect 2025 1567 2198 1572
rect 193 1562 222 1567
rect 513 1562 646 1567
rect 641 1557 646 1562
rect 745 1562 814 1567
rect 745 1557 750 1562
rect 417 1552 454 1557
rect 521 1552 622 1557
rect 641 1552 750 1557
rect 809 1557 814 1562
rect 897 1562 926 1567
rect 1201 1562 1358 1567
rect 1401 1562 1662 1567
rect 1785 1562 2030 1567
rect 2193 1562 2278 1567
rect 2369 1562 2398 1567
rect 2673 1562 2790 1567
rect 2817 1562 2982 1567
rect 3185 1562 3254 1567
rect 3305 1562 3470 1567
rect 3585 1562 3646 1567
rect 3793 1562 3822 1567
rect 3945 1562 4110 1567
rect 897 1557 902 1562
rect 2273 1557 2374 1562
rect 2817 1557 2822 1562
rect 809 1552 902 1557
rect 1297 1552 1318 1557
rect 1537 1552 1566 1557
rect 1577 1552 1878 1557
rect 2041 1552 2254 1557
rect 2737 1552 2822 1557
rect 2841 1552 2870 1557
rect 3177 1552 3342 1557
rect 1337 1547 1422 1552
rect 3337 1547 3342 1552
rect 3409 1552 3438 1557
rect 3521 1552 3550 1557
rect 3777 1552 3806 1557
rect 3945 1552 3998 1557
rect 3409 1547 3414 1552
rect 161 1542 374 1547
rect 385 1542 542 1547
rect 561 1542 590 1547
rect 769 1542 790 1547
rect 929 1542 1134 1547
rect 1217 1542 1342 1547
rect 1417 1542 1966 1547
rect 2289 1542 2326 1547
rect 2345 1542 2454 1547
rect 2473 1542 2526 1547
rect 2545 1542 2654 1547
rect 2689 1542 2750 1547
rect 2865 1542 2942 1547
rect 3089 1542 3158 1547
rect 3201 1542 3286 1547
rect 3337 1542 3414 1547
rect 3537 1542 3614 1547
rect 3689 1542 3774 1547
rect 3817 1542 3926 1547
rect 4001 1542 4062 1547
rect 369 1537 374 1542
rect 113 1532 150 1537
rect 145 1527 150 1532
rect 209 1532 262 1537
rect 369 1532 398 1537
rect 529 1532 566 1537
rect 641 1532 734 1537
rect 209 1527 214 1532
rect 393 1527 534 1532
rect 641 1527 646 1532
rect 145 1522 214 1527
rect 553 1522 646 1527
rect 729 1527 734 1532
rect 729 1522 758 1527
rect 769 1517 774 1542
rect 2137 1537 2270 1542
rect 2345 1537 2350 1542
rect 833 1532 862 1537
rect 1313 1532 1406 1537
rect 1497 1532 1542 1537
rect 1801 1532 1822 1537
rect 1985 1532 2094 1537
rect 2113 1532 2142 1537
rect 2265 1532 2350 1537
rect 2449 1537 2454 1542
rect 2545 1537 2550 1542
rect 2449 1532 2550 1537
rect 2649 1537 2654 1542
rect 2649 1532 3046 1537
rect 3241 1532 3294 1537
rect 3489 1532 3630 1537
rect 3881 1532 3942 1537
rect 1561 1527 1782 1532
rect 1841 1527 1990 1532
rect 2089 1527 2094 1532
rect 953 1522 1038 1527
rect 1105 1522 1126 1527
rect 1145 1522 1294 1527
rect 953 1517 958 1522
rect 233 1512 278 1517
rect 353 1512 398 1517
rect 521 1512 558 1517
rect 569 1512 598 1517
rect 633 1512 774 1517
rect 785 1512 822 1517
rect 857 1512 958 1517
rect 1033 1517 1038 1522
rect 1145 1517 1150 1522
rect 1033 1512 1150 1517
rect 1289 1517 1294 1522
rect 1345 1522 1566 1527
rect 1777 1522 1846 1527
rect 2089 1522 2438 1527
rect 2537 1522 2670 1527
rect 2793 1522 2854 1527
rect 2913 1522 3222 1527
rect 3329 1522 3438 1527
rect 3793 1522 3822 1527
rect 1345 1517 1350 1522
rect 2433 1517 2542 1522
rect 3969 1517 3974 1537
rect 1289 1512 1350 1517
rect 1433 1512 2182 1517
rect 2249 1512 2406 1517
rect 2561 1512 2622 1517
rect 2697 1512 3062 1517
rect 3081 1512 3126 1517
rect 3153 1512 3198 1517
rect 3353 1512 3406 1517
rect 3793 1512 3838 1517
rect 3969 1512 3990 1517
rect 4009 1512 4134 1517
rect 3985 1507 3990 1512
rect 249 1502 414 1507
rect 513 1502 542 1507
rect 553 1502 590 1507
rect 689 1502 830 1507
rect 841 1502 886 1507
rect 969 1502 1022 1507
rect 1089 1502 1126 1507
rect 1161 1502 1278 1507
rect 1345 1502 1406 1507
rect 1449 1502 1598 1507
rect 1617 1502 1678 1507
rect 1745 1502 2166 1507
rect 2185 1502 2214 1507
rect 2225 1502 2574 1507
rect 2857 1502 3022 1507
rect 3297 1502 3470 1507
rect 3825 1502 3878 1507
rect 3985 1502 4078 1507
rect 1273 1497 1350 1502
rect 561 1492 606 1497
rect 641 1492 686 1497
rect 753 1492 1062 1497
rect 1721 1492 2150 1497
rect 2161 1492 2286 1497
rect 2361 1492 2390 1497
rect 2713 1492 2918 1497
rect 1537 1487 1630 1492
rect 2145 1487 2150 1492
rect 2913 1487 2918 1492
rect 3001 1492 3030 1497
rect 3177 1492 3462 1497
rect 3841 1492 3958 1497
rect 3001 1487 3006 1492
rect 537 1482 742 1487
rect 857 1482 982 1487
rect 993 1482 1046 1487
rect 1105 1482 1238 1487
rect 1257 1482 1286 1487
rect 1305 1482 1382 1487
rect 1401 1482 1494 1487
rect 1513 1482 1542 1487
rect 1625 1482 1694 1487
rect 1105 1477 1110 1482
rect 433 1472 518 1477
rect 601 1472 1110 1477
rect 1233 1477 1238 1482
rect 1401 1477 1406 1482
rect 1233 1472 1406 1477
rect 1489 1477 1494 1482
rect 1689 1477 1694 1482
rect 1865 1482 1902 1487
rect 2145 1482 2230 1487
rect 2849 1482 2894 1487
rect 2913 1482 3006 1487
rect 3329 1482 3382 1487
rect 3473 1482 3558 1487
rect 3665 1482 3742 1487
rect 1865 1477 1870 1482
rect 3665 1477 3670 1482
rect 1489 1472 1614 1477
rect 1689 1472 1870 1477
rect 1889 1472 1998 1477
rect 2105 1472 2190 1477
rect 2409 1472 2694 1477
rect 3145 1472 3670 1477
rect 3737 1477 3742 1482
rect 3737 1472 3918 1477
rect 433 1467 438 1472
rect 409 1462 438 1467
rect 513 1467 518 1472
rect 2409 1467 2414 1472
rect 513 1462 694 1467
rect 705 1462 742 1467
rect 753 1462 798 1467
rect 841 1462 878 1467
rect 953 1462 990 1467
rect 1009 1462 1054 1467
rect 1121 1462 1238 1467
rect 1417 1462 1638 1467
rect 2177 1462 2414 1467
rect 2689 1467 2694 1472
rect 2689 1462 2798 1467
rect 2841 1462 3126 1467
rect 3649 1462 3726 1467
rect 689 1447 694 1462
rect 1233 1457 1422 1462
rect 2433 1457 2518 1462
rect 2841 1457 2846 1462
rect 793 1452 1110 1457
rect 1513 1452 1566 1457
rect 1633 1452 1670 1457
rect 2409 1452 2438 1457
rect 2513 1452 2678 1457
rect 2817 1452 2846 1457
rect 3121 1457 3126 1462
rect 3361 1457 3494 1462
rect 3721 1457 3726 1462
rect 3849 1462 3942 1467
rect 3849 1457 3854 1462
rect 3121 1452 3230 1457
rect 3337 1452 3366 1457
rect 3489 1452 3518 1457
rect 3721 1452 3854 1457
rect 793 1447 798 1452
rect 1105 1447 1214 1452
rect 1513 1447 1518 1452
rect 2241 1447 2390 1452
rect 2673 1447 2822 1452
rect 249 1442 390 1447
rect 417 1442 438 1447
rect 473 1442 502 1447
rect 689 1442 798 1447
rect 833 1442 1086 1447
rect 1209 1442 1518 1447
rect 1553 1442 1686 1447
rect 1769 1442 2246 1447
rect 2385 1442 2502 1447
rect 2857 1442 2950 1447
rect 3385 1442 3454 1447
rect 3481 1442 3518 1447
rect 3537 1442 3606 1447
rect 3873 1442 3894 1447
rect 3913 1442 3974 1447
rect 249 1437 254 1442
rect 209 1432 254 1437
rect 385 1437 390 1442
rect 3161 1437 3278 1442
rect 3537 1437 3542 1442
rect 385 1432 534 1437
rect 817 1432 854 1437
rect 937 1432 982 1437
rect 1041 1432 1094 1437
rect 1145 1432 1190 1437
rect 1561 1432 1590 1437
rect 2257 1432 2406 1437
rect 2705 1432 2742 1437
rect 2753 1432 2814 1437
rect 2865 1432 3166 1437
rect 3273 1432 3302 1437
rect 3417 1432 3542 1437
rect 3601 1437 3606 1442
rect 3601 1432 3670 1437
rect 3681 1432 3750 1437
rect 3817 1432 3870 1437
rect 3889 1432 4014 1437
rect 129 1422 166 1427
rect 313 1422 358 1427
rect 369 1422 462 1427
rect 561 1422 590 1427
rect 681 1422 734 1427
rect 905 1422 950 1427
rect 1017 1422 1126 1427
rect 1185 1422 1550 1427
rect 1577 1422 1622 1427
rect 1673 1422 1766 1427
rect 1873 1422 1918 1427
rect 1937 1422 2030 1427
rect 369 1417 374 1422
rect 1185 1417 1190 1422
rect 1937 1417 1942 1422
rect 265 1412 374 1417
rect 385 1412 430 1417
rect 649 1412 678 1417
rect 897 1412 958 1417
rect 977 1412 1046 1417
rect 1065 1412 1094 1417
rect 1145 1412 1190 1417
rect 1665 1412 1694 1417
rect 1777 1412 1942 1417
rect 2025 1417 2030 1422
rect 2065 1422 2150 1427
rect 2169 1422 2198 1427
rect 2209 1422 2358 1427
rect 2425 1422 2486 1427
rect 2521 1422 2678 1427
rect 2025 1412 2054 1417
rect 249 1402 366 1407
rect 673 1402 678 1412
rect 977 1407 982 1412
rect 1089 1407 1094 1412
rect 1689 1407 1782 1412
rect 2065 1407 2070 1422
rect 2145 1417 2150 1422
rect 2521 1417 2526 1422
rect 2145 1412 2526 1417
rect 2673 1407 2678 1422
rect 2729 1417 2734 1427
rect 2889 1422 3022 1427
rect 3113 1422 3150 1427
rect 3177 1422 3238 1427
rect 3529 1422 3590 1427
rect 3657 1422 3702 1427
rect 3713 1422 3934 1427
rect 3257 1417 3510 1422
rect 2729 1412 2750 1417
rect 2897 1412 2950 1417
rect 3033 1412 3102 1417
rect 3153 1412 3262 1417
rect 3505 1412 3566 1417
rect 3577 1412 3646 1417
rect 3729 1412 3790 1417
rect 4017 1412 4054 1417
rect 3729 1407 3734 1412
rect 793 1402 982 1407
rect 1049 1402 1094 1407
rect 1345 1402 1390 1407
rect 1881 1402 2070 1407
rect 2089 1402 2142 1407
rect 2241 1402 2526 1407
rect 2673 1402 3678 1407
rect 3729 1402 3758 1407
rect 3817 1402 3862 1407
rect 3953 1402 4030 1407
rect 345 1392 494 1397
rect 617 1392 670 1397
rect 713 1392 806 1397
rect 961 1392 1038 1397
rect 1209 1392 1294 1397
rect 1377 1392 1470 1397
rect 1721 1392 1758 1397
rect 1809 1392 1878 1397
rect 1985 1392 2070 1397
rect 2201 1392 2286 1397
rect 2361 1392 2566 1397
rect 2609 1392 2662 1397
rect 2673 1392 2742 1397
rect 2753 1392 2790 1397
rect 2881 1392 2942 1397
rect 3033 1392 3070 1397
rect 3193 1392 3374 1397
rect 3481 1392 3574 1397
rect 3737 1392 3774 1397
rect 3889 1392 3982 1397
rect 417 1382 462 1387
rect 593 1382 790 1387
rect 921 1382 958 1387
rect 1161 1382 1262 1387
rect 1273 1382 1318 1387
rect 1425 1382 1510 1387
rect 1833 1382 1894 1387
rect 2041 1382 3222 1387
rect 3305 1382 3334 1387
rect 3457 1382 3486 1387
rect 3513 1382 3534 1387
rect 3561 1382 3606 1387
rect 3681 1382 4038 1387
rect 3217 1377 3310 1382
rect 3681 1377 3686 1382
rect 513 1372 550 1377
rect 657 1372 686 1377
rect 705 1372 774 1377
rect 793 1372 814 1377
rect 1305 1372 1550 1377
rect 1913 1372 2014 1377
rect 2033 1372 2062 1377
rect 2145 1372 2614 1377
rect 2625 1372 2678 1377
rect 2745 1372 2774 1377
rect 2785 1372 2806 1377
rect 2833 1372 2902 1377
rect 3049 1372 3198 1377
rect 3345 1372 3406 1377
rect 3537 1372 3574 1377
rect 3593 1372 3686 1377
rect 3737 1372 3766 1377
rect 3785 1372 3862 1377
rect 3873 1372 3902 1377
rect 3961 1372 3982 1377
rect 1913 1367 1918 1372
rect 361 1362 462 1367
rect 497 1362 534 1367
rect 665 1362 862 1367
rect 977 1362 1086 1367
rect 1153 1362 1206 1367
rect 1217 1362 1254 1367
rect 1385 1362 1446 1367
rect 1569 1362 1806 1367
rect 1825 1362 1918 1367
rect 2009 1367 2014 1372
rect 2921 1367 3030 1372
rect 2009 1362 2102 1367
rect 2121 1362 2414 1367
rect 2473 1362 2494 1367
rect 2529 1362 2926 1367
rect 3025 1362 3622 1367
rect 3721 1362 4086 1367
rect 977 1357 982 1362
rect 361 1352 646 1357
rect 681 1352 726 1357
rect 737 1352 782 1357
rect 945 1352 982 1357
rect 1081 1357 1086 1362
rect 1569 1357 1574 1362
rect 1081 1352 1110 1357
rect 1281 1352 1366 1357
rect 1521 1352 1574 1357
rect 1801 1357 1806 1362
rect 3617 1357 3726 1362
rect 1801 1352 1878 1357
rect 1897 1352 2086 1357
rect 2169 1352 2398 1357
rect 2489 1352 2518 1357
rect 2553 1352 2582 1357
rect 2617 1352 2670 1357
rect 2793 1352 2886 1357
rect 2905 1352 3054 1357
rect 3081 1352 3238 1357
rect 3537 1352 3598 1357
rect 3745 1352 3870 1357
rect 1281 1347 1286 1352
rect 337 1342 382 1347
rect 401 1342 542 1347
rect 609 1342 838 1347
rect 937 1342 1014 1347
rect 1025 1342 1134 1347
rect 1257 1342 1286 1347
rect 1361 1347 1366 1352
rect 2393 1347 2494 1352
rect 3337 1347 3438 1352
rect 3537 1347 3542 1352
rect 3865 1347 3870 1352
rect 3969 1352 3998 1357
rect 3969 1347 3974 1352
rect 1361 1342 1390 1347
rect 1649 1342 1750 1347
rect 1849 1342 1990 1347
rect 2049 1342 2254 1347
rect 2337 1342 2366 1347
rect 2545 1342 2606 1347
rect 2641 1342 2694 1347
rect 2721 1342 2790 1347
rect 2865 1342 2894 1347
rect 2945 1342 2966 1347
rect 3041 1342 3134 1347
rect 3145 1342 3190 1347
rect 3217 1342 3342 1347
rect 3433 1342 3542 1347
rect 3553 1342 3630 1347
rect 3729 1342 3758 1347
rect 3777 1342 3846 1347
rect 3865 1342 3974 1347
rect 4017 1342 4062 1347
rect 401 1337 406 1342
rect 2249 1337 2342 1342
rect 297 1332 406 1337
rect 449 1332 494 1337
rect 513 1332 534 1337
rect 721 1332 750 1337
rect 785 1332 1022 1337
rect 1065 1332 1318 1337
rect 1329 1332 1414 1337
rect 1505 1332 2078 1337
rect 2377 1332 2534 1337
rect 2601 1332 2822 1337
rect 2873 1332 2918 1337
rect 2953 1332 2990 1337
rect 3177 1332 3246 1337
rect 3353 1332 3414 1337
rect 3633 1332 3678 1337
rect 4009 1332 4102 1337
rect 513 1327 518 1332
rect 2073 1327 2214 1332
rect 2377 1327 2382 1332
rect 2529 1327 2606 1332
rect 465 1322 502 1327
rect 513 1322 542 1327
rect 921 1322 974 1327
rect 993 1322 1046 1327
rect 1481 1322 1542 1327
rect 1729 1322 2014 1327
rect 2025 1322 2054 1327
rect 2209 1322 2382 1327
rect 2625 1322 2678 1327
rect 2841 1322 2870 1327
rect 3529 1322 3574 1327
rect 3713 1322 3782 1327
rect 3929 1322 4118 1327
rect 129 1312 174 1317
rect 249 1312 318 1317
rect 337 1312 454 1317
rect 473 1312 534 1317
rect 641 1312 750 1317
rect 793 1312 814 1317
rect 1313 1312 1502 1317
rect 1585 1312 1822 1317
rect 1833 1312 1862 1317
rect 1881 1312 1934 1317
rect 2081 1312 2150 1317
rect 2161 1312 2190 1317
rect 2465 1312 2502 1317
rect 2545 1312 2654 1317
rect 249 1307 254 1312
rect 161 1302 254 1307
rect 313 1307 318 1312
rect 2145 1307 2150 1312
rect 313 1302 630 1307
rect 873 1302 934 1307
rect 993 1302 1030 1307
rect 1769 1302 2078 1307
rect 2145 1302 2222 1307
rect 2241 1302 2446 1307
rect 2529 1302 2574 1307
rect 2625 1302 2630 1312
rect 2673 1307 2678 1322
rect 2913 1317 3006 1322
rect 2705 1312 2790 1317
rect 2889 1312 2918 1317
rect 3001 1312 3222 1317
rect 3329 1312 3382 1317
rect 3489 1312 3566 1317
rect 3593 1312 3694 1317
rect 3785 1312 3918 1317
rect 4017 1312 4070 1317
rect 4113 1312 4118 1322
rect 3593 1307 3598 1312
rect 2673 1302 2726 1307
rect 2945 1302 2990 1307
rect 3473 1302 3526 1307
rect 3545 1302 3598 1307
rect 3689 1307 3694 1312
rect 3689 1302 3750 1307
rect 3769 1302 3822 1307
rect 3905 1302 3958 1307
rect 265 1292 718 1297
rect 1025 1292 1198 1297
rect 1217 1292 1382 1297
rect 1545 1292 1638 1297
rect 1817 1292 2038 1297
rect 2073 1292 2174 1297
rect 1217 1287 1222 1292
rect 385 1282 478 1287
rect 729 1282 878 1287
rect 993 1282 1054 1287
rect 1137 1282 1222 1287
rect 1377 1287 1382 1292
rect 1697 1287 1798 1292
rect 2241 1287 2246 1302
rect 2441 1292 2446 1302
rect 2609 1292 2846 1297
rect 3497 1292 3518 1297
rect 3537 1292 3742 1297
rect 4033 1292 4070 1297
rect 2441 1287 2590 1292
rect 1377 1282 1406 1287
rect 1425 1282 1526 1287
rect 1673 1282 1702 1287
rect 1793 1282 2246 1287
rect 2265 1282 2422 1287
rect 2585 1282 2742 1287
rect 2857 1282 3158 1287
rect 3753 1282 3814 1287
rect 473 1277 478 1282
rect 633 1277 734 1282
rect 1241 1277 1358 1282
rect 1425 1277 1430 1282
rect 1521 1277 1654 1282
rect 2265 1277 2270 1282
rect 473 1272 638 1277
rect 1169 1272 1246 1277
rect 1353 1272 1430 1277
rect 1649 1272 2270 1277
rect 2417 1277 2422 1282
rect 2737 1277 2862 1282
rect 2417 1272 2718 1277
rect 3873 1272 3958 1277
rect 1049 1267 1174 1272
rect 3873 1267 3878 1272
rect 297 1262 366 1267
rect 297 1257 302 1262
rect 169 1252 302 1257
rect 361 1257 366 1262
rect 377 1262 454 1267
rect 657 1262 686 1267
rect 377 1257 382 1262
rect 361 1252 382 1257
rect 449 1257 454 1262
rect 681 1257 686 1262
rect 849 1262 1054 1267
rect 1185 1262 1342 1267
rect 1433 1262 2246 1267
rect 2265 1262 3014 1267
rect 3137 1262 3214 1267
rect 3233 1262 3270 1267
rect 3801 1262 3878 1267
rect 3953 1267 3958 1272
rect 3953 1262 3982 1267
rect 849 1257 854 1262
rect 1337 1257 1438 1262
rect 2241 1257 2246 1262
rect 3137 1257 3142 1262
rect 449 1252 582 1257
rect 681 1252 854 1257
rect 873 1252 902 1257
rect 897 1247 902 1252
rect 1065 1252 1318 1257
rect 1457 1252 2174 1257
rect 2241 1252 2318 1257
rect 2393 1252 2446 1257
rect 2521 1252 2694 1257
rect 3113 1252 3142 1257
rect 3209 1257 3214 1262
rect 3209 1252 3302 1257
rect 3417 1252 3518 1257
rect 3889 1252 3982 1257
rect 4009 1252 4078 1257
rect 1065 1247 1070 1252
rect 97 1242 246 1247
rect 393 1242 438 1247
rect 897 1242 1070 1247
rect 1089 1242 1118 1247
rect 1201 1242 1230 1247
rect 265 1237 366 1242
rect 1113 1237 1206 1242
rect 1313 1237 1318 1252
rect 2769 1247 2926 1252
rect 1401 1242 1470 1247
rect 1481 1242 1918 1247
rect 2065 1242 2134 1247
rect 2193 1242 2270 1247
rect 2649 1242 2774 1247
rect 2921 1242 3430 1247
rect 1913 1237 2070 1242
rect 209 1232 270 1237
rect 361 1232 390 1237
rect 1257 1232 1302 1237
rect 1313 1232 1702 1237
rect 1801 1232 1830 1237
rect 1849 1232 1894 1237
rect 2089 1232 2230 1237
rect 2369 1232 2438 1237
rect 2593 1232 2646 1237
rect 2785 1232 2910 1237
rect 3137 1232 3998 1237
rect 1697 1227 1806 1232
rect 2905 1227 3142 1232
rect 89 1222 142 1227
rect 185 1222 230 1227
rect 281 1222 326 1227
rect 401 1222 446 1227
rect 601 1222 646 1227
rect 681 1222 702 1227
rect 825 1222 870 1227
rect 985 1222 1078 1227
rect 1129 1222 1206 1227
rect 1241 1222 1430 1227
rect 1449 1222 1478 1227
rect 1473 1217 1478 1222
rect 1553 1222 1678 1227
rect 1969 1222 2062 1227
rect 2081 1222 2158 1227
rect 2209 1222 2270 1227
rect 2337 1222 2366 1227
rect 2777 1222 2886 1227
rect 3209 1222 3358 1227
rect 3401 1222 3430 1227
rect 1553 1217 1558 1222
rect 1969 1217 1974 1222
rect 273 1212 302 1217
rect 385 1212 422 1217
rect 577 1212 622 1217
rect 849 1212 934 1217
rect 1065 1212 1102 1217
rect 1193 1212 1238 1217
rect 1273 1212 1334 1217
rect 1473 1212 1558 1217
rect 1577 1212 1670 1217
rect 1697 1212 1766 1217
rect 1945 1212 1974 1217
rect 2057 1217 2062 1222
rect 3425 1217 3430 1222
rect 3513 1222 3542 1227
rect 3569 1222 3590 1227
rect 3513 1217 3518 1222
rect 2057 1212 2134 1217
rect 2457 1212 2574 1217
rect 2153 1207 2246 1212
rect 2457 1207 2462 1212
rect 137 1202 350 1207
rect 569 1202 606 1207
rect 841 1202 910 1207
rect 1145 1202 1206 1207
rect 1369 1202 1406 1207
rect 1617 1202 1694 1207
rect 1857 1202 2158 1207
rect 2241 1202 2462 1207
rect 2569 1207 2574 1212
rect 2681 1212 2758 1217
rect 2865 1212 3006 1217
rect 3073 1212 3142 1217
rect 3257 1212 3310 1217
rect 3425 1212 3518 1217
rect 2681 1207 2686 1212
rect 2753 1207 2846 1212
rect 3073 1207 3078 1212
rect 2569 1202 2686 1207
rect 2841 1202 2910 1207
rect 3009 1202 3078 1207
rect 169 1192 222 1197
rect 257 1192 550 1197
rect 617 1192 782 1197
rect 857 1192 950 1197
rect 977 1192 1014 1197
rect 1073 1192 1102 1197
rect 1129 1192 1222 1197
rect 1321 1192 1446 1197
rect 1529 1192 1614 1197
rect 1689 1192 1726 1197
rect 1745 1192 1838 1197
rect 1857 1192 1862 1202
rect 3137 1197 3142 1212
rect 3209 1202 3286 1207
rect 3681 1202 3686 1227
rect 3697 1202 3702 1227
rect 3729 1222 3758 1227
rect 3753 1217 3758 1222
rect 3841 1222 3870 1227
rect 3977 1222 4030 1227
rect 3841 1217 3846 1222
rect 3753 1212 3846 1217
rect 3881 1212 3926 1217
rect 3977 1202 4014 1207
rect 1873 1192 1950 1197
rect 2113 1192 2166 1197
rect 2193 1192 2230 1197
rect 2433 1192 2582 1197
rect 2697 1192 2798 1197
rect 2809 1192 2838 1197
rect 1745 1187 1750 1192
rect 297 1182 390 1187
rect 417 1182 510 1187
rect 529 1182 686 1187
rect 681 1177 686 1182
rect 793 1182 894 1187
rect 977 1182 998 1187
rect 1169 1182 1286 1187
rect 1401 1182 1750 1187
rect 1833 1187 1838 1192
rect 2833 1187 2838 1192
rect 2921 1192 2998 1197
rect 2921 1187 2926 1192
rect 1833 1182 2062 1187
rect 2145 1182 2182 1187
rect 2249 1182 2350 1187
rect 2369 1182 2430 1187
rect 2441 1182 2470 1187
rect 2529 1182 2574 1187
rect 2833 1182 2926 1187
rect 2993 1187 2998 1192
rect 3089 1192 3118 1197
rect 3137 1192 3190 1197
rect 3233 1192 3278 1197
rect 3393 1192 3454 1197
rect 3473 1192 3558 1197
rect 3737 1192 3798 1197
rect 3929 1192 4022 1197
rect 3089 1187 3094 1192
rect 3473 1187 3478 1192
rect 2993 1182 3094 1187
rect 3113 1182 3478 1187
rect 3553 1187 3558 1192
rect 3553 1182 3870 1187
rect 3913 1182 4038 1187
rect 793 1177 798 1182
rect 2249 1177 2254 1182
rect 513 1172 550 1177
rect 633 1172 662 1177
rect 681 1172 798 1177
rect 1225 1172 1390 1177
rect 1465 1172 2254 1177
rect 2345 1177 2350 1182
rect 2345 1172 2782 1177
rect 3121 1172 3158 1177
rect 3225 1172 3366 1177
rect 3425 1172 3750 1177
rect 3769 1172 4054 1177
rect 1385 1167 1470 1172
rect 129 1162 182 1167
rect 553 1162 630 1167
rect 1281 1162 1326 1167
rect 1529 1162 1822 1167
rect 1897 1162 1934 1167
rect 2129 1162 2438 1167
rect 2801 1162 2958 1167
rect 2977 1162 2998 1167
rect 3169 1162 3198 1167
rect 3497 1162 3550 1167
rect 3561 1162 3590 1167
rect 3601 1162 3710 1167
rect 3753 1162 3790 1167
rect 4009 1162 4110 1167
rect 2457 1157 2686 1162
rect 2801 1157 2806 1162
rect 81 1152 134 1157
rect 361 1152 406 1157
rect 553 1152 598 1157
rect 713 1152 822 1157
rect 873 1152 894 1157
rect 913 1152 1038 1157
rect 1329 1152 1446 1157
rect 1489 1152 1830 1157
rect 129 1147 134 1152
rect 97 1142 118 1147
rect 129 1142 182 1147
rect 273 1142 390 1147
rect 113 1112 118 1142
rect 401 1137 406 1152
rect 913 1147 918 1152
rect 593 1142 702 1147
rect 697 1137 702 1142
rect 809 1142 918 1147
rect 1033 1147 1038 1152
rect 1825 1147 1830 1152
rect 1945 1152 2118 1157
rect 2249 1152 2462 1157
rect 2681 1152 2806 1157
rect 2953 1157 2958 1162
rect 3281 1157 3350 1162
rect 2953 1152 3286 1157
rect 3345 1152 3494 1157
rect 3513 1152 3582 1157
rect 3665 1152 3694 1157
rect 3833 1152 3942 1157
rect 4001 1152 4094 1157
rect 1945 1147 1950 1152
rect 2113 1147 2254 1152
rect 3489 1147 3494 1152
rect 1033 1142 1062 1147
rect 1081 1142 1190 1147
rect 1201 1142 1318 1147
rect 1537 1142 1798 1147
rect 1825 1142 1950 1147
rect 2273 1142 2670 1147
rect 809 1137 814 1142
rect 1313 1137 1542 1142
rect 2817 1137 2822 1147
rect 2849 1142 2942 1147
rect 3001 1142 3030 1147
rect 3185 1142 3246 1147
rect 3297 1142 3334 1147
rect 3433 1142 3478 1147
rect 3489 1142 3622 1147
rect 2937 1137 3006 1142
rect 3617 1137 3622 1142
rect 3745 1142 3774 1147
rect 3793 1142 3854 1147
rect 3865 1142 3918 1147
rect 4017 1142 4078 1147
rect 3745 1137 3750 1142
rect 385 1132 406 1137
rect 385 1122 390 1132
rect 641 1127 646 1137
rect 697 1132 814 1137
rect 833 1132 902 1137
rect 1009 1132 1030 1137
rect 641 1122 670 1127
rect 833 1122 838 1132
rect 1009 1127 1014 1132
rect 857 1122 1014 1127
rect 1025 1127 1030 1132
rect 1153 1132 1294 1137
rect 1561 1132 1606 1137
rect 1713 1132 1766 1137
rect 1969 1132 1998 1137
rect 2025 1132 2142 1137
rect 2161 1132 2238 1137
rect 2817 1132 2862 1137
rect 3193 1132 3262 1137
rect 3313 1132 3486 1137
rect 3497 1132 3526 1137
rect 3617 1132 3750 1137
rect 3857 1132 3886 1137
rect 3969 1132 4014 1137
rect 1153 1127 1158 1132
rect 2025 1127 2030 1132
rect 1025 1122 1158 1127
rect 1193 1122 1550 1127
rect 1545 1117 1550 1122
rect 1617 1122 1702 1127
rect 1617 1117 1622 1122
rect 321 1112 366 1117
rect 433 1112 478 1117
rect 497 1112 622 1117
rect 1177 1112 1214 1117
rect 1257 1112 1310 1117
rect 1545 1112 1622 1117
rect 1697 1117 1702 1122
rect 1777 1122 1806 1127
rect 2001 1122 2030 1127
rect 2137 1127 2142 1132
rect 2257 1127 2382 1132
rect 2417 1127 2606 1132
rect 2137 1122 2262 1127
rect 2377 1122 2422 1127
rect 2601 1122 2630 1127
rect 2657 1122 2710 1127
rect 2945 1122 3494 1127
rect 1777 1117 1782 1122
rect 2809 1117 2894 1122
rect 3521 1117 3526 1132
rect 3537 1122 3598 1127
rect 3993 1122 4126 1127
rect 1697 1112 1782 1117
rect 1841 1112 1862 1117
rect 1985 1112 2166 1117
rect 2193 1112 2310 1117
rect 2321 1112 2366 1117
rect 2433 1112 2518 1117
rect 2537 1112 2582 1117
rect 2785 1112 2814 1117
rect 2889 1112 2974 1117
rect 3201 1112 3254 1117
rect 3337 1112 3414 1117
rect 3521 1112 3558 1117
rect 3833 1112 3878 1117
rect 3985 1112 4030 1117
rect 2305 1107 2310 1112
rect 465 1102 574 1107
rect 689 1102 814 1107
rect 849 1102 894 1107
rect 913 1102 1158 1107
rect 1905 1102 2118 1107
rect 2153 1102 2190 1107
rect 2305 1102 2334 1107
rect 2369 1102 2638 1107
rect 2665 1102 2726 1107
rect 2809 1102 2838 1107
rect 2849 1102 2878 1107
rect 2993 1102 3182 1107
rect 3209 1102 3350 1107
rect 3361 1102 3518 1107
rect 3873 1102 3910 1107
rect 3945 1102 4030 1107
rect 689 1097 694 1102
rect 465 1092 494 1097
rect 585 1092 694 1097
rect 809 1097 814 1102
rect 913 1097 918 1102
rect 809 1092 918 1097
rect 1153 1097 1158 1102
rect 1769 1097 1886 1102
rect 2369 1097 2374 1102
rect 2993 1097 2998 1102
rect 1153 1092 1502 1097
rect 1561 1092 1686 1097
rect 1745 1092 1774 1097
rect 1881 1092 2054 1097
rect 2169 1092 2270 1097
rect 2313 1092 2374 1097
rect 2409 1092 2582 1097
rect 2697 1092 2726 1097
rect 2777 1092 2814 1097
rect 2833 1092 2862 1097
rect 2913 1092 2998 1097
rect 3177 1097 3182 1102
rect 3177 1092 3278 1097
rect 3457 1092 3638 1097
rect 2577 1087 2702 1092
rect 473 1082 542 1087
rect 577 1082 686 1087
rect 705 1082 1078 1087
rect 1113 1082 1134 1087
rect 1801 1082 2182 1087
rect 2433 1082 2470 1087
rect 2505 1082 2558 1087
rect 2937 1082 3246 1087
rect 1153 1077 1222 1082
rect 1297 1077 1518 1082
rect 1577 1077 1686 1082
rect 345 1072 446 1077
rect 601 1072 1158 1077
rect 1217 1072 1302 1077
rect 1513 1072 1542 1077
rect 1553 1072 1582 1077
rect 1681 1072 1758 1077
rect 2129 1072 2390 1077
rect 2401 1072 2734 1077
rect 2809 1072 2998 1077
rect 3665 1072 3694 1077
rect 3953 1072 3998 1077
rect 345 1067 350 1072
rect 321 1062 350 1067
rect 441 1067 446 1072
rect 1777 1067 2134 1072
rect 441 1062 1206 1067
rect 1313 1062 1782 1067
rect 2145 1062 2182 1067
rect 2241 1062 2526 1067
rect 2521 1057 2526 1062
rect 2649 1062 3062 1067
rect 2649 1057 2654 1062
rect 3057 1057 3062 1062
rect 3169 1062 3198 1067
rect 3401 1062 3550 1067
rect 3169 1057 3174 1062
rect 3401 1057 3406 1062
rect 649 1052 1270 1057
rect 1313 1052 2486 1057
rect 2521 1052 2654 1057
rect 2673 1052 2694 1057
rect 2761 1052 2902 1057
rect 3009 1052 3038 1057
rect 3057 1052 3174 1057
rect 3377 1052 3406 1057
rect 3545 1057 3550 1062
rect 3545 1052 3574 1057
rect 3625 1052 3678 1057
rect 3785 1052 3862 1057
rect 1313 1047 1318 1052
rect 2897 1047 3014 1052
rect 3425 1047 3526 1052
rect 329 1042 454 1047
rect 633 1042 1318 1047
rect 1625 1042 1694 1047
rect 1761 1042 2502 1047
rect 2721 1042 2878 1047
rect 3353 1042 3430 1047
rect 3521 1042 3614 1047
rect 3633 1042 3790 1047
rect 1465 1037 1534 1042
rect 209 1032 302 1037
rect 545 1032 710 1037
rect 785 1032 1038 1037
rect 1073 1032 1470 1037
rect 1529 1032 1582 1037
rect 1673 1032 1718 1037
rect 1777 1032 1830 1037
rect 2049 1032 2094 1037
rect 2137 1032 2198 1037
rect 2385 1032 2542 1037
rect 2617 1032 2646 1037
rect 2657 1032 2974 1037
rect 3329 1032 3766 1037
rect 209 1027 214 1032
rect 121 1022 174 1027
rect 185 1022 214 1027
rect 297 1027 302 1032
rect 1849 1027 2030 1032
rect 2193 1027 2390 1032
rect 297 1022 326 1027
rect 481 1022 526 1027
rect 729 1022 774 1027
rect 873 1022 910 1027
rect 961 1022 982 1027
rect 1057 1022 1110 1027
rect 1201 1022 1230 1027
rect 1481 1022 1854 1027
rect 2025 1022 2174 1027
rect 2409 1022 2462 1027
rect 2481 1022 2782 1027
rect 2817 1022 2910 1027
rect 3017 1022 3078 1027
rect 3393 1022 3526 1027
rect 3593 1022 3734 1027
rect 4025 1022 4150 1027
rect 1225 1017 1230 1022
rect 1297 1017 1486 1022
rect 233 1012 406 1017
rect 545 1012 606 1017
rect 689 1012 982 1017
rect 1225 1012 1302 1017
rect 1505 1012 1534 1017
rect 1665 1012 1726 1017
rect 1737 1012 1766 1017
rect 1777 1012 2326 1017
rect 2345 1012 2622 1017
rect 2729 1012 2774 1017
rect 2841 1012 2862 1017
rect 2873 1012 3014 1017
rect 3089 1012 3150 1017
rect 3321 1012 3366 1017
rect 3385 1012 3470 1017
rect 425 1007 526 1012
rect 169 1002 206 1007
rect 385 1002 430 1007
rect 521 1002 654 1007
rect 721 1002 806 1007
rect 897 1002 958 1007
rect 1057 1002 1174 1007
rect 1321 1002 1478 1007
rect 1505 1002 1566 1007
rect 1657 1002 1694 1007
rect 1745 1002 2046 1007
rect 2145 1002 2286 1007
rect 1321 997 1326 1002
rect 161 992 398 997
rect 449 992 478 997
rect 513 992 566 997
rect 609 992 646 997
rect 753 992 774 997
rect 873 992 934 997
rect 1233 992 1326 997
rect 1473 997 1478 1002
rect 2321 997 2326 1012
rect 3009 1007 3094 1012
rect 3609 1007 3614 1017
rect 3721 1012 3742 1017
rect 3961 1012 4006 1017
rect 2401 1002 2430 1007
rect 2505 1002 2542 1007
rect 2625 1002 2654 1007
rect 2833 1002 2902 1007
rect 2921 1002 2990 1007
rect 3193 1002 3238 1007
rect 3257 1002 3334 1007
rect 3345 1002 3462 1007
rect 3529 1002 3598 1007
rect 3609 1002 3734 1007
rect 2537 997 2630 1002
rect 1473 992 1822 997
rect 1945 992 2230 997
rect 2321 992 2446 997
rect 2497 992 2518 997
rect 2665 992 2782 997
rect 2817 992 2894 997
rect 3009 992 3086 997
rect 3313 992 3430 997
rect 3505 992 3550 997
rect 3585 992 3662 997
rect 3753 992 3814 997
rect 4017 992 4078 997
rect 1817 987 1950 992
rect 745 982 822 987
rect 905 982 942 987
rect 1337 982 1462 987
rect 1697 982 1742 987
rect 1761 982 1798 987
rect 1969 982 2006 987
rect 2081 982 2134 987
rect 2161 982 2190 987
rect 2201 982 2294 987
rect 2377 982 2422 987
rect 2433 982 2462 987
rect 2577 982 2702 987
rect 2793 982 2846 987
rect 2873 982 2918 987
rect 2961 982 3022 987
rect 3105 982 3286 987
rect 3305 982 3398 987
rect 3409 982 3438 987
rect 3561 982 3590 987
rect 3625 982 3670 987
rect 3681 982 3758 987
rect 337 977 414 982
rect 553 977 726 982
rect 1569 977 1678 982
rect 1969 977 1974 982
rect 2417 977 2422 982
rect 3105 977 3110 982
rect 105 972 342 977
rect 409 972 438 977
rect 529 972 558 977
rect 721 972 846 977
rect 865 972 894 977
rect 889 967 894 972
rect 953 972 1070 977
rect 1273 972 1574 977
rect 1673 972 1774 977
rect 1785 972 1814 977
rect 1833 972 1974 977
rect 1985 972 2078 977
rect 2097 972 2270 977
rect 2305 972 2406 977
rect 2417 972 2630 977
rect 2705 972 2742 977
rect 2761 972 2822 977
rect 2833 972 2862 977
rect 3081 972 3110 977
rect 3281 977 3286 982
rect 3393 977 3398 982
rect 3281 972 3382 977
rect 3393 972 3438 977
rect 3537 972 3582 977
rect 3793 972 3822 977
rect 953 967 958 972
rect 1833 967 1838 972
rect 2817 967 2822 972
rect 2881 967 3006 972
rect 3129 967 3262 972
rect 3601 967 3774 972
rect 353 962 726 967
rect 889 962 958 967
rect 1073 962 1198 967
rect 1217 962 1246 967
rect 1353 962 1414 967
rect 1465 962 1494 967
rect 1585 962 1838 967
rect 2001 962 2414 967
rect 2497 962 2590 967
rect 2601 962 2622 967
rect 2697 962 2790 967
rect 2817 962 2886 967
rect 3001 962 3030 967
rect 3041 962 3134 967
rect 3257 962 3326 967
rect 3369 962 3406 967
rect 3433 962 3606 967
rect 3769 962 3822 967
rect 233 957 334 962
rect 1241 957 1358 962
rect 209 952 238 957
rect 329 952 374 957
rect 505 952 542 957
rect 553 952 638 957
rect 737 952 766 957
rect 1433 952 1462 957
rect 1601 952 1654 957
rect 1705 952 1758 957
rect 1769 952 2046 957
rect 2065 952 2670 957
rect 2713 952 3446 957
rect 3585 952 3614 957
rect 3665 952 3886 957
rect 633 947 742 952
rect 3441 947 3590 952
rect 81 942 110 947
rect 185 942 230 947
rect 289 942 502 947
rect 569 942 614 947
rect 849 942 958 947
rect 1017 942 1126 947
rect 1289 942 1318 947
rect 1473 942 1590 947
rect 225 937 230 942
rect 1313 937 1318 942
rect 1401 937 1478 942
rect 1585 937 1590 942
rect 1705 942 1830 947
rect 1921 942 2334 947
rect 2401 942 2430 947
rect 1705 937 1710 942
rect 1825 937 1926 942
rect 2425 937 2430 942
rect 2521 942 2710 947
rect 2729 942 2774 947
rect 2801 942 3078 947
rect 3177 942 3310 947
rect 3321 942 3422 947
rect 3657 942 3686 947
rect 3817 942 3934 947
rect 2521 937 2526 942
rect 161 932 206 937
rect 225 932 310 937
rect 345 932 366 937
rect 585 932 726 937
rect 1033 932 1214 937
rect 1225 932 1294 937
rect 1313 932 1406 937
rect 1585 932 1710 937
rect 1729 932 1806 937
rect 1945 932 1982 937
rect 2041 932 2406 937
rect 2425 932 2526 937
rect 2545 932 2574 937
rect 2681 932 2710 937
rect 209 922 238 927
rect 249 922 294 927
rect 129 912 230 917
rect 305 877 310 932
rect 329 922 358 927
rect 369 922 414 927
rect 481 922 534 927
rect 553 922 582 927
rect 1065 922 1254 927
rect 1817 922 1910 927
rect 1937 922 2030 927
rect 2065 922 2150 927
rect 2161 922 2390 927
rect 2401 917 2406 932
rect 2745 927 2750 937
rect 2761 932 2870 937
rect 2865 927 2870 932
rect 3025 932 3054 937
rect 3065 932 3134 937
rect 3225 932 3254 937
rect 3025 927 3030 932
rect 3249 927 3254 932
rect 3345 932 3374 937
rect 3385 932 3534 937
rect 3345 927 3350 932
rect 3809 927 3958 932
rect 2593 922 2662 927
rect 2729 922 2750 927
rect 2785 922 2846 927
rect 2865 922 3030 927
rect 3105 922 3198 927
rect 3249 922 3350 927
rect 3393 922 3414 927
rect 3785 922 3814 927
rect 3953 922 3982 927
rect 3105 917 3110 922
rect 337 912 430 917
rect 449 912 566 917
rect 617 912 662 917
rect 777 912 902 917
rect 921 912 942 917
rect 1193 912 1238 917
rect 1273 912 1358 917
rect 777 907 782 912
rect 409 902 782 907
rect 897 907 902 912
rect 1273 907 1278 912
rect 897 902 1278 907
rect 1353 907 1358 912
rect 1425 912 1710 917
rect 1777 912 1830 917
rect 1921 912 1950 917
rect 1985 912 2006 917
rect 2041 912 2102 917
rect 2137 912 2254 917
rect 2401 912 2526 917
rect 2561 912 2590 917
rect 2641 912 2686 917
rect 2793 912 2822 917
rect 3049 912 3110 917
rect 3489 912 3534 917
rect 3633 912 3678 917
rect 3825 912 3894 917
rect 3913 912 4046 917
rect 1425 907 1430 912
rect 1353 902 1430 907
rect 1705 907 1710 912
rect 2521 907 2526 912
rect 1705 902 1766 907
rect 1801 902 1822 907
rect 1841 902 1966 907
rect 2105 902 2358 907
rect 2521 902 3038 907
rect 3121 902 3702 907
rect 3809 902 3838 907
rect 1993 897 2086 902
rect 3033 897 3126 902
rect 353 892 406 897
rect 449 892 478 897
rect 609 892 638 897
rect 857 892 974 897
rect 1177 892 1206 897
rect 1313 892 1342 897
rect 1441 892 1998 897
rect 2081 892 2326 897
rect 2417 892 2670 897
rect 2681 892 2710 897
rect 2809 892 2870 897
rect 3281 892 3310 897
rect 3465 892 3494 897
rect 3625 892 3870 897
rect 473 887 614 892
rect 1201 887 1318 892
rect 2321 887 2422 892
rect 793 882 878 887
rect 921 882 1166 887
rect 1833 882 1934 887
rect 2009 882 2214 887
rect 2249 882 2302 887
rect 2537 882 2574 887
rect 2633 882 2662 887
rect 2745 882 2838 887
rect 3113 882 3190 887
rect 3417 882 3478 887
rect 3601 882 3638 887
rect 3657 882 3774 887
rect 1433 877 1814 882
rect 305 872 822 877
rect 945 872 974 877
rect 1257 872 1438 877
rect 1809 872 2566 877
rect 2577 872 2622 877
rect 2649 872 2670 877
rect 2777 872 2910 877
rect 3273 872 3406 877
rect 3513 872 3558 877
rect 3697 872 3790 877
rect 1449 862 1782 867
rect 1793 862 2102 867
rect 2113 862 2142 867
rect 2169 862 2230 867
rect 2281 862 2318 867
rect 2921 862 2990 867
rect 3217 862 3334 867
rect 3401 862 3502 867
rect 3569 862 3838 867
rect 3857 862 3934 867
rect 1777 857 1782 862
rect 3497 857 3574 862
rect 3857 857 3862 862
rect 329 852 366 857
rect 593 852 854 857
rect 873 852 1206 857
rect 1225 852 1270 857
rect 1385 852 1438 857
rect 1609 852 1670 857
rect 1777 852 1814 857
rect 1841 852 1862 857
rect 1945 852 2366 857
rect 2449 852 2502 857
rect 2521 852 2622 857
rect 2721 852 2766 857
rect 3009 852 3046 857
rect 3153 852 3278 857
rect 3377 852 3406 857
rect 3817 852 3862 857
rect 3929 857 3934 862
rect 3929 852 4046 857
rect 873 847 878 852
rect 385 842 574 847
rect 817 842 878 847
rect 1201 847 1206 852
rect 1457 847 1590 852
rect 2521 847 2526 852
rect 1201 842 1350 847
rect 1417 842 1462 847
rect 1585 842 1886 847
rect 1921 842 2526 847
rect 2617 847 2622 852
rect 3377 847 3382 852
rect 2617 842 2710 847
rect 2825 842 2886 847
rect 2985 842 3166 847
rect 3329 842 3382 847
rect 3401 847 3406 852
rect 3705 847 3822 852
rect 3401 842 3710 847
rect 3841 842 3886 847
rect 385 837 390 842
rect 177 832 390 837
rect 569 837 574 842
rect 569 832 1302 837
rect 1297 827 1302 832
rect 1361 832 1982 837
rect 2073 832 2318 837
rect 2329 832 2606 837
rect 2993 832 3206 837
rect 3233 832 3270 837
rect 3289 832 3382 837
rect 3729 832 3782 837
rect 3801 832 3918 837
rect 1361 827 1366 832
rect 129 822 174 827
rect 433 822 486 827
rect 497 822 542 827
rect 673 822 718 827
rect 865 822 894 827
rect 1057 822 1102 827
rect 1153 822 1214 827
rect 1249 822 1278 827
rect 1297 822 1366 827
rect 1465 822 1510 827
rect 1681 822 1774 827
rect 1785 822 1814 827
rect 1897 822 1958 827
rect 1969 822 2086 827
rect 2129 822 2230 827
rect 2305 822 2342 827
rect 2393 822 2430 827
rect 2713 822 2894 827
rect 3001 822 3158 827
rect 3177 822 3198 827
rect 3225 822 3286 827
rect 3473 822 3542 827
rect 193 817 358 822
rect 2449 817 2526 822
rect 3473 817 3478 822
rect 81 812 198 817
rect 353 812 454 817
rect 545 812 574 817
rect 761 812 814 817
rect 849 812 1014 817
rect 1113 812 1262 817
rect 1489 812 1678 817
rect 1785 812 1878 817
rect 1913 812 2454 817
rect 2521 812 2742 817
rect 2977 812 3246 817
rect 3449 812 3478 817
rect 3537 817 3542 822
rect 3577 822 3710 827
rect 3769 822 3830 827
rect 4017 822 4070 827
rect 3577 817 3582 822
rect 3537 812 3582 817
rect 3705 817 3710 822
rect 3705 812 3894 817
rect 161 802 334 807
rect 1081 802 1110 807
rect 1105 797 1110 802
rect 1169 802 1366 807
rect 1641 802 1710 807
rect 1737 802 1766 807
rect 1865 802 1894 807
rect 2025 802 2086 807
rect 2097 802 2174 807
rect 2377 802 2510 807
rect 2665 802 2734 807
rect 2761 802 2806 807
rect 2913 802 2974 807
rect 3017 802 3094 807
rect 3105 802 3414 807
rect 3737 802 3854 807
rect 3913 802 3966 807
rect 1169 797 1174 802
rect 1761 797 1870 802
rect 2169 797 2262 802
rect 2529 797 2622 802
rect 3409 797 3414 802
rect 201 792 230 797
rect 345 792 590 797
rect 625 792 662 797
rect 705 792 782 797
rect 849 792 966 797
rect 1105 792 1174 797
rect 1217 792 1382 797
rect 1433 792 1486 797
rect 1897 792 2014 797
rect 2113 792 2150 797
rect 225 787 350 792
rect 2257 787 2262 797
rect 2281 792 2534 797
rect 2617 792 2734 797
rect 2817 792 3238 797
rect 3409 792 3526 797
rect 3593 792 3686 797
rect 3857 792 4134 797
rect 2729 787 2822 792
rect 521 782 894 787
rect 961 782 1006 787
rect 1193 782 1342 787
rect 1753 782 1878 787
rect 1985 782 2118 787
rect 2145 782 2174 787
rect 2257 782 2414 787
rect 2521 782 2606 787
rect 2681 782 2710 787
rect 2881 782 3198 787
rect 3209 782 3334 787
rect 3345 782 3486 787
rect 3681 782 3710 787
rect 3881 782 3998 787
rect 4041 782 4070 787
rect 257 772 278 777
rect 321 772 382 777
rect 553 772 870 777
rect 1097 772 1126 777
rect 1137 772 1190 777
rect 1345 772 1550 777
rect 1649 772 1702 777
rect 1825 772 1878 777
rect 1961 772 2110 777
rect 2545 772 2566 777
rect 2577 772 2614 777
rect 2785 772 2814 777
rect 2889 772 2958 777
rect 2993 772 3046 777
rect 3137 772 3454 777
rect 3665 772 3702 777
rect 3817 772 3982 777
rect 377 767 382 772
rect 473 767 558 772
rect 889 767 1078 772
rect 1209 767 1326 772
rect 2273 767 2398 772
rect 2577 767 2582 772
rect 297 762 358 767
rect 377 762 478 767
rect 577 762 894 767
rect 1073 762 1214 767
rect 1321 762 1374 767
rect 1561 762 1814 767
rect 1889 762 1950 767
rect 2017 762 2278 767
rect 2393 762 2582 767
rect 2841 762 2886 767
rect 2937 762 2982 767
rect 3169 762 3198 767
rect 3217 762 3278 767
rect 3393 762 3438 767
rect 3449 762 3518 767
rect 3625 762 3886 767
rect 3937 762 3982 767
rect 1369 757 1566 762
rect 1809 757 1894 762
rect 1945 757 2022 762
rect 569 752 646 757
rect 825 752 854 757
rect 865 752 1014 757
rect 1033 752 1350 757
rect 1649 752 1694 757
rect 2041 752 2158 757
rect 2289 752 2382 757
rect 2513 752 2574 757
rect 2625 752 2662 757
rect 2673 752 2782 757
rect 2945 752 2966 757
rect 3017 752 3046 757
rect 3241 752 3318 757
rect 3385 752 3694 757
rect 3713 752 3790 757
rect 3889 752 3950 757
rect 641 747 830 752
rect 3041 747 3046 752
rect 177 742 302 747
rect 497 742 558 747
rect 593 742 622 747
rect 849 742 886 747
rect 993 742 1030 747
rect 1073 742 1206 747
rect 1241 742 1270 747
rect 1265 737 1270 742
rect 1361 742 1462 747
rect 1513 742 1726 747
rect 1865 742 1894 747
rect 1961 742 2702 747
rect 2753 742 2846 747
rect 2969 742 3030 747
rect 3041 742 3094 747
rect 3137 742 3166 747
rect 3185 742 3382 747
rect 3409 742 3478 747
rect 3593 742 3678 747
rect 1361 737 1366 742
rect 145 732 278 737
rect 457 732 486 737
rect 609 727 614 737
rect 705 732 750 737
rect 769 732 910 737
rect 929 732 974 737
rect 1017 732 1150 737
rect 1177 732 1214 737
rect 1265 732 1366 737
rect 1481 732 2054 737
rect 2265 732 2326 737
rect 2545 732 2582 737
rect 2689 732 2726 737
rect 2745 732 2982 737
rect 2993 732 3190 737
rect 3201 732 3246 737
rect 3305 732 3366 737
rect 2049 727 2166 732
rect 2993 727 2998 732
rect 177 722 206 727
rect 473 722 542 727
rect 569 722 614 727
rect 729 722 830 727
rect 977 722 1046 727
rect 1137 722 1190 727
rect 1537 722 1582 727
rect 1593 722 1726 727
rect 1833 722 1878 727
rect 1985 722 2030 727
rect 2161 722 2646 727
rect 2705 722 2790 727
rect 2817 722 2910 727
rect 2969 722 2998 727
rect 3017 722 3070 727
rect 3329 722 3398 727
rect 3713 722 3718 752
rect 3729 742 3798 747
rect 3889 742 3974 747
rect 4009 742 4094 747
rect 3833 732 3878 737
rect 3985 732 4030 737
rect 3769 722 3806 727
rect 849 717 918 722
rect 225 712 270 717
rect 345 712 390 717
rect 513 712 582 717
rect 801 712 854 717
rect 913 712 1126 717
rect 801 707 806 712
rect 1121 707 1126 712
rect 1201 712 1822 717
rect 1889 712 2326 717
rect 2521 712 3630 717
rect 3657 712 3686 717
rect 3801 712 3862 717
rect 1201 707 1206 712
rect 1817 707 1894 712
rect 2321 707 2414 712
rect 377 702 510 707
rect 561 702 806 707
rect 817 702 902 707
rect 969 702 1038 707
rect 1121 702 1206 707
rect 1481 702 1526 707
rect 1561 702 1614 707
rect 1625 702 1670 707
rect 1705 702 1750 707
rect 2001 702 2078 707
rect 2209 702 2254 707
rect 2409 702 2566 707
rect 2593 702 2694 707
rect 2801 702 2830 707
rect 2873 702 2966 707
rect 3025 702 3078 707
rect 3385 702 3454 707
rect 433 692 606 697
rect 673 692 702 697
rect 809 692 886 697
rect 937 692 974 697
rect 993 692 1062 697
rect 1673 692 1734 697
rect 1881 692 2198 697
rect 2257 692 2398 697
rect 2513 692 3358 697
rect 393 682 638 687
rect 729 682 1670 687
rect 1665 677 1670 682
rect 1761 682 1830 687
rect 1945 682 2030 687
rect 2377 682 2438 687
rect 2721 682 2926 687
rect 3001 682 3038 687
rect 3473 682 3734 687
rect 1761 677 1766 682
rect 2473 677 2598 682
rect 3473 677 3478 682
rect 465 672 1118 677
rect 1665 672 1766 677
rect 1793 672 1846 677
rect 1441 667 1566 672
rect 569 662 1446 667
rect 1561 662 1590 667
rect 1841 657 1846 672
rect 2305 672 2366 677
rect 2305 667 2310 672
rect 2041 662 2310 667
rect 2361 667 2366 672
rect 2449 672 2478 677
rect 2593 672 2686 677
rect 2697 672 3086 677
rect 2449 667 2454 672
rect 3081 667 3086 672
rect 3225 672 3478 677
rect 3729 677 3734 682
rect 3729 672 3758 677
rect 3225 667 3230 672
rect 2361 662 2454 667
rect 2513 662 2582 667
rect 2729 662 2766 667
rect 2793 662 2998 667
rect 3081 662 3230 667
rect 2041 657 2046 662
rect 3281 657 3446 662
rect 321 652 446 657
rect 585 652 758 657
rect 857 652 958 657
rect 321 647 326 652
rect 185 642 326 647
rect 441 647 446 652
rect 753 647 862 652
rect 953 647 958 652
rect 1041 652 1150 657
rect 1041 647 1046 652
rect 441 642 574 647
rect 705 642 734 647
rect 881 642 910 647
rect 953 642 1046 647
rect 569 637 710 642
rect 1145 637 1150 652
rect 1457 652 1614 657
rect 1801 652 1822 657
rect 1841 652 2046 657
rect 2737 652 2798 657
rect 2825 652 2886 657
rect 3001 652 3062 657
rect 3257 652 3286 657
rect 3441 652 3758 657
rect 1457 647 1462 652
rect 1353 642 1462 647
rect 2329 642 2526 647
rect 2569 642 2606 647
rect 2705 642 2774 647
rect 2817 642 2838 647
rect 2993 642 3046 647
rect 3249 642 3542 647
rect 3737 642 3846 647
rect 1353 637 1358 642
rect 3537 637 3542 642
rect 3633 637 3742 642
rect 249 632 438 637
rect 761 632 830 637
rect 841 632 934 637
rect 1065 632 1126 637
rect 1145 632 1358 637
rect 1481 632 1534 637
rect 2241 632 2358 637
rect 2529 632 2566 637
rect 2681 632 3214 637
rect 3241 632 3326 637
rect 3385 632 3478 637
rect 3537 632 3638 637
rect 3761 632 3902 637
rect 3945 632 3990 637
rect 145 622 174 627
rect 249 622 294 627
rect 345 622 398 627
rect 441 622 486 627
rect 529 622 574 627
rect 617 622 662 627
rect 833 622 870 627
rect 905 622 950 627
rect 1025 622 1070 627
rect 1393 617 1398 627
rect 1465 622 1510 627
rect 1529 622 1566 627
rect 1585 622 1630 627
rect 1649 622 1678 627
rect 2073 622 2190 627
rect 2289 622 2342 627
rect 2393 622 2470 627
rect 2553 622 2590 627
rect 2657 622 2694 627
rect 2769 622 2846 627
rect 2929 622 2990 627
rect 3001 622 3102 627
rect 3209 622 3294 627
rect 3361 622 3422 627
rect 3457 622 3518 627
rect 3657 622 3718 627
rect 3785 622 3830 627
rect 3881 622 3942 627
rect 2393 617 2398 622
rect 161 612 238 617
rect 489 612 542 617
rect 745 612 814 617
rect 873 612 902 617
rect 985 612 1014 617
rect 1121 612 1190 617
rect 233 607 494 612
rect 897 607 990 612
rect 1121 607 1126 612
rect 137 602 174 607
rect 513 602 590 607
rect 649 602 726 607
rect 849 602 878 607
rect 1089 602 1126 607
rect 1185 607 1190 612
rect 1377 612 1398 617
rect 1513 612 1534 617
rect 1601 612 1718 617
rect 1737 612 1886 617
rect 1905 612 1942 617
rect 1961 612 2054 617
rect 2369 612 2398 617
rect 2465 617 2470 622
rect 4145 617 4150 627
rect 2465 612 2494 617
rect 2505 612 2614 617
rect 2905 612 2942 617
rect 2961 612 3038 617
rect 3281 612 3326 617
rect 3369 612 3430 617
rect 3441 612 3494 617
rect 3537 612 3638 617
rect 3745 612 3798 617
rect 3833 612 3862 617
rect 3953 612 4150 617
rect 1185 602 1214 607
rect 1297 602 1366 607
rect 649 597 654 602
rect 113 592 254 597
rect 281 592 502 597
rect 577 592 654 597
rect 721 597 726 602
rect 753 597 854 602
rect 721 592 758 597
rect 977 592 1054 597
rect 1137 592 1190 597
rect 665 582 766 587
rect 881 582 958 587
rect 129 577 374 582
rect 881 577 886 582
rect 81 572 134 577
rect 369 572 398 577
rect 521 572 798 577
rect 857 572 886 577
rect 953 577 958 582
rect 953 572 1062 577
rect 1377 572 1382 612
rect 1737 607 1742 612
rect 1393 602 1742 607
rect 1881 607 1886 612
rect 1961 607 1966 612
rect 1881 602 1966 607
rect 2049 607 2054 612
rect 2225 607 2326 612
rect 2689 607 2830 612
rect 2961 607 2966 612
rect 3441 607 3446 612
rect 3537 607 3542 612
rect 2049 602 2230 607
rect 2321 602 2694 607
rect 2825 602 2966 607
rect 3057 602 3198 607
rect 3265 602 3302 607
rect 3441 602 3470 607
rect 3481 602 3542 607
rect 3633 607 3638 612
rect 3857 607 3958 612
rect 3633 602 3702 607
rect 3057 597 3062 602
rect 1497 592 1550 597
rect 1633 592 1662 597
rect 1969 592 2006 597
rect 2065 592 2126 597
rect 2233 592 2310 597
rect 2377 592 2414 597
rect 2497 592 2542 597
rect 2561 592 2622 597
rect 2705 592 3062 597
rect 3193 597 3198 602
rect 3193 592 3222 597
rect 3233 592 3382 597
rect 3393 592 3494 597
rect 3585 592 3678 597
rect 3705 592 3734 597
rect 3857 592 3910 597
rect 4017 592 4078 597
rect 1721 587 1814 592
rect 3081 587 3174 592
rect 3393 587 3398 592
rect 3489 587 3494 592
rect 1577 582 1726 587
rect 1809 582 1902 587
rect 1953 582 1990 587
rect 2041 582 2350 587
rect 2393 582 2582 587
rect 2625 582 2758 587
rect 2985 582 3086 587
rect 3169 582 3398 587
rect 3441 582 3478 587
rect 3489 582 3694 587
rect 3817 582 3878 587
rect 3897 582 4006 587
rect 2777 577 2966 582
rect 1625 572 1670 577
rect 1737 572 1798 577
rect 2313 572 2478 577
rect 2497 572 2646 577
rect 2745 572 2782 577
rect 2961 572 3782 577
rect 3881 572 3926 577
rect 1057 567 1062 572
rect 2497 567 2502 572
rect 2641 567 2726 572
rect 169 562 222 567
rect 265 562 574 567
rect 681 562 958 567
rect 985 562 1046 567
rect 1057 562 1510 567
rect 1617 562 1910 567
rect 2361 562 2502 567
rect 2593 562 2622 567
rect 2721 562 3406 567
rect 569 557 686 562
rect 3401 557 3406 562
rect 3465 562 3542 567
rect 3593 562 3646 567
rect 3673 562 3766 567
rect 3865 562 3918 567
rect 3465 557 3470 562
rect 337 552 358 557
rect 441 552 550 557
rect 705 552 742 557
rect 753 552 862 557
rect 889 552 950 557
rect 1721 552 1846 557
rect 2209 552 2302 557
rect 2353 552 2398 557
rect 2489 552 2734 557
rect 753 547 758 552
rect 2729 547 2734 552
rect 2833 552 2862 557
rect 3097 552 3150 557
rect 3401 552 3470 557
rect 3505 552 3542 557
rect 3697 552 3822 557
rect 3889 552 3918 557
rect 3929 552 4102 557
rect 2833 547 2838 552
rect 161 542 230 547
rect 601 542 758 547
rect 809 542 870 547
rect 1217 542 1246 547
rect 1505 542 1606 547
rect 1737 542 1766 547
rect 1817 542 1862 547
rect 1929 542 2030 547
rect 2049 542 2214 547
rect 2313 542 2366 547
rect 2481 542 2710 547
rect 2729 542 2838 547
rect 2985 542 3134 547
rect 3193 542 3342 547
rect 3489 542 3518 547
rect 3689 542 3742 547
rect 3913 542 3990 547
rect 1505 537 1510 542
rect 1929 537 1934 542
rect 201 532 238 537
rect 305 532 350 537
rect 593 527 598 537
rect 1001 532 1030 537
rect 1057 532 1094 537
rect 1289 532 1358 537
rect 1489 532 1510 537
rect 1769 532 1934 537
rect 2025 537 2030 542
rect 2313 537 2318 542
rect 2025 532 2318 537
rect 2337 527 2342 537
rect 2433 532 2518 537
rect 2617 532 2686 537
rect 2913 532 2974 537
rect 3113 532 3190 537
rect 3201 532 3254 537
rect 3521 532 3574 537
rect 3625 532 3654 537
rect 3865 532 4070 537
rect 497 522 574 527
rect 593 522 670 527
rect 953 522 998 527
rect 1033 522 1110 527
rect 1129 522 1246 527
rect 1409 522 1454 527
rect 1513 522 1606 527
rect 1737 522 1782 527
rect 1905 522 1942 527
rect 2337 522 2366 527
rect 2521 522 2550 527
rect 2809 522 2830 527
rect 2849 522 3078 527
rect 3121 522 3174 527
rect 3329 522 3358 527
rect 3377 522 3678 527
rect 3713 522 3862 527
rect 3897 522 4054 527
rect 497 517 502 522
rect 129 512 174 517
rect 201 512 390 517
rect 409 512 454 517
rect 473 512 502 517
rect 569 517 574 522
rect 1129 517 1134 522
rect 569 512 598 517
rect 649 512 694 517
rect 713 512 814 517
rect 873 512 902 517
rect 929 512 966 517
rect 1065 512 1134 517
rect 1241 517 1246 522
rect 1985 517 2094 522
rect 2217 517 2318 522
rect 2545 517 2550 522
rect 3713 517 3718 522
rect 1241 512 1342 517
rect 1457 512 1502 517
rect 1593 512 1646 517
rect 1721 512 1766 517
rect 1961 512 1990 517
rect 2089 512 2174 517
rect 2193 512 2222 517
rect 2313 512 2486 517
rect 2545 512 2822 517
rect 3041 512 3166 517
rect 3265 512 3334 517
rect 3513 512 3566 517
rect 3609 512 3718 517
rect 3857 512 3950 517
rect 385 497 390 512
rect 713 507 718 512
rect 689 502 718 507
rect 809 507 814 512
rect 2841 507 3022 512
rect 809 502 838 507
rect 969 502 990 507
rect 1041 502 1110 507
rect 1129 502 1230 507
rect 1633 502 1830 507
rect 1945 502 2846 507
rect 3017 502 3062 507
rect 3169 502 3198 507
rect 3345 502 3406 507
rect 521 497 694 502
rect 1417 497 1614 502
rect 3057 497 3174 502
rect 385 492 526 497
rect 833 492 1422 497
rect 1609 492 1926 497
rect 1937 492 1982 497
rect 2025 492 2070 497
rect 2273 492 2326 497
rect 2577 492 3038 497
rect 2089 487 2278 492
rect 2345 487 2558 492
rect 545 482 710 487
rect 729 482 822 487
rect 993 482 1086 487
rect 1433 482 2094 487
rect 2297 482 2350 487
rect 2553 482 2942 487
rect 3057 482 3326 487
rect 817 477 894 482
rect 993 477 998 482
rect 1121 477 1318 482
rect 2961 477 3062 482
rect 3321 477 3326 482
rect 889 472 998 477
rect 1097 472 1126 477
rect 1313 472 1342 477
rect 1537 472 1582 477
rect 1617 472 1646 477
rect 1993 472 2054 477
rect 2065 472 2710 477
rect 2721 472 2758 477
rect 2769 472 2966 477
rect 3321 472 3382 477
rect 1361 467 1430 472
rect 1665 467 1974 472
rect 2705 467 2710 472
rect 3081 467 3198 472
rect 553 462 782 467
rect 841 462 870 467
rect 1017 462 1366 467
rect 1425 462 1670 467
rect 1969 462 2462 467
rect 2705 462 2766 467
rect 2889 462 3086 467
rect 3193 462 3462 467
rect 3481 462 3798 467
rect 2537 457 2686 462
rect 2761 457 2894 462
rect 753 452 1006 457
rect 1001 447 1006 452
rect 1097 452 1414 457
rect 1585 452 1902 457
rect 1921 452 2398 457
rect 2457 452 2494 457
rect 2513 452 2542 457
rect 2681 452 2742 457
rect 2913 452 2958 457
rect 3025 452 3270 457
rect 3481 452 3486 462
rect 1097 447 1102 452
rect 1409 447 1574 452
rect 3369 447 3486 452
rect 3793 447 3798 462
rect 465 442 558 447
rect 593 442 630 447
rect 817 442 974 447
rect 1001 442 1102 447
rect 1121 442 1174 447
rect 1569 442 1878 447
rect 1953 442 1982 447
rect 2393 442 2838 447
rect 2913 442 2998 447
rect 3009 442 3318 447
rect 3345 442 3374 447
rect 3641 442 3774 447
rect 3793 442 3822 447
rect 1249 437 1390 442
rect 1977 437 2398 442
rect 3641 437 3646 442
rect 441 432 518 437
rect 577 432 614 437
rect 873 432 918 437
rect 1225 432 1254 437
rect 1385 432 1414 437
rect 1529 432 1566 437
rect 1585 432 1798 437
rect 1865 432 1886 437
rect 1905 432 1942 437
rect 2417 432 2438 437
rect 2545 432 2686 437
rect 2945 432 3046 437
rect 3129 432 3238 437
rect 3321 432 3646 437
rect 3769 437 3774 442
rect 3769 432 4014 437
rect 937 427 1030 432
rect 1585 427 1590 432
rect 2545 427 2550 432
rect 2945 427 2950 432
rect 193 422 222 427
rect 281 422 326 427
rect 409 422 454 427
rect 537 422 574 427
rect 601 422 670 427
rect 777 422 942 427
rect 1025 422 1590 427
rect 1601 422 1638 427
rect 1801 422 1862 427
rect 1961 422 2038 427
rect 2153 422 2182 427
rect 2257 422 2334 427
rect 2393 422 2550 427
rect 2569 422 2614 427
rect 2841 422 2950 427
rect 2977 422 3030 427
rect 3057 422 3134 427
rect 3201 422 3254 427
rect 3265 422 3542 427
rect 3657 422 3814 427
rect 1657 417 1734 422
rect 1881 417 1966 422
rect 2033 417 2038 422
rect 3025 417 3030 422
rect 209 412 238 417
rect 337 412 478 417
rect 689 412 742 417
rect 785 412 846 417
rect 913 412 1014 417
rect 1377 412 1662 417
rect 1729 412 1886 417
rect 2033 412 2142 417
rect 2385 412 2478 417
rect 2553 412 2654 417
rect 2705 412 2758 417
rect 2937 412 3014 417
rect 3025 412 3054 417
rect 3241 412 3526 417
rect 233 407 342 412
rect 1273 407 1358 412
rect 3129 407 3222 412
rect 3537 407 3542 422
rect 3553 412 3710 417
rect 129 402 206 407
rect 545 402 646 407
rect 993 402 1038 407
rect 1177 402 1278 407
rect 1353 402 1414 407
rect 1497 402 1542 407
rect 1609 402 1694 407
rect 1817 402 2022 407
rect 2433 402 2470 407
rect 2545 402 2574 407
rect 2681 402 2766 407
rect 2801 402 3134 407
rect 3217 402 3478 407
rect 3537 402 3846 407
rect 1817 397 1822 402
rect 3473 397 3478 402
rect 161 392 302 397
rect 337 392 438 397
rect 529 392 574 397
rect 753 392 806 397
rect 817 392 854 397
rect 865 392 918 397
rect 953 392 1014 397
rect 1289 392 1366 397
rect 1393 392 1430 397
rect 1713 392 1822 397
rect 1841 392 1878 397
rect 1929 392 1958 397
rect 1977 392 2094 397
rect 2161 392 2286 397
rect 2449 392 2494 397
rect 2625 392 2654 397
rect 2905 392 2958 397
rect 2969 392 3014 397
rect 3145 392 3206 397
rect 3265 392 3334 397
rect 3385 392 3454 397
rect 3473 392 3558 397
rect 3625 392 3662 397
rect 3673 392 3734 397
rect 3833 392 3910 397
rect 4009 392 4086 397
rect 1561 387 1718 392
rect 657 382 710 387
rect 737 382 1230 387
rect 1377 382 1566 387
rect 2161 382 2166 392
rect 345 377 638 382
rect 1825 377 1950 382
rect 2001 377 2166 382
rect 2281 377 2286 392
rect 2329 382 2414 387
rect 2441 382 2470 387
rect 2481 382 2774 387
rect 2857 382 2950 387
rect 2985 382 3126 387
rect 3169 382 3430 387
rect 3641 382 3702 387
rect 3889 382 3926 387
rect 3953 382 4062 387
rect 2329 377 2334 382
rect 281 372 350 377
rect 633 372 670 377
rect 665 367 670 372
rect 801 372 1102 377
rect 1385 372 1406 377
rect 1417 372 1446 377
rect 1577 372 1830 377
rect 1945 372 2006 377
rect 2281 372 2334 377
rect 2409 377 2414 382
rect 2481 377 2486 382
rect 3721 377 3870 382
rect 2409 372 2486 377
rect 2577 372 3006 377
rect 3049 372 3262 377
rect 3561 372 3598 377
rect 3609 372 3638 377
rect 3657 372 3726 377
rect 3865 372 3974 377
rect 801 367 806 372
rect 1441 367 1582 372
rect 2577 367 2582 372
rect 3281 367 3366 372
rect 361 362 646 367
rect 665 362 806 367
rect 841 362 974 367
rect 985 362 1022 367
rect 1073 362 1126 367
rect 1145 362 1358 367
rect 1601 362 1662 367
rect 1841 362 1934 367
rect 2017 362 2582 367
rect 2593 362 3286 367
rect 3361 362 3606 367
rect 3657 362 3854 367
rect 1145 357 1150 362
rect 193 352 598 357
rect 825 352 862 357
rect 913 352 958 357
rect 1001 352 1150 357
rect 1353 357 1358 362
rect 1657 357 1846 362
rect 1353 352 1638 357
rect 1865 352 1886 357
rect 1945 352 1998 357
rect 2049 352 2094 357
rect 2137 352 2510 357
rect 2665 352 2750 357
rect 2849 352 2950 357
rect 3017 352 3158 357
rect 3217 352 3262 357
rect 3321 352 3350 357
rect 3585 352 3694 357
rect 3817 352 4030 357
rect 913 347 918 352
rect 329 342 366 347
rect 449 342 622 347
rect 737 342 918 347
rect 937 342 974 347
rect 1033 342 1094 347
rect 1129 342 1254 347
rect 1273 342 1350 347
rect 1361 342 1422 347
rect 1513 342 1582 347
rect 1697 342 1750 347
rect 1833 342 1886 347
rect 1969 342 2006 347
rect 2073 342 2134 347
rect 2177 342 2206 347
rect 2249 342 2326 347
rect 2385 342 2590 347
rect 2689 342 2766 347
rect 2833 342 2862 347
rect 2905 342 2982 347
rect 3025 342 3078 347
rect 3225 342 3254 347
rect 3273 342 3342 347
rect 3457 342 3662 347
rect 3673 342 3734 347
rect 3801 342 3910 347
rect 3921 342 3982 347
rect 201 332 238 337
rect 249 332 294 337
rect 993 332 1062 337
rect 1153 332 1270 337
rect 1289 332 1382 337
rect 585 327 742 332
rect 817 327 958 332
rect 161 322 222 327
rect 241 322 590 327
rect 737 322 822 327
rect 953 322 982 327
rect 1113 322 1190 327
rect 1209 322 1318 327
rect 1553 322 1558 342
rect 1617 332 1670 337
rect 1985 332 2086 337
rect 2289 332 2334 337
rect 2425 332 2446 337
rect 2577 332 2614 337
rect 2633 332 2678 337
rect 2729 332 2790 337
rect 2985 332 3030 337
rect 3089 332 3350 337
rect 3505 332 3582 337
rect 3681 332 3814 337
rect 3865 332 4038 337
rect 1689 327 1782 332
rect 1569 322 1694 327
rect 1777 322 1806 327
rect 1841 322 1902 327
rect 1921 322 1958 327
rect 2009 322 2142 327
rect 2161 322 2270 327
rect 2297 322 2326 327
rect 2441 322 2446 332
rect 3025 327 3094 332
rect 2465 322 2742 327
rect 2937 322 3006 327
rect 3225 322 3262 327
rect 3545 322 3862 327
rect 3897 322 3926 327
rect 4001 322 4046 327
rect 1001 317 1094 322
rect 1569 317 1574 322
rect 153 312 214 317
rect 225 312 286 317
rect 601 312 726 317
rect 833 312 1006 317
rect 1089 312 1134 317
rect 1177 312 1230 317
rect 1329 312 1406 317
rect 1481 312 1526 317
rect 1545 312 1574 317
rect 1649 312 1694 317
rect 1705 312 1750 317
rect 1801 312 1846 317
rect 1857 312 1862 322
rect 2161 317 2166 322
rect 1961 312 2166 317
rect 2265 317 2270 322
rect 4001 317 4006 322
rect 2265 312 2686 317
rect 833 307 838 312
rect 1225 307 1334 312
rect 2681 307 2686 312
rect 2753 312 2926 317
rect 3009 312 3630 317
rect 3641 312 3782 317
rect 3809 312 4006 317
rect 4025 312 4094 317
rect 2753 307 2758 312
rect 2921 307 3014 312
rect 233 302 262 307
rect 273 302 518 307
rect 593 302 630 307
rect 721 302 838 307
rect 857 302 1062 307
rect 1073 302 1150 307
rect 1169 302 1206 307
rect 1353 302 1398 307
rect 1481 302 2406 307
rect 2417 302 2454 307
rect 2529 302 2574 307
rect 2617 302 2662 307
rect 2681 302 2758 307
rect 3033 302 3070 307
rect 3545 302 3582 307
rect 3649 302 3686 307
rect 3801 302 3846 307
rect 3905 302 3982 307
rect 3089 297 3206 302
rect 3249 297 3398 302
rect 209 292 238 297
rect 465 292 998 297
rect 1121 292 1190 297
rect 1249 292 1758 297
rect 1793 292 1894 297
rect 1953 292 2046 297
rect 2057 292 2118 297
rect 2369 292 2470 297
rect 2481 292 2550 297
rect 2897 292 3094 297
rect 3201 292 3254 297
rect 3393 292 3462 297
rect 3497 292 3670 297
rect 233 287 238 292
rect 337 287 470 292
rect 2137 287 2350 292
rect 2569 287 2662 292
rect 233 282 342 287
rect 489 282 742 287
rect 785 282 1110 287
rect 1137 282 1174 287
rect 1561 282 1958 287
rect 2025 282 2142 287
rect 2345 282 2382 287
rect 2481 282 2574 287
rect 2657 282 3382 287
rect 3505 282 3534 287
rect 737 277 742 282
rect 1193 277 1374 282
rect 1425 277 1566 282
rect 2377 277 2486 282
rect 3377 277 3510 282
rect 361 272 430 277
rect 449 272 726 277
rect 737 272 1198 277
rect 1369 272 1398 277
rect 361 267 366 272
rect 281 262 366 267
rect 425 267 430 272
rect 1425 267 1430 277
rect 1585 272 1742 277
rect 1753 272 1830 277
rect 1841 272 1918 277
rect 2001 272 2358 277
rect 2505 272 2646 277
rect 2641 267 2646 272
rect 2937 272 3190 277
rect 3281 272 3358 277
rect 3561 272 3902 277
rect 2937 267 2942 272
rect 425 262 1006 267
rect 1057 262 1430 267
rect 1441 262 1550 267
rect 1609 262 1766 267
rect 1785 262 1814 267
rect 1865 262 1950 267
rect 1961 262 2022 267
rect 2089 262 2318 267
rect 2401 262 2622 267
rect 2641 262 2942 267
rect 2961 262 3414 267
rect 3513 262 3566 267
rect 3873 262 3910 267
rect 1441 257 1446 262
rect 377 252 454 257
rect 521 252 662 257
rect 745 252 926 257
rect 1009 252 1046 257
rect 1161 252 1190 257
rect 1233 252 1382 257
rect 1393 252 1446 257
rect 1529 252 1750 257
rect 1777 252 2614 257
rect 3065 252 3310 257
rect 3457 252 3670 257
rect 3689 252 3710 257
rect 3833 252 3886 257
rect 657 247 750 252
rect 1041 247 1166 252
rect 1377 247 1382 252
rect 2633 247 2702 252
rect 2961 247 3046 252
rect 409 242 638 247
rect 769 242 854 247
rect 929 242 1022 247
rect 1281 242 1358 247
rect 1377 242 2054 247
rect 2073 242 2638 247
rect 2697 242 2966 247
rect 3041 242 3478 247
rect 3561 242 3702 247
rect 3761 242 3838 247
rect 1281 237 1286 242
rect 425 232 534 237
rect 561 232 630 237
rect 761 232 1054 237
rect 1089 232 1142 237
rect 1225 232 1286 237
rect 1353 232 1390 237
rect 1465 232 1606 237
rect 1641 232 1782 237
rect 1801 232 2638 237
rect 2657 232 2686 237
rect 2977 232 3006 237
rect 3017 232 3350 237
rect 3489 232 3822 237
rect 3905 232 3966 237
rect 561 227 566 232
rect 3345 227 3478 232
rect 3905 227 3910 232
rect 249 222 566 227
rect 577 222 614 227
rect 633 222 1582 227
rect 1681 222 2070 227
rect 2113 222 2310 227
rect 2393 222 2478 227
rect 2537 222 2590 227
rect 2641 222 2726 227
rect 2753 222 2798 227
rect 2873 222 3254 227
rect 3265 222 3318 227
rect 3473 222 3638 227
rect 3713 222 3742 227
rect 3785 222 3830 227
rect 3849 222 3910 227
rect 3921 222 3974 227
rect 4033 222 4086 227
rect 1601 217 1686 222
rect 3249 217 3254 222
rect 3633 217 3638 222
rect 217 212 606 217
rect 729 212 934 217
rect 969 212 1054 217
rect 1065 212 1126 217
rect 1161 212 1294 217
rect 1393 212 1606 217
rect 1705 212 1806 217
rect 1841 212 1926 217
rect 1937 212 2046 217
rect 2073 212 2294 217
rect 2417 212 2446 217
rect 2553 212 2582 217
rect 2705 212 2742 217
rect 3025 212 3054 217
rect 3129 212 3238 217
rect 3249 212 3502 217
rect 3553 212 3574 217
rect 3633 212 3726 217
rect 3825 212 4046 217
rect 1393 207 1398 212
rect 2441 207 2558 212
rect 2577 207 2582 212
rect 425 202 702 207
rect 713 202 782 207
rect 873 202 1110 207
rect 1281 202 1398 207
rect 1433 202 1798 207
rect 1889 202 2302 207
rect 2313 202 2334 207
rect 2577 202 2694 207
rect 2809 202 2894 207
rect 3233 202 3238 212
rect 3569 207 3574 212
rect 3361 202 3486 207
rect 3529 202 3694 207
rect 3745 202 3854 207
rect 3881 202 3926 207
rect 4017 202 4038 207
rect 1793 197 1894 202
rect 3233 197 3342 202
rect 113 192 190 197
rect 345 192 374 197
rect 457 192 510 197
rect 529 192 558 197
rect 113 187 118 192
rect 73 182 118 187
rect 185 187 190 192
rect 553 187 558 192
rect 633 192 670 197
rect 681 192 742 197
rect 865 192 894 197
rect 993 192 1030 197
rect 1089 192 1174 197
rect 1185 192 1486 197
rect 1497 192 1590 197
rect 1665 192 1710 197
rect 1737 192 1774 197
rect 1913 192 1950 197
rect 2033 192 2094 197
rect 2169 192 2230 197
rect 2409 192 2430 197
rect 2489 192 2566 197
rect 2633 192 2662 197
rect 2721 192 2758 197
rect 2865 192 3022 197
rect 3049 192 3118 197
rect 3145 192 3206 197
rect 3337 192 3510 197
rect 3769 192 3870 197
rect 3897 192 4014 197
rect 633 187 638 192
rect 2561 187 2638 192
rect 185 182 238 187
rect 553 182 638 187
rect 657 182 886 187
rect 1121 182 1246 187
rect 1577 182 1718 187
rect 1793 182 1838 187
rect 1929 182 2022 187
rect 2049 182 2118 187
rect 2145 182 2206 187
rect 2417 182 2454 187
rect 2897 182 3134 187
rect 3161 182 3334 187
rect 3345 182 3678 187
rect 1265 177 1430 182
rect 3673 177 3678 182
rect 3889 182 3974 187
rect 3889 177 3894 182
rect 129 172 174 177
rect 665 172 830 177
rect 825 167 830 172
rect 897 172 1158 177
rect 1169 172 1270 177
rect 1425 172 1454 177
rect 1617 172 1734 177
rect 1753 172 2078 177
rect 2137 172 2246 177
rect 2545 172 2694 177
rect 2969 172 3070 177
rect 3185 172 3278 177
rect 3321 172 3398 177
rect 3505 172 3534 177
rect 3673 172 3894 177
rect 897 167 902 172
rect 1153 167 1158 172
rect 1729 167 1734 172
rect 2545 167 2550 172
rect 593 162 654 167
rect 777 162 806 167
rect 825 162 902 167
rect 1073 162 1134 167
rect 1153 162 1614 167
rect 1625 162 1662 167
rect 1729 162 1990 167
rect 2001 162 2118 167
rect 2129 162 2174 167
rect 2201 162 2262 167
rect 2281 162 2502 167
rect 2521 162 2550 167
rect 2689 167 2694 172
rect 3393 167 3510 172
rect 2689 162 2862 167
rect 2913 162 2942 167
rect 3001 162 3062 167
rect 3073 162 3342 167
rect 649 157 782 162
rect 2281 157 2286 162
rect 1129 152 1182 157
rect 1265 152 1398 157
rect 1617 152 2286 157
rect 2497 157 2502 162
rect 2497 152 2678 157
rect 3073 152 3078 162
rect 3329 152 3654 157
rect 3913 152 3950 157
rect 2817 147 3078 152
rect 3649 147 3654 152
rect 153 142 566 147
rect 665 142 982 147
rect 1153 142 1190 147
rect 1201 142 1342 147
rect 1409 142 2822 147
rect 3249 142 3318 147
rect 801 132 830 137
rect 825 127 830 132
rect 993 132 1174 137
rect 993 127 998 132
rect 825 122 998 127
rect 1185 127 1190 142
rect 1337 137 1414 142
rect 3249 137 3254 142
rect 3313 137 3318 142
rect 3473 142 3502 147
rect 3649 142 3702 147
rect 3809 142 4038 147
rect 3473 137 3478 142
rect 1273 132 1318 137
rect 1633 127 1638 137
rect 1681 132 1878 137
rect 2097 132 2742 137
rect 2833 132 3254 137
rect 3265 132 3294 137
rect 3313 132 3478 137
rect 3505 132 3542 137
rect 3953 132 4062 137
rect 4081 132 4118 137
rect 1897 127 1974 132
rect 2737 127 2838 132
rect 1185 122 1294 127
rect 1417 122 1518 127
rect 1633 122 1902 127
rect 1969 122 2494 127
rect 2545 122 2598 127
rect 2593 117 2598 122
rect 2689 122 2718 127
rect 2857 122 2990 127
rect 2689 117 2694 122
rect 2985 117 2990 122
rect 3073 122 3102 127
rect 3073 117 3078 122
rect 225 112 270 117
rect 345 112 390 117
rect 513 112 790 117
rect 785 107 790 112
rect 1425 112 1622 117
rect 1633 112 1678 117
rect 1793 112 1838 117
rect 1913 112 1958 117
rect 2033 112 2078 117
rect 2121 112 2150 117
rect 2273 112 2526 117
rect 2593 112 2694 117
rect 2745 112 2790 117
rect 2985 112 3078 117
rect 785 102 1174 107
rect 1169 97 1174 102
rect 1425 97 1430 112
rect 2145 107 2278 112
rect 1449 102 1478 107
rect 1169 92 1430 97
rect 1473 97 1478 102
rect 1657 102 1686 107
rect 1721 102 1902 107
rect 1657 97 1662 102
rect 1473 92 1662 97
rect 1897 97 1902 102
rect 1969 102 1990 107
rect 2297 102 2574 107
rect 1969 97 1974 102
rect 1897 92 1974 97
rect 1985 97 1990 102
rect 2569 97 2574 102
rect 2801 102 2846 107
rect 2801 97 2806 102
rect 1985 92 2286 97
rect 2281 87 2286 92
rect 2521 92 2550 97
rect 2569 92 2806 97
rect 2841 97 2846 102
rect 3113 102 3622 107
rect 3113 97 3118 102
rect 2841 92 3118 97
rect 2521 87 2526 92
rect 2281 82 2526 87
rect 1585 72 1966 77
rect 1585 57 1590 72
rect 1961 67 1966 72
rect 1961 62 2382 67
rect 289 52 1590 57
rect 2377 57 2382 62
rect 2401 57 2406 67
rect 2377 52 2406 57
rect 1601 42 2694 47
rect 1745 22 1774 27
rect 1769 17 1774 22
rect 2705 22 2742 27
rect 2705 17 2710 22
rect 1769 12 2710 17
use top_level_VIA1  top_level_VIA1_0
timestamp 1682952543
transform 1 0 24 0 1 4117
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_1
timestamp 1682952543
transform 1 0 4201 0 1 4117
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_2
timestamp 1682952543
transform 1 0 48 0 1 4093
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_3
timestamp 1682952543
transform 1 0 4177 0 1 4093
box -10 -10 10 10
use top_level_VIA0  top_level_VIA0_0
timestamp 1682952543
transform 1 0 24 0 1 4070
box -10 -3 10 3
use M2_M1  M2_M1_0
timestamp 1682952543
transform 1 0 132 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1
timestamp 1682952543
transform 1 0 164 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1682952543
transform 1 0 172 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1682952543
transform 1 0 188 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1682952543
transform 1 0 84 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_46
timestamp 1682952543
transform 1 0 132 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_47
timestamp 1682952543
transform 1 0 172 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_91
timestamp 1682952543
transform 1 0 180 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1682952543
transform 1 0 164 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1682952543
transform 1 0 180 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_92
timestamp 1682952543
transform 1 0 220 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1682952543
transform 1 0 236 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1682952543
transform 1 0 236 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1682952543
transform 1 0 252 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1682952543
transform 1 0 292 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1682952543
transform 1 0 252 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_6
timestamp 1682952543
transform 1 0 292 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1682952543
transform 1 0 348 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1682952543
transform 1 0 244 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_61
timestamp 1682952543
transform 1 0 244 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_94
timestamp 1682952543
transform 1 0 268 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1682952543
transform 1 0 340 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_62
timestamp 1682952543
transform 1 0 300 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_95
timestamp 1682952543
transform 1 0 372 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_10
timestamp 1682952543
transform 1 0 396 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_8
timestamp 1682952543
transform 1 0 396 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_11
timestamp 1682952543
transform 1 0 436 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1682952543
transform 1 0 436 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1682952543
transform 1 0 492 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1682952543
transform 1 0 412 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_101
timestamp 1682952543
transform 1 0 436 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1682952543
transform 1 0 516 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1682952543
transform 1 0 556 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1682952543
transform 1 0 516 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_12
timestamp 1682952543
transform 1 0 556 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_13
timestamp 1682952543
transform 1 0 612 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1682952543
transform 1 0 508 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1682952543
transform 1 0 532 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_63
timestamp 1682952543
transform 1 0 532 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_14
timestamp 1682952543
transform 1 0 676 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1682952543
transform 1 0 716 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1682952543
transform 1 0 636 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_64
timestamp 1682952543
transform 1 0 636 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_16
timestamp 1682952543
transform 1 0 732 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_17
timestamp 1682952543
transform 1 0 780 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1682952543
transform 1 0 812 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_65
timestamp 1682952543
transform 1 0 812 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_101
timestamp 1682952543
transform 1 0 836 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_14
timestamp 1682952543
transform 1 0 852 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1682952543
transform 1 0 892 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_18
timestamp 1682952543
transform 1 0 852 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_19
timestamp 1682952543
transform 1 0 860 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1682952543
transform 1 0 892 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_50
timestamp 1682952543
transform 1 0 916 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_102
timestamp 1682952543
transform 1 0 940 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_66
timestamp 1682952543
transform 1 0 876 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1682952543
transform 1 0 940 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1682952543
transform 1 0 956 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_51
timestamp 1682952543
transform 1 0 956 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_22
timestamp 1682952543
transform 1 0 996 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_103
timestamp 1682952543
transform 1 0 1044 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_68
timestamp 1682952543
transform 1 0 1044 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_23
timestamp 1682952543
transform 1 0 1100 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1682952543
transform 1 0 1156 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1682952543
transform 1 0 1076 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_102
timestamp 1682952543
transform 1 0 1076 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1682952543
transform 1 0 1180 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1682952543
transform 1 0 1220 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_18
timestamp 1682952543
transform 1 0 1292 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1682952543
transform 1 0 1332 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_25
timestamp 1682952543
transform 1 0 1180 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1682952543
transform 1 0 1220 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1682952543
transform 1 0 1276 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1682952543
transform 1 0 1292 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_29
timestamp 1682952543
transform 1 0 1300 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1682952543
transform 1 0 1332 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1682952543
transform 1 0 1396 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1682952543
transform 1 0 1452 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1682952543
transform 1 0 1172 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_69
timestamp 1682952543
transform 1 0 1172 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_106
timestamp 1682952543
transform 1 0 1196 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1682952543
transform 1 0 1284 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_70
timestamp 1682952543
transform 1 0 1220 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1682952543
transform 1 0 1196 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_108
timestamp 1682952543
transform 1 0 1380 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_71
timestamp 1682952543
transform 1 0 1380 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_109
timestamp 1682952543
transform 1 0 1476 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_72
timestamp 1682952543
transform 1 0 1460 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1682952543
transform 1 0 1476 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1682952543
transform 1 0 1548 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1682952543
transform 1 0 1588 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_33
timestamp 1682952543
transform 1 0 1548 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1682952543
transform 1 0 1580 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1682952543
transform 1 0 1588 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_110
timestamp 1682952543
transform 1 0 1500 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_74
timestamp 1682952543
transform 1 0 1500 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_111
timestamp 1682952543
transform 1 0 1604 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1682952543
transform 1 0 1644 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_22
timestamp 1682952543
transform 1 0 1660 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1682952543
transform 1 0 1700 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_36
timestamp 1682952543
transform 1 0 1660 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1682952543
transform 1 0 1668 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1682952543
transform 1 0 1700 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1682952543
transform 1 0 1748 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_75
timestamp 1682952543
transform 1 0 1748 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_39
timestamp 1682952543
transform 1 0 1764 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1682952543
transform 1 0 1772 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_40
timestamp 1682952543
transform 1 0 1836 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_36
timestamp 1682952543
transform 1 0 1860 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_114
timestamp 1682952543
transform 1 0 1860 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1682952543
transform 1 0 1860 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1682952543
transform 1 0 1972 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_41
timestamp 1682952543
transform 1 0 1884 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_37
timestamp 1682952543
transform 1 0 1892 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_42
timestamp 1682952543
transform 1 0 1940 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1682952543
transform 1 0 1964 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_78
timestamp 1682952543
transform 1 0 1964 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1682952543
transform 1 0 2004 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1682952543
transform 1 0 2028 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1682952543
transform 1 0 2020 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1682952543
transform 1 0 2020 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1682952543
transform 1 0 2020 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1682952543
transform 1 0 2076 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1682952543
transform 1 0 1996 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_79
timestamp 1682952543
transform 1 0 1996 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1682952543
transform 1 0 2164 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1682952543
transform 1 0 2100 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_45
timestamp 1682952543
transform 1 0 2124 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_39
timestamp 1682952543
transform 1 0 2140 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_46
timestamp 1682952543
transform 1 0 2180 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1682952543
transform 1 0 2188 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1682952543
transform 1 0 2204 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1682952543
transform 1 0 2236 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_117
timestamp 1682952543
transform 1 0 2100 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_80
timestamp 1682952543
transform 1 0 2100 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_118
timestamp 1682952543
transform 1 0 2196 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_52
timestamp 1682952543
transform 1 0 2204 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1682952543
transform 1 0 2244 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_119
timestamp 1682952543
transform 1 0 2284 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_50
timestamp 1682952543
transform 1 0 2364 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1682952543
transform 1 0 2316 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_81
timestamp 1682952543
transform 1 0 2316 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1682952543
transform 1 0 2340 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1682952543
transform 1 0 2364 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_51
timestamp 1682952543
transform 1 0 2420 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_84
timestamp 1682952543
transform 1 0 2428 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_104
timestamp 1682952543
transform 1 0 2420 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_52
timestamp 1682952543
transform 1 0 2484 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1682952543
transform 1 0 2444 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1682952543
transform 1 0 2436 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_53
timestamp 1682952543
transform 1 0 2532 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1682952543
transform 1 0 2612 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_40
timestamp 1682952543
transform 1 0 2660 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_55
timestamp 1682952543
transform 1 0 2668 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1682952543
transform 1 0 2588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_24
timestamp 1682952543
transform 1 0 2692 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_123
timestamp 1682952543
transform 1 0 2684 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_124
timestamp 1682952543
transform 1 0 2692 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_25
timestamp 1682952543
transform 1 0 2724 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_56
timestamp 1682952543
transform 1 0 2700 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_57
timestamp 1682952543
transform 1 0 2708 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1682952543
transform 1 0 2724 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1682952543
transform 1 0 2780 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_41
timestamp 1682952543
transform 1 0 2804 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_54
timestamp 1682952543
transform 1 0 2740 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_125
timestamp 1682952543
transform 1 0 2804 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_85
timestamp 1682952543
transform 1 0 2780 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1682952543
transform 1 0 2804 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_26
timestamp 1682952543
transform 1 0 2820 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_126
timestamp 1682952543
transform 1 0 2820 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_27
timestamp 1682952543
transform 1 0 2852 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_60
timestamp 1682952543
transform 1 0 2836 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1682952543
transform 1 0 2852 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1682952543
transform 1 0 2884 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1682952543
transform 1 0 2932 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_55
timestamp 1682952543
transform 1 0 2844 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1682952543
transform 1 0 2884 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_127
timestamp 1682952543
transform 1 0 2932 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1682952543
transform 1 0 2836 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1682952543
transform 1 0 2852 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1682952543
transform 1 0 2948 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_63
timestamp 1682952543
transform 1 0 2964 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_29
timestamp 1682952543
transform 1 0 2980 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_64
timestamp 1682952543
transform 1 0 2980 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_57
timestamp 1682952543
transform 1 0 2972 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_65
timestamp 1682952543
transform 1 0 3028 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_43
timestamp 1682952543
transform 1 0 3076 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1682952543
transform 1 0 3028 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_128
timestamp 1682952543
transform 1 0 3076 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_66
timestamp 1682952543
transform 1 0 3100 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1682952543
transform 1 0 3116 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_59
timestamp 1682952543
transform 1 0 3108 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_68
timestamp 1682952543
transform 1 0 3164 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1682952543
transform 1 0 3212 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1682952543
transform 1 0 3164 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_129
timestamp 1682952543
transform 1 0 3212 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_0
timestamp 1682952543
transform 1 0 3308 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1682952543
transform 1 0 3332 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1682952543
transform 1 0 3284 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1682952543
transform 1 0 3340 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1682952543
transform 1 0 3252 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_69
timestamp 1682952543
transform 1 0 3276 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_70
timestamp 1682952543
transform 1 0 3332 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1682952543
transform 1 0 3340 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1682952543
transform 1 0 3252 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_89
timestamp 1682952543
transform 1 0 3268 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1682952543
transform 1 0 3284 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1682952543
transform 1 0 3300 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1682952543
transform 1 0 3252 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1682952543
transform 1 0 3356 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_131
timestamp 1682952543
transform 1 0 3348 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_33
timestamp 1682952543
transform 1 0 3460 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_72
timestamp 1682952543
transform 1 0 3396 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1682952543
transform 1 0 3452 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1682952543
transform 1 0 3460 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1682952543
transform 1 0 3372 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_92
timestamp 1682952543
transform 1 0 3372 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_133
timestamp 1682952543
transform 1 0 3468 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_107
timestamp 1682952543
transform 1 0 3452 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1682952543
transform 1 0 3780 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_75
timestamp 1682952543
transform 1 0 3532 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1682952543
transform 1 0 3572 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_77
timestamp 1682952543
transform 1 0 3636 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1682952543
transform 1 0 3668 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1682952543
transform 1 0 3708 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1682952543
transform 1 0 3764 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1682952543
transform 1 0 3828 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_82
timestamp 1682952543
transform 1 0 3860 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1682952543
transform 1 0 3492 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_93
timestamp 1682952543
transform 1 0 3492 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1682952543
transform 1 0 3492 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_135
timestamp 1682952543
transform 1 0 3588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_109
timestamp 1682952543
transform 1 0 3588 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_136
timestamp 1682952543
transform 1 0 3684 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_110
timestamp 1682952543
transform 1 0 3684 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1682952543
transform 1 0 3748 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_137
timestamp 1682952543
transform 1 0 3780 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1682952543
transform 1 0 3884 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1682952543
transform 1 0 3876 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1682952543
transform 1 0 3780 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1682952543
transform 1 0 3828 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1682952543
transform 1 0 3868 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1682952543
transform 1 0 3900 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_84
timestamp 1682952543
transform 1 0 3924 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1682952543
transform 1 0 3980 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1682952543
transform 1 0 3988 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1682952543
transform 1 0 3900 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1682952543
transform 1 0 4036 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_88
timestamp 1682952543
transform 1 0 4092 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1682952543
transform 1 0 3996 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1682952543
transform 1 0 4012 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_97
timestamp 1682952543
transform 1 0 3996 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1682952543
transform 1 0 4036 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1682952543
transform 1 0 3980 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_113
timestamp 1682952543
transform 1 0 4012 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_89
timestamp 1682952543
transform 1 0 4116 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1682952543
transform 1 0 4108 0 1 4005
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_1
timestamp 1682952543
transform 1 0 4201 0 1 4070
box -10 -3 10 3
use top_level_VIA0  top_level_VIA0_2
timestamp 1682952543
transform 1 0 48 0 1 3970
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_0
timestamp 1682952543
transform 1 0 72 0 1 3970
box -8 -3 104 105
use AOI22X1  AOI22X1_0
timestamp 1682952543
transform -1 0 208 0 1 3970
box -8 -3 46 105
use FILL  FILL_0
timestamp 1682952543
transform 1 0 208 0 1 3970
box -8 -3 16 105
use FILL  FILL_1
timestamp 1682952543
transform 1 0 216 0 1 3970
box -8 -3 16 105
use FILL  FILL_2
timestamp 1682952543
transform 1 0 224 0 1 3970
box -8 -3 16 105
use FILL  FILL_3
timestamp 1682952543
transform 1 0 232 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_114
timestamp 1682952543
transform 1 0 268 0 1 3975
box -3 -3 3 3
use INVX2  INVX2_0
timestamp 1682952543
transform 1 0 240 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1682952543
transform 1 0 256 0 1 3970
box -8 -3 104 105
use FILL  FILL_4
timestamp 1682952543
transform 1 0 352 0 1 3970
box -8 -3 16 105
use FILL  FILL_5
timestamp 1682952543
transform 1 0 360 0 1 3970
box -8 -3 16 105
use FILL  FILL_6
timestamp 1682952543
transform 1 0 368 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_1
timestamp 1682952543
transform 1 0 376 0 1 3970
box -9 -3 26 105
use FILL  FILL_7
timestamp 1682952543
transform 1 0 392 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_115
timestamp 1682952543
transform 1 0 412 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_2
timestamp 1682952543
transform 1 0 400 0 1 3970
box -8 -3 104 105
use FILL  FILL_8
timestamp 1682952543
transform 1 0 496 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1682952543
transform 1 0 504 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1682952543
transform 1 0 520 0 1 3970
box -8 -3 104 105
use FILL  FILL_9
timestamp 1682952543
transform 1 0 616 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_116
timestamp 1682952543
transform 1 0 716 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_4
timestamp 1682952543
transform 1 0 624 0 1 3970
box -8 -3 104 105
use FILL  FILL_10
timestamp 1682952543
transform 1 0 720 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1682952543
transform -1 0 824 0 1 3970
box -8 -3 104 105
use FILL  FILL_11
timestamp 1682952543
transform 1 0 824 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_117
timestamp 1682952543
transform 1 0 860 0 1 3975
box -3 -3 3 3
use INVX2  INVX2_3
timestamp 1682952543
transform 1 0 832 0 1 3970
box -9 -3 26 105
use FILL  FILL_12
timestamp 1682952543
transform 1 0 848 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1682952543
transform -1 0 952 0 1 3970
box -8 -3 104 105
use FILL  FILL_13
timestamp 1682952543
transform 1 0 952 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1682952543
transform -1 0 1056 0 1 3970
box -8 -3 104 105
use FILL  FILL_14
timestamp 1682952543
transform 1 0 1056 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1682952543
transform 1 0 1064 0 1 3970
box -8 -3 104 105
use FILL  FILL_15
timestamp 1682952543
transform 1 0 1160 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_4
timestamp 1682952543
transform 1 0 1168 0 1 3970
box -9 -3 26 105
use M3_M2  M3_M2_118
timestamp 1682952543
transform 1 0 1284 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_9
timestamp 1682952543
transform 1 0 1184 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_5
timestamp 1682952543
transform 1 0 1280 0 1 3970
box -9 -3 26 105
use M3_M2  M3_M2_119
timestamp 1682952543
transform 1 0 1324 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_10
timestamp 1682952543
transform -1 0 1392 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1682952543
transform -1 0 1488 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1682952543
transform 1 0 1488 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_6
timestamp 1682952543
transform -1 0 1600 0 1 3970
box -9 -3 26 105
use FILL  FILL_16
timestamp 1682952543
transform 1 0 1600 0 1 3970
box -8 -3 16 105
use FILL  FILL_17
timestamp 1682952543
transform 1 0 1608 0 1 3970
box -8 -3 16 105
use FILL  FILL_18
timestamp 1682952543
transform 1 0 1616 0 1 3970
box -8 -3 16 105
use FILL  FILL_19
timestamp 1682952543
transform 1 0 1624 0 1 3970
box -8 -3 16 105
use FILL  FILL_20
timestamp 1682952543
transform 1 0 1632 0 1 3970
box -8 -3 16 105
use FILL  FILL_21
timestamp 1682952543
transform 1 0 1640 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_7
timestamp 1682952543
transform 1 0 1648 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1682952543
transform -1 0 1760 0 1 3970
box -8 -3 104 105
use FILL  FILL_22
timestamp 1682952543
transform 1 0 1760 0 1 3970
box -8 -3 16 105
use FILL  FILL_23
timestamp 1682952543
transform 1 0 1768 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_120
timestamp 1682952543
transform 1 0 1852 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_14
timestamp 1682952543
transform -1 0 1872 0 1 3970
box -8 -3 104 105
use M3_M2  M3_M2_121
timestamp 1682952543
transform 1 0 1884 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_122
timestamp 1682952543
transform 1 0 1916 0 1 3975
box -3 -3 3 3
use FILL  FILL_24
timestamp 1682952543
transform 1 0 1872 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_123
timestamp 1682952543
transform 1 0 1956 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_15
timestamp 1682952543
transform -1 0 1976 0 1 3970
box -8 -3 104 105
use FILL  FILL_25
timestamp 1682952543
transform 1 0 1976 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1682952543
transform 1 0 1984 0 1 3970
box -8 -3 104 105
use FILL  FILL_26
timestamp 1682952543
transform 1 0 2080 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1682952543
transform 1 0 2088 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_8
timestamp 1682952543
transform -1 0 2200 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1682952543
transform -1 0 2296 0 1 3970
box -8 -3 104 105
use FILL  FILL_27
timestamp 1682952543
transform 1 0 2296 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_124
timestamp 1682952543
transform 1 0 2340 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_19
timestamp 1682952543
transform 1 0 2304 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_9
timestamp 1682952543
transform 1 0 2400 0 1 3970
box -9 -3 26 105
use FILL  FILL_28
timestamp 1682952543
transform 1 0 2416 0 1 3970
box -8 -3 16 105
use FILL  FILL_29
timestamp 1682952543
transform 1 0 2424 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_125
timestamp 1682952543
transform 1 0 2444 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_20
timestamp 1682952543
transform 1 0 2432 0 1 3970
box -8 -3 104 105
use FILL  FILL_30
timestamp 1682952543
transform 1 0 2528 0 1 3970
box -8 -3 16 105
use FILL  FILL_76
timestamp 1682952543
transform 1 0 2536 0 1 3970
box -8 -3 16 105
use FILL  FILL_77
timestamp 1682952543
transform 1 0 2544 0 1 3970
box -8 -3 16 105
use FILL  FILL_78
timestamp 1682952543
transform 1 0 2552 0 1 3970
box -8 -3 16 105
use FILL  FILL_80
timestamp 1682952543
transform 1 0 2560 0 1 3970
box -8 -3 16 105
use FILL  FILL_82
timestamp 1682952543
transform 1 0 2568 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_126
timestamp 1682952543
transform 1 0 2588 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_28
timestamp 1682952543
transform 1 0 2576 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_21
timestamp 1682952543
transform -1 0 2688 0 1 3970
box -9 -3 26 105
use FILL  FILL_83
timestamp 1682952543
transform 1 0 2688 0 1 3970
box -8 -3 16 105
use FILL  FILL_84
timestamp 1682952543
transform 1 0 2696 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_22
timestamp 1682952543
transform 1 0 2704 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1682952543
transform -1 0 2816 0 1 3970
box -8 -3 104 105
use M3_M2  M3_M2_127
timestamp 1682952543
transform 1 0 2828 0 1 3975
box -3 -3 3 3
use FILL  FILL_85
timestamp 1682952543
transform 1 0 2816 0 1 3970
box -8 -3 16 105
use FILL  FILL_86
timestamp 1682952543
transform 1 0 2824 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_23
timestamp 1682952543
transform 1 0 2832 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1682952543
transform -1 0 2944 0 1 3970
box -8 -3 104 105
use FILL  FILL_87
timestamp 1682952543
transform 1 0 2944 0 1 3970
box -8 -3 16 105
use FILL  FILL_95
timestamp 1682952543
transform 1 0 2952 0 1 3970
box -8 -3 16 105
use FILL  FILL_96
timestamp 1682952543
transform 1 0 2960 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_128
timestamp 1682952543
transform 1 0 2988 0 1 3975
box -3 -3 3 3
use INVX2  INVX2_26
timestamp 1682952543
transform -1 0 2984 0 1 3970
box -9 -3 26 105
use FILL  FILL_97
timestamp 1682952543
transform 1 0 2984 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_129
timestamp 1682952543
transform 1 0 3092 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_32
timestamp 1682952543
transform -1 0 3088 0 1 3970
box -8 -3 104 105
use FILL  FILL_98
timestamp 1682952543
transform 1 0 3088 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_27
timestamp 1682952543
transform -1 0 3112 0 1 3970
box -9 -3 26 105
use FILL  FILL_99
timestamp 1682952543
transform 1 0 3112 0 1 3970
box -8 -3 16 105
use FILL  FILL_100
timestamp 1682952543
transform 1 0 3120 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1682952543
transform -1 0 3224 0 1 3970
box -8 -3 104 105
use FILL  FILL_101
timestamp 1682952543
transform 1 0 3224 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_130
timestamp 1682952543
transform 1 0 3244 0 1 3975
box -3 -3 3 3
use FILL  FILL_102
timestamp 1682952543
transform 1 0 3232 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_131
timestamp 1682952543
transform 1 0 3260 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_34
timestamp 1682952543
transform 1 0 3240 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_28
timestamp 1682952543
transform -1 0 3352 0 1 3970
box -9 -3 26 105
use FILL  FILL_103
timestamp 1682952543
transform 1 0 3352 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1682952543
transform 1 0 3360 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_32
timestamp 1682952543
transform -1 0 3472 0 1 3970
box -9 -3 26 105
use FILL  FILL_105
timestamp 1682952543
transform 1 0 3472 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_132
timestamp 1682952543
transform 1 0 3548 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_38
timestamp 1682952543
transform 1 0 3480 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1682952543
transform 1 0 3576 0 1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1682952543
transform 1 0 3672 0 1 3970
box -8 -3 104 105
use M3_M2  M3_M2_133
timestamp 1682952543
transform 1 0 3852 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_41
timestamp 1682952543
transform 1 0 3768 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_33
timestamp 1682952543
transform -1 0 3880 0 1 3970
box -9 -3 26 105
use M3_M2  M3_M2_134
timestamp 1682952543
transform 1 0 3892 0 1 3975
box -3 -3 3 3
use FILL  FILL_106
timestamp 1682952543
transform 1 0 3880 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1682952543
transform 1 0 3888 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_34
timestamp 1682952543
transform -1 0 4000 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1682952543
transform 1 0 4000 0 1 3970
box -8 -3 104 105
use INVX2  INVX2_35
timestamp 1682952543
transform -1 0 4112 0 1 3970
box -9 -3 26 105
use FILL  FILL_107
timestamp 1682952543
transform 1 0 4112 0 1 3970
box -8 -3 16 105
use FILL  FILL_108
timestamp 1682952543
transform 1 0 4120 0 1 3970
box -8 -3 16 105
use FILL  FILL_109
timestamp 1682952543
transform 1 0 4128 0 1 3970
box -8 -3 16 105
use FILL  FILL_110
timestamp 1682952543
transform 1 0 4136 0 1 3970
box -8 -3 16 105
use FILL  FILL_111
timestamp 1682952543
transform 1 0 4144 0 1 3970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_3
timestamp 1682952543
transform 1 0 4177 0 1 3970
box -10 -3 10 3
use M3_M2  M3_M2_183
timestamp 1682952543
transform 1 0 84 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_146
timestamp 1682952543
transform 1 0 84 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_184
timestamp 1682952543
transform 1 0 196 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_147
timestamp 1682952543
transform 1 0 180 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1682952543
transform 1 0 196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1682952543
transform 1 0 116 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1682952543
transform 1 0 164 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1682952543
transform 1 0 172 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_185
timestamp 1682952543
transform 1 0 292 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_149
timestamp 1682952543
transform 1 0 292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1682952543
transform 1 0 228 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1682952543
transform 1 0 276 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1682952543
transform 1 0 284 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1682952543
transform 1 0 300 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_272
timestamp 1682952543
transform 1 0 276 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_273
timestamp 1682952543
transform 1 0 308 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_314
timestamp 1682952543
transform 1 0 324 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_186
timestamp 1682952543
transform 1 0 332 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_311
timestamp 1682952543
transform 1 0 324 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1682952543
transform 1 0 348 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1682952543
transform 1 0 356 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_150
timestamp 1682952543
transform 1 0 348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_151
timestamp 1682952543
transform 1 0 356 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1682952543
transform 1 0 340 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_151
timestamp 1682952543
transform 1 0 388 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1682952543
transform 1 0 428 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_152
timestamp 1682952543
transform 1 0 388 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_153
timestamp 1682952543
transform 1 0 396 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1682952543
transform 1 0 412 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1682952543
transform 1 0 356 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_249
timestamp 1682952543
transform 1 0 364 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_228
timestamp 1682952543
transform 1 0 420 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1682952543
transform 1 0 468 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_155
timestamp 1682952543
transform 1 0 428 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1682952543
transform 1 0 436 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1682952543
transform 1 0 452 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_158
timestamp 1682952543
transform 1 0 468 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1682952543
transform 1 0 372 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1682952543
transform 1 0 388 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1682952543
transform 1 0 404 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1682952543
transform 1 0 420 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_321
timestamp 1682952543
transform 1 0 436 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_322
timestamp 1682952543
transform 1 0 460 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_274
timestamp 1682952543
transform 1 0 396 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1682952543
transform 1 0 420 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1682952543
transform 1 0 468 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_323
timestamp 1682952543
transform 1 0 476 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_276
timestamp 1682952543
transform 1 0 460 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_312
timestamp 1682952543
transform 1 0 364 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_313
timestamp 1682952543
transform 1 0 388 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_314
timestamp 1682952543
transform 1 0 404 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_315
timestamp 1682952543
transform 1 0 436 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1682952543
transform 1 0 452 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1682952543
transform 1 0 492 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1682952543
transform 1 0 500 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_159
timestamp 1682952543
transform 1 0 500 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1682952543
transform 1 0 508 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1682952543
transform 1 0 508 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_324
timestamp 1682952543
transform 1 0 516 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_277
timestamp 1682952543
transform 1 0 508 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1682952543
transform 1 0 556 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_161
timestamp 1682952543
transform 1 0 556 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1682952543
transform 1 0 556 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_326
timestamp 1682952543
transform 1 0 564 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_338
timestamp 1682952543
transform 1 0 556 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_327
timestamp 1682952543
transform 1 0 580 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_339
timestamp 1682952543
transform 1 0 572 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1682952543
transform 1 0 612 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_162
timestamp 1682952543
transform 1 0 596 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1682952543
transform 1 0 604 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1682952543
transform 1 0 620 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_252
timestamp 1682952543
transform 1 0 604 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_328
timestamp 1682952543
transform 1 0 612 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1682952543
transform 1 0 620 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1682952543
transform 1 0 644 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1682952543
transform 1 0 716 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1682952543
transform 1 0 788 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1682952543
transform 1 0 828 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_159
timestamp 1682952543
transform 1 0 852 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1682952543
transform 1 0 820 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1682952543
transform 1 0 884 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_165
timestamp 1682952543
transform 1 0 644 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1682952543
transform 1 0 660 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1682952543
transform 1 0 668 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1682952543
transform 1 0 692 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_169
timestamp 1682952543
transform 1 0 708 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1682952543
transform 1 0 732 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_171
timestamp 1682952543
transform 1 0 756 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1682952543
transform 1 0 764 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1682952543
transform 1 0 788 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1682952543
transform 1 0 804 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_175
timestamp 1682952543
transform 1 0 828 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1682952543
transform 1 0 836 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_177
timestamp 1682952543
transform 1 0 852 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_178
timestamp 1682952543
transform 1 0 860 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_179
timestamp 1682952543
transform 1 0 884 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_329
timestamp 1682952543
transform 1 0 628 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1682952543
transform 1 0 652 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1682952543
transform 1 0 668 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1682952543
transform 1 0 676 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_340
timestamp 1682952543
transform 1 0 628 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1682952543
transform 1 0 692 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_333
timestamp 1682952543
transform 1 0 700 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1682952543
transform 1 0 716 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1682952543
transform 1 0 732 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_278
timestamp 1682952543
transform 1 0 716 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1682952543
transform 1 0 740 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_336
timestamp 1682952543
transform 1 0 748 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1682952543
transform 1 0 764 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_256
timestamp 1682952543
transform 1 0 772 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_338
timestamp 1682952543
transform 1 0 780 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1682952543
transform 1 0 788 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1682952543
transform 1 0 812 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1682952543
transform 1 0 828 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1682952543
transform 1 0 844 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_341
timestamp 1682952543
transform 1 0 700 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1682952543
transform 1 0 732 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1682952543
transform 1 0 756 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1682952543
transform 1 0 812 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_316
timestamp 1682952543
transform 1 0 788 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_344
timestamp 1682952543
transform 1 0 812 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1682952543
transform 1 0 852 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_143
timestamp 1682952543
transform 1 0 964 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1682952543
transform 1 0 916 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1682952543
transform 1 0 932 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1682952543
transform 1 0 940 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_343
timestamp 1682952543
transform 1 0 860 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1682952543
transform 1 0 868 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1682952543
transform 1 0 892 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_258
timestamp 1682952543
transform 1 0 900 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1682952543
transform 1 0 948 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_230
timestamp 1682952543
transform 1 0 964 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_161
timestamp 1682952543
transform 1 0 980 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_144
timestamp 1682952543
transform 1 0 980 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1682952543
transform 1 0 972 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1682952543
transform 1 0 908 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1682952543
transform 1 0 924 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_348
timestamp 1682952543
transform 1 0 940 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_349
timestamp 1682952543
transform 1 0 964 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_280
timestamp 1682952543
transform 1 0 892 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1682952543
transform 1 0 868 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1682952543
transform 1 0 836 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1682952543
transform 1 0 940 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1682952543
transform 1 0 932 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1682952543
transform 1 0 996 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_184
timestamp 1682952543
transform 1 0 1012 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1682952543
transform 1 0 1004 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_347
timestamp 1682952543
transform 1 0 1004 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_190
timestamp 1682952543
transform 1 0 1036 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_185
timestamp 1682952543
transform 1 0 1036 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1682952543
transform 1 0 1052 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1682952543
transform 1 0 1060 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1682952543
transform 1 0 1020 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1682952543
transform 1 0 1028 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1682952543
transform 1 0 1044 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_259
timestamp 1682952543
transform 1 0 1052 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_354
timestamp 1682952543
transform 1 0 1068 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1682952543
transform 1 0 1020 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1682952543
transform 1 0 1028 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1682952543
transform 1 0 1068 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_138
timestamp 1682952543
transform 1 0 1092 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_191
timestamp 1682952543
transform 1 0 1108 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_188
timestamp 1682952543
transform 1 0 1100 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_189
timestamp 1682952543
transform 1 0 1108 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_190
timestamp 1682952543
transform 1 0 1116 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1682952543
transform 1 0 1132 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1682952543
transform 1 0 1148 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1682952543
transform 1 0 1108 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1682952543
transform 1 0 1124 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1682952543
transform 1 0 1140 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_260
timestamp 1682952543
transform 1 0 1148 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1682952543
transform 1 0 1140 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1682952543
transform 1 0 1204 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1682952543
transform 1 0 1172 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1682952543
transform 1 0 1244 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1682952543
transform 1 0 1276 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1682952543
transform 1 0 1340 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1682952543
transform 1 0 1276 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_145
timestamp 1682952543
transform 1 0 1284 0 1 3945
box -2 -2 2 2
use M3_M2  M3_M2_194
timestamp 1682952543
transform 1 0 1300 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1682952543
transform 1 0 1316 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_193
timestamp 1682952543
transform 1 0 1180 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1682952543
transform 1 0 1196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1682952543
transform 1 0 1204 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1682952543
transform 1 0 1212 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_197
timestamp 1682952543
transform 1 0 1244 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1682952543
transform 1 0 1172 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1682952543
transform 1 0 1188 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_261
timestamp 1682952543
transform 1 0 1196 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1682952543
transform 1 0 1252 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_198
timestamp 1682952543
transform 1 0 1260 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_234
timestamp 1682952543
transform 1 0 1268 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_199
timestamp 1682952543
transform 1 0 1276 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1682952543
transform 1 0 1292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1682952543
transform 1 0 1300 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_202
timestamp 1682952543
transform 1 0 1332 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1682952543
transform 1 0 1340 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1682952543
transform 1 0 1204 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1682952543
transform 1 0 1220 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1682952543
transform 1 0 1236 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1682952543
transform 1 0 1252 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1682952543
transform 1 0 1268 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_282
timestamp 1682952543
transform 1 0 1180 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1682952543
transform 1 0 1196 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1682952543
transform 1 0 1268 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1682952543
transform 1 0 1236 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_365
timestamp 1682952543
transform 1 0 1300 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1682952543
transform 1 0 1308 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1682952543
transform 1 0 1324 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1682952543
transform 1 0 1340 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1682952543
transform 1 0 1300 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_359
timestamp 1682952543
transform 1 0 1284 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1682952543
transform 1 0 1340 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_196
timestamp 1682952543
transform 1 0 1388 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_204
timestamp 1682952543
transform 1 0 1364 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_205
timestamp 1682952543
transform 1 0 1380 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1682952543
transform 1 0 1388 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1682952543
transform 1 0 1404 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1682952543
transform 1 0 1420 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1682952543
transform 1 0 1428 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1682952543
transform 1 0 1372 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_360
timestamp 1682952543
transform 1 0 1364 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_262
timestamp 1682952543
transform 1 0 1404 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_370
timestamp 1682952543
transform 1 0 1412 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1682952543
transform 1 0 1428 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_286
timestamp 1682952543
transform 1 0 1428 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_372
timestamp 1682952543
transform 1 0 1452 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_235
timestamp 1682952543
transform 1 0 1468 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_373
timestamp 1682952543
transform 1 0 1468 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_361
timestamp 1682952543
transform 1 0 1468 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1682952543
transform 1 0 1580 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_197
timestamp 1682952543
transform 1 0 1540 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1682952543
transform 1 0 1588 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_210
timestamp 1682952543
transform 1 0 1508 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1682952543
transform 1 0 1524 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1682952543
transform 1 0 1540 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_213
timestamp 1682952543
transform 1 0 1548 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_236
timestamp 1682952543
transform 1 0 1556 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_214
timestamp 1682952543
transform 1 0 1564 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1682952543
transform 1 0 1580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1682952543
transform 1 0 1588 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_165
timestamp 1682952543
transform 1 0 1652 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1682952543
transform 1 0 1668 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1682952543
transform 1 0 1708 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1682952543
transform 1 0 1764 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_217
timestamp 1682952543
transform 1 0 1636 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1682952543
transform 1 0 1652 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_199
timestamp 1682952543
transform 1 0 1748 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_219
timestamp 1682952543
transform 1 0 1748 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1682952543
transform 1 0 1516 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_375
timestamp 1682952543
transform 1 0 1532 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1682952543
transform 1 0 1548 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1682952543
transform 1 0 1572 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1682952543
transform 1 0 1588 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1682952543
transform 1 0 1604 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1682952543
transform 1 0 1620 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1682952543
transform 1 0 1628 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1682952543
transform 1 0 1644 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1682952543
transform 1 0 1660 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_384
timestamp 1682952543
transform 1 0 1668 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1682952543
transform 1 0 1724 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1682952543
transform 1 0 1764 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_287
timestamp 1682952543
transform 1 0 1508 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1682952543
transform 1 0 1524 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_325
timestamp 1682952543
transform 1 0 1540 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1682952543
transform 1 0 1572 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1682952543
transform 1 0 1564 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_362
timestamp 1682952543
transform 1 0 1516 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_363
timestamp 1682952543
transform 1 0 1548 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1682952543
transform 1 0 1604 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_328
timestamp 1682952543
transform 1 0 1620 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1682952543
transform 1 0 1628 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_288
timestamp 1682952543
transform 1 0 1668 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1682952543
transform 1 0 1724 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_290
timestamp 1682952543
transform 1 0 1764 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_140
timestamp 1682952543
transform 1 0 1836 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_220
timestamp 1682952543
transform 1 0 1804 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1682952543
transform 1 0 1812 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1682952543
transform 1 0 1828 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1682952543
transform 1 0 1796 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_263
timestamp 1682952543
transform 1 0 1812 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1682952543
transform 1 0 1844 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_388
timestamp 1682952543
transform 1 0 1820 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1682952543
transform 1 0 1836 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1682952543
transform 1 0 1844 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_329
timestamp 1682952543
transform 1 0 1836 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1682952543
transform 1 0 1940 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_223
timestamp 1682952543
transform 1 0 1940 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1682952543
transform 1 0 1908 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_365
timestamp 1682952543
transform 1 0 1884 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1682952543
transform 1 0 2004 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_224
timestamp 1682952543
transform 1 0 1972 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_141
timestamp 1682952543
transform 1 0 2076 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1682952543
transform 1 0 2068 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1682952543
transform 1 0 2084 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1682952543
transform 1 0 2132 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_225
timestamp 1682952543
transform 1 0 2068 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1682952543
transform 1 0 2020 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1682952543
transform 1 0 2052 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1682952543
transform 1 0 2116 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_291
timestamp 1682952543
transform 1 0 2116 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1682952543
transform 1 0 2196 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_226
timestamp 1682952543
transform 1 0 2188 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_366
timestamp 1682952543
transform 1 0 2180 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_395
timestamp 1682952543
transform 1 0 2196 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_349
timestamp 1682952543
transform 1 0 2196 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1682952543
transform 1 0 2236 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_238
timestamp 1682952543
transform 1 0 2212 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_227
timestamp 1682952543
transform 1 0 2220 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1682952543
transform 1 0 2236 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1682952543
transform 1 0 2244 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1682952543
transform 1 0 2212 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_205
timestamp 1682952543
transform 1 0 2316 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1682952543
transform 1 0 2372 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_230
timestamp 1682952543
transform 1 0 2340 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1682952543
transform 1 0 2356 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_232
timestamp 1682952543
transform 1 0 2372 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1682952543
transform 1 0 2252 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1682952543
transform 1 0 2260 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1682952543
transform 1 0 2316 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_264
timestamp 1682952543
transform 1 0 2356 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_400
timestamp 1682952543
transform 1 0 2364 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_401
timestamp 1682952543
transform 1 0 2380 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_292
timestamp 1682952543
transform 1 0 2292 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_330
timestamp 1682952543
transform 1 0 2252 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_350
timestamp 1682952543
transform 1 0 2268 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_207
timestamp 1682952543
transform 1 0 2396 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_233
timestamp 1682952543
transform 1 0 2396 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1682952543
transform 1 0 2404 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_265
timestamp 1682952543
transform 1 0 2404 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1682952543
transform 1 0 2444 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_235
timestamp 1682952543
transform 1 0 2428 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1682952543
transform 1 0 2444 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1682952543
transform 1 0 2452 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1682952543
transform 1 0 2420 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1682952543
transform 1 0 2436 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_266
timestamp 1682952543
transform 1 0 2452 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_331
timestamp 1682952543
transform 1 0 2444 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1682952543
transform 1 0 2420 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_209
timestamp 1682952543
transform 1 0 2500 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1682952543
transform 1 0 2476 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_238
timestamp 1682952543
transform 1 0 2484 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1682952543
transform 1 0 2500 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1682952543
transform 1 0 2476 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1682952543
transform 1 0 2532 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_210
timestamp 1682952543
transform 1 0 2556 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_241
timestamp 1682952543
transform 1 0 2556 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1682952543
transform 1 0 2548 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_211
timestamp 1682952543
transform 1 0 2676 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_242
timestamp 1682952543
transform 1 0 2572 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1682952543
transform 1 0 2588 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1682952543
transform 1 0 2604 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1682952543
transform 1 0 2620 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1682952543
transform 1 0 2636 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_406
timestamp 1682952543
transform 1 0 2564 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_293
timestamp 1682952543
transform 1 0 2564 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_407
timestamp 1682952543
transform 1 0 2588 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1682952543
transform 1 0 2612 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_294
timestamp 1682952543
transform 1 0 2588 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_267
timestamp 1682952543
transform 1 0 2620 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_409
timestamp 1682952543
transform 1 0 2676 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_295
timestamp 1682952543
transform 1 0 2700 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1682952543
transform 1 0 2596 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1682952543
transform 1 0 2628 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_334
timestamp 1682952543
transform 1 0 2708 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1682952543
transform 1 0 2740 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_247
timestamp 1682952543
transform 1 0 2740 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1682952543
transform 1 0 2732 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_144
timestamp 1682952543
transform 1 0 2788 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_212
timestamp 1682952543
transform 1 0 2764 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1682952543
transform 1 0 2780 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1682952543
transform 1 0 2860 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_248
timestamp 1682952543
transform 1 0 2764 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1682952543
transform 1 0 2780 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1682952543
transform 1 0 2788 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_251
timestamp 1682952543
transform 1 0 2804 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1682952543
transform 1 0 2828 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_411
timestamp 1682952543
transform 1 0 2772 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1682952543
transform 1 0 2788 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1682952543
transform 1 0 2812 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_296
timestamp 1682952543
transform 1 0 2772 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1682952543
transform 1 0 2812 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1682952543
transform 1 0 2788 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1682952543
transform 1 0 2836 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1682952543
transform 1 0 2868 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1682952543
transform 1 0 2844 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1682952543
transform 1 0 2860 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_255
timestamp 1682952543
transform 1 0 2868 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1682952543
transform 1 0 2836 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1682952543
transform 1 0 2852 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_146
timestamp 1682952543
transform 1 0 2932 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1682952543
transform 1 0 2924 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_256
timestamp 1682952543
transform 1 0 2892 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1682952543
transform 1 0 2908 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1682952543
transform 1 0 2884 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_241
timestamp 1682952543
transform 1 0 2916 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_258
timestamp 1682952543
transform 1 0 2924 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1682952543
transform 1 0 2932 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1682952543
transform 1 0 2916 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_367
timestamp 1682952543
transform 1 0 2892 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_418
timestamp 1682952543
transform 1 0 2940 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_147
timestamp 1682952543
transform 1 0 3076 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_171
timestamp 1682952543
transform 1 0 2988 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1682952543
transform 1 0 3004 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1682952543
transform 1 0 3124 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1682952543
transform 1 0 3172 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_260
timestamp 1682952543
transform 1 0 2972 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1682952543
transform 1 0 2988 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1682952543
transform 1 0 3076 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_263
timestamp 1682952543
transform 1 0 3092 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1682952543
transform 1 0 3108 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_265
timestamp 1682952543
transform 1 0 3124 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1682952543
transform 1 0 3140 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1682952543
transform 1 0 2964 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1682952543
transform 1 0 2980 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1682952543
transform 1 0 2996 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_422
timestamp 1682952543
transform 1 0 3028 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_298
timestamp 1682952543
transform 1 0 2980 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_299
timestamp 1682952543
transform 1 0 3012 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_368
timestamp 1682952543
transform 1 0 3036 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_423
timestamp 1682952543
transform 1 0 3100 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1682952543
transform 1 0 3116 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_352
timestamp 1682952543
transform 1 0 3116 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_425
timestamp 1682952543
transform 1 0 3164 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1682952543
transform 1 0 3220 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1682952543
transform 1 0 3228 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1682952543
transform 1 0 3236 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1682952543
transform 1 0 3244 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_173
timestamp 1682952543
transform 1 0 3252 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1682952543
transform 1 0 3300 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_174
timestamp 1682952543
transform 1 0 3292 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1682952543
transform 1 0 3340 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1682952543
transform 1 0 3300 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1682952543
transform 1 0 3340 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_269
timestamp 1682952543
transform 1 0 3260 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1682952543
transform 1 0 3276 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1682952543
transform 1 0 3292 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1682952543
transform 1 0 3300 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1682952543
transform 1 0 3316 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_274
timestamp 1682952543
transform 1 0 3332 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1682952543
transform 1 0 3340 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1682952543
transform 1 0 3252 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1682952543
transform 1 0 3260 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1682952543
transform 1 0 3268 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1682952543
transform 1 0 3284 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1682952543
transform 1 0 3300 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1682952543
transform 1 0 3324 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_434
timestamp 1682952543
transform 1 0 3340 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_300
timestamp 1682952543
transform 1 0 3284 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_301
timestamp 1682952543
transform 1 0 3324 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_353
timestamp 1682952543
transform 1 0 3340 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_435
timestamp 1682952543
transform 1 0 3356 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_219
timestamp 1682952543
transform 1 0 3372 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_276
timestamp 1682952543
transform 1 0 3372 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1682952543
transform 1 0 3388 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_278
timestamp 1682952543
transform 1 0 3404 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1682952543
transform 1 0 3492 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1682952543
transform 1 0 3396 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_268
timestamp 1682952543
transform 1 0 3404 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1682952543
transform 1 0 3516 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_280
timestamp 1682952543
transform 1 0 3508 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1682952543
transform 1 0 3412 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1682952543
transform 1 0 3444 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_269
timestamp 1682952543
transform 1 0 3508 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1682952543
transform 1 0 3388 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_303
timestamp 1682952543
transform 1 0 3404 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1682952543
transform 1 0 3444 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1682952543
transform 1 0 3396 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1682952543
transform 1 0 3372 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1682952543
transform 1 0 3388 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1682952543
transform 1 0 3420 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1682952543
transform 1 0 3556 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1682952543
transform 1 0 3588 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1682952543
transform 1 0 3548 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1682952543
transform 1 0 3572 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_242
timestamp 1682952543
transform 1 0 3524 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_281
timestamp 1682952543
transform 1 0 3532 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1682952543
transform 1 0 3548 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_283
timestamp 1682952543
transform 1 0 3556 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1682952543
transform 1 0 3572 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1682952543
transform 1 0 3580 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1682952543
transform 1 0 3596 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_285
timestamp 1682952543
transform 1 0 3588 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1682952543
transform 1 0 3596 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1682952543
transform 1 0 3524 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_440
timestamp 1682952543
transform 1 0 3556 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1682952543
transform 1 0 3564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1682952543
transform 1 0 3580 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_371
timestamp 1682952543
transform 1 0 3516 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_305
timestamp 1682952543
transform 1 0 3556 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_443
timestamp 1682952543
transform 1 0 3596 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_306
timestamp 1682952543
transform 1 0 3596 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1682952543
transform 1 0 3660 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_287
timestamp 1682952543
transform 1 0 3628 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_244
timestamp 1682952543
transform 1 0 3636 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1682952543
transform 1 0 3716 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_288
timestamp 1682952543
transform 1 0 3644 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1682952543
transform 1 0 3660 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1682952543
transform 1 0 3668 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1682952543
transform 1 0 3684 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1682952543
transform 1 0 3700 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1682952543
transform 1 0 3636 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1682952543
transform 1 0 3652 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_354
timestamp 1682952543
transform 1 0 3628 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_245
timestamp 1682952543
transform 1 0 3708 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_293
timestamp 1682952543
transform 1 0 3716 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_446
timestamp 1682952543
transform 1 0 3692 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1682952543
transform 1 0 3708 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1682952543
transform 1 0 3724 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_223
timestamp 1682952543
transform 1 0 3732 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1682952543
transform 1 0 3764 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_294
timestamp 1682952543
transform 1 0 3732 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1682952543
transform 1 0 3748 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_307
timestamp 1682952543
transform 1 0 3692 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_308
timestamp 1682952543
transform 1 0 3724 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1682952543
transform 1 0 3684 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_449
timestamp 1682952543
transform 1 0 3796 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_355
timestamp 1682952543
transform 1 0 3748 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_356
timestamp 1682952543
transform 1 0 3764 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_373
timestamp 1682952543
transform 1 0 3820 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_180
timestamp 1682952543
transform 1 0 3900 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1682952543
transform 1 0 3860 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1682952543
transform 1 0 3884 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_296
timestamp 1682952543
transform 1 0 3852 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1682952543
transform 1 0 3868 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1682952543
transform 1 0 3876 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1682952543
transform 1 0 3932 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_298
timestamp 1682952543
transform 1 0 3884 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1682952543
transform 1 0 3892 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1682952543
transform 1 0 3908 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1682952543
transform 1 0 3924 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1682952543
transform 1 0 3932 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1682952543
transform 1 0 3844 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1682952543
transform 1 0 3852 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1682952543
transform 1 0 3860 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1682952543
transform 1 0 3876 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_357
timestamp 1682952543
transform 1 0 3852 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_270
timestamp 1682952543
transform 1 0 3884 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_454
timestamp 1682952543
transform 1 0 3892 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1682952543
transform 1 0 3916 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_271
timestamp 1682952543
transform 1 0 3924 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1682952543
transform 1 0 3892 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_303
timestamp 1682952543
transform 1 0 3948 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1682952543
transform 1 0 3956 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_310
timestamp 1682952543
transform 1 0 3972 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1682952543
transform 1 0 4004 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1682952543
transform 1 0 3988 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_304
timestamp 1682952543
transform 1 0 3996 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1682952543
transform 1 0 4012 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1682952543
transform 1 0 3988 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1682952543
transform 1 0 4004 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_181
timestamp 1682952543
transform 1 0 4044 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1682952543
transform 1 0 4068 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_306
timestamp 1682952543
transform 1 0 4068 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_248
timestamp 1682952543
transform 1 0 4116 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_459
timestamp 1682952543
transform 1 0 4092 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1682952543
transform 1 0 4148 0 1 3925
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_4
timestamp 1682952543
transform 1 0 24 0 1 3870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_21
timestamp 1682952543
transform 1 0 72 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_10
timestamp 1682952543
transform -1 0 184 0 -1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1682952543
transform 1 0 184 0 -1 3970
box -8 -3 104 105
use AOI22X1  AOI22X1_1
timestamp 1682952543
transform 1 0 280 0 -1 3970
box -8 -3 46 105
use FILL  FILL_31
timestamp 1682952543
transform 1 0 320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_32
timestamp 1682952543
transform 1 0 328 0 -1 3970
box -8 -3 16 105
use FILL  FILL_33
timestamp 1682952543
transform 1 0 336 0 -1 3970
box -8 -3 16 105
use FILL  FILL_34
timestamp 1682952543
transform 1 0 344 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1682952543
transform 1 0 352 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_0
timestamp 1682952543
transform 1 0 392 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_1
timestamp 1682952543
transform 1 0 432 0 -1 3970
box -8 -3 46 105
use FILL  FILL_35
timestamp 1682952543
transform 1 0 472 0 -1 3970
box -8 -3 16 105
use FILL  FILL_36
timestamp 1682952543
transform 1 0 480 0 -1 3970
box -8 -3 16 105
use FILL  FILL_37
timestamp 1682952543
transform 1 0 488 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_3
timestamp 1682952543
transform 1 0 496 0 -1 3970
box -8 -3 46 105
use FILL  FILL_38
timestamp 1682952543
transform 1 0 536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_39
timestamp 1682952543
transform 1 0 544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_40
timestamp 1682952543
transform 1 0 552 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_11
timestamp 1682952543
transform -1 0 576 0 -1 3970
box -9 -3 26 105
use FILL  FILL_41
timestamp 1682952543
transform 1 0 576 0 -1 3970
box -8 -3 16 105
use FILL  FILL_42
timestamp 1682952543
transform 1 0 584 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_374
timestamp 1682952543
transform 1 0 604 0 1 3875
box -3 -3 3 3
use AOI22X1  AOI22X1_4
timestamp 1682952543
transform 1 0 592 0 -1 3970
box -8 -3 46 105
use M3_M2  M3_M2_375
timestamp 1682952543
transform 1 0 660 0 1 3875
box -3 -3 3 3
use AOI22X1  AOI22X1_5
timestamp 1682952543
transform -1 0 672 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_12
timestamp 1682952543
transform 1 0 672 0 -1 3970
box -9 -3 26 105
use M3_M2  M3_M2_376
timestamp 1682952543
transform 1 0 708 0 1 3875
box -3 -3 3 3
use OAI22X1  OAI22X1_2
timestamp 1682952543
transform 1 0 688 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_6
timestamp 1682952543
transform -1 0 768 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_13
timestamp 1682952543
transform 1 0 768 0 -1 3970
box -9 -3 26 105
use OAI22X1  OAI22X1_3
timestamp 1682952543
transform 1 0 784 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_7
timestamp 1682952543
transform 1 0 824 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_4
timestamp 1682952543
transform 1 0 864 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_8
timestamp 1682952543
transform -1 0 944 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_14
timestamp 1682952543
transform 1 0 944 0 -1 3970
box -9 -3 26 105
use M3_M2  M3_M2_377
timestamp 1682952543
transform 1 0 980 0 1 3875
box -3 -3 3 3
use NOR2X1  NOR2X1_0
timestamp 1682952543
transform 1 0 960 0 -1 3970
box -8 -3 32 105
use FILL  FILL_43
timestamp 1682952543
transform 1 0 984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_44
timestamp 1682952543
transform 1 0 992 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_378
timestamp 1682952543
transform 1 0 1028 0 1 3875
box -3 -3 3 3
use NOR2X1  NOR2X1_1
timestamp 1682952543
transform 1 0 1000 0 -1 3970
box -8 -3 32 105
use AOI22X1  AOI22X1_9
timestamp 1682952543
transform 1 0 1024 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_15
timestamp 1682952543
transform 1 0 1064 0 -1 3970
box -9 -3 26 105
use FILL  FILL_45
timestamp 1682952543
transform 1 0 1080 0 -1 3970
box -8 -3 16 105
use FILL  FILL_46
timestamp 1682952543
transform 1 0 1088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_47
timestamp 1682952543
transform 1 0 1096 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_10
timestamp 1682952543
transform 1 0 1104 0 -1 3970
box -8 -3 46 105
use FILL  FILL_48
timestamp 1682952543
transform 1 0 1144 0 -1 3970
box -8 -3 16 105
use FILL  FILL_49
timestamp 1682952543
transform 1 0 1152 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_5
timestamp 1682952543
transform -1 0 1200 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1682952543
transform 1 0 1200 0 -1 3970
box -8 -3 46 105
use M3_M2  M3_M2_379
timestamp 1682952543
transform 1 0 1252 0 1 3875
box -3 -3 3 3
use OAI22X1  OAI22X1_6
timestamp 1682952543
transform -1 0 1280 0 -1 3970
box -8 -3 46 105
use NOR2X1  NOR2X1_2
timestamp 1682952543
transform 1 0 1280 0 -1 3970
box -8 -3 32 105
use AOI22X1  AOI22X1_12
timestamp 1682952543
transform -1 0 1344 0 -1 3970
box -8 -3 46 105
use FILL  FILL_50
timestamp 1682952543
transform 1 0 1344 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_13
timestamp 1682952543
transform 1 0 1352 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_14
timestamp 1682952543
transform -1 0 1432 0 -1 3970
box -8 -3 46 105
use FILL  FILL_51
timestamp 1682952543
transform 1 0 1432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_52
timestamp 1682952543
transform 1 0 1440 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_16
timestamp 1682952543
transform 1 0 1448 0 -1 3970
box -9 -3 26 105
use FILL  FILL_53
timestamp 1682952543
transform 1 0 1464 0 -1 3970
box -8 -3 16 105
use FILL  FILL_54
timestamp 1682952543
transform 1 0 1472 0 -1 3970
box -8 -3 16 105
use FILL  FILL_55
timestamp 1682952543
transform 1 0 1480 0 -1 3970
box -8 -3 16 105
use FILL  FILL_56
timestamp 1682952543
transform 1 0 1488 0 -1 3970
box -8 -3 16 105
use FILL  FILL_57
timestamp 1682952543
transform 1 0 1496 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_380
timestamp 1682952543
transform 1 0 1532 0 1 3875
box -3 -3 3 3
use OAI22X1  OAI22X1_7
timestamp 1682952543
transform 1 0 1504 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_8
timestamp 1682952543
transform 1 0 1544 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_15
timestamp 1682952543
transform -1 0 1624 0 -1 3970
box -8 -3 46 105
use AOI22X1  AOI22X1_16
timestamp 1682952543
transform 1 0 1624 0 -1 3970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1682952543
transform -1 0 1760 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_17
timestamp 1682952543
transform -1 0 1776 0 -1 3970
box -9 -3 26 105
use FILL  FILL_58
timestamp 1682952543
transform 1 0 1776 0 -1 3970
box -8 -3 16 105
use FILL  FILL_59
timestamp 1682952543
transform 1 0 1784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_60
timestamp 1682952543
transform 1 0 1792 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_17
timestamp 1682952543
transform -1 0 1840 0 -1 3970
box -8 -3 46 105
use FILL  FILL_61
timestamp 1682952543
transform 1 0 1840 0 -1 3970
box -8 -3 16 105
use FILL  FILL_62
timestamp 1682952543
transform 1 0 1848 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1682952543
transform -1 0 1952 0 -1 3970
box -8 -3 104 105
use FILL  FILL_63
timestamp 1682952543
transform 1 0 1952 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1682952543
transform 1 0 1960 0 -1 3970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1682952543
transform 1 0 2056 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_18
timestamp 1682952543
transform 1 0 2152 0 -1 3970
box -9 -3 26 105
use FILL  FILL_64
timestamp 1682952543
transform 1 0 2168 0 -1 3970
box -8 -3 16 105
use FILL  FILL_65
timestamp 1682952543
transform 1 0 2176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_66
timestamp 1682952543
transform 1 0 2184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_67
timestamp 1682952543
transform 1 0 2192 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_9
timestamp 1682952543
transform -1 0 2240 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_19
timestamp 1682952543
transform 1 0 2240 0 -1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1682952543
transform -1 0 2352 0 -1 3970
box -8 -3 104 105
use OAI22X1  OAI22X1_10
timestamp 1682952543
transform -1 0 2392 0 -1 3970
box -8 -3 46 105
use FILL  FILL_68
timestamp 1682952543
transform 1 0 2392 0 -1 3970
box -8 -3 16 105
use FILL  FILL_69
timestamp 1682952543
transform 1 0 2400 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_11
timestamp 1682952543
transform -1 0 2448 0 -1 3970
box -8 -3 46 105
use FILL  FILL_70
timestamp 1682952543
transform 1 0 2448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_71
timestamp 1682952543
transform 1 0 2456 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_12
timestamp 1682952543
transform -1 0 2504 0 -1 3970
box -8 -3 46 105
use FILL  FILL_72
timestamp 1682952543
transform 1 0 2504 0 -1 3970
box -8 -3 16 105
use FILL  FILL_73
timestamp 1682952543
transform 1 0 2512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_74
timestamp 1682952543
transform 1 0 2520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_75
timestamp 1682952543
transform 1 0 2528 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_381
timestamp 1682952543
transform 1 0 2556 0 1 3875
box -3 -3 3 3
use INVX2  INVX2_20
timestamp 1682952543
transform 1 0 2536 0 -1 3970
box -9 -3 26 105
use FILL  FILL_79
timestamp 1682952543
transform 1 0 2552 0 -1 3970
box -8 -3 16 105
use FILL  FILL_81
timestamp 1682952543
transform 1 0 2560 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_24
timestamp 1682952543
transform 1 0 2568 0 -1 3970
box -9 -3 26 105
use OAI22X1  OAI22X1_13
timestamp 1682952543
transform 1 0 2584 0 -1 3970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1682952543
transform 1 0 2624 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_25
timestamp 1682952543
transform 1 0 2720 0 -1 3970
box -9 -3 26 105
use FILL  FILL_88
timestamp 1682952543
transform 1 0 2736 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_14
timestamp 1682952543
transform 1 0 2744 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_15
timestamp 1682952543
transform 1 0 2784 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_16
timestamp 1682952543
transform -1 0 2864 0 -1 3970
box -8 -3 46 105
use FILL  FILL_89
timestamp 1682952543
transform 1 0 2864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_90
timestamp 1682952543
transform 1 0 2872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_91
timestamp 1682952543
transform 1 0 2880 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_17
timestamp 1682952543
transform 1 0 2888 0 -1 3970
box -8 -3 46 105
use FILL  FILL_92
timestamp 1682952543
transform 1 0 2928 0 -1 3970
box -8 -3 16 105
use FILL  FILL_93
timestamp 1682952543
transform 1 0 2936 0 -1 3970
box -8 -3 16 105
use FILL  FILL_94
timestamp 1682952543
transform 1 0 2944 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_18
timestamp 1682952543
transform 1 0 2952 0 -1 3970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_35
timestamp 1682952543
transform -1 0 3088 0 -1 3970
box -8 -3 104 105
use OAI22X1  OAI22X1_19
timestamp 1682952543
transform 1 0 3088 0 -1 3970
box -8 -3 46 105
use M3_M2  M3_M2_382
timestamp 1682952543
transform 1 0 3164 0 1 3875
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1682952543
transform 1 0 3228 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_36
timestamp 1682952543
transform 1 0 3128 0 -1 3970
box -8 -3 104 105
use M3_M2  M3_M2_384
timestamp 1682952543
transform 1 0 3244 0 1 3875
box -3 -3 3 3
use INVX2  INVX2_29
timestamp 1682952543
transform -1 0 3240 0 -1 3970
box -9 -3 26 105
use INVX2  INVX2_30
timestamp 1682952543
transform 1 0 3240 0 -1 3970
box -9 -3 26 105
use OAI22X1  OAI22X1_20
timestamp 1682952543
transform 1 0 3256 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_21
timestamp 1682952543
transform 1 0 3296 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_31
timestamp 1682952543
transform 1 0 3336 0 -1 3970
box -9 -3 26 105
use FILL  FILL_104
timestamp 1682952543
transform 1 0 3352 0 -1 3970
box -8 -3 16 105
use FILL  FILL_112
timestamp 1682952543
transform 1 0 3360 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_22
timestamp 1682952543
transform 1 0 3368 0 -1 3970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1682952543
transform -1 0 3504 0 -1 3970
box -8 -3 104 105
use FILL  FILL_113
timestamp 1682952543
transform 1 0 3504 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_23
timestamp 1682952543
transform -1 0 3552 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_24
timestamp 1682952543
transform 1 0 3552 0 -1 3970
box -8 -3 46 105
use FILL  FILL_114
timestamp 1682952543
transform 1 0 3592 0 -1 3970
box -8 -3 16 105
use FILL  FILL_115
timestamp 1682952543
transform 1 0 3600 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_36
timestamp 1682952543
transform 1 0 3608 0 -1 3970
box -9 -3 26 105
use OAI22X1  OAI22X1_25
timestamp 1682952543
transform -1 0 3664 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_37
timestamp 1682952543
transform 1 0 3664 0 -1 3970
box -9 -3 26 105
use OAI22X1  OAI22X1_26
timestamp 1682952543
transform 1 0 3680 0 -1 3970
box -8 -3 46 105
use INVX2  INVX2_38
timestamp 1682952543
transform -1 0 3736 0 -1 3970
box -9 -3 26 105
use M3_M2  M3_M2_385
timestamp 1682952543
transform 1 0 3788 0 1 3875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_45
timestamp 1682952543
transform 1 0 3736 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_39
timestamp 1682952543
transform 1 0 3832 0 -1 3970
box -9 -3 26 105
use OAI22X1  OAI22X1_27
timestamp 1682952543
transform 1 0 3848 0 -1 3970
box -8 -3 46 105
use OAI22X1  OAI22X1_28
timestamp 1682952543
transform 1 0 3888 0 -1 3970
box -8 -3 46 105
use FILL  FILL_116
timestamp 1682952543
transform 1 0 3928 0 -1 3970
box -8 -3 16 105
use FILL  FILL_117
timestamp 1682952543
transform 1 0 3936 0 -1 3970
box -8 -3 16 105
use FILL  FILL_118
timestamp 1682952543
transform 1 0 3944 0 -1 3970
box -8 -3 16 105
use FILL  FILL_119
timestamp 1682952543
transform 1 0 3952 0 -1 3970
box -8 -3 16 105
use FILL  FILL_120
timestamp 1682952543
transform 1 0 3960 0 -1 3970
box -8 -3 16 105
use FILL  FILL_121
timestamp 1682952543
transform 1 0 3968 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_29
timestamp 1682952543
transform 1 0 3976 0 -1 3970
box -8 -3 46 105
use FILL  FILL_122
timestamp 1682952543
transform 1 0 4016 0 -1 3970
box -8 -3 16 105
use FILL  FILL_123
timestamp 1682952543
transform 1 0 4024 0 -1 3970
box -8 -3 16 105
use FILL  FILL_124
timestamp 1682952543
transform 1 0 4032 0 -1 3970
box -8 -3 16 105
use FILL  FILL_125
timestamp 1682952543
transform 1 0 4040 0 -1 3970
box -8 -3 16 105
use FILL  FILL_126
timestamp 1682952543
transform 1 0 4048 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1682952543
transform 1 0 4056 0 -1 3970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_5
timestamp 1682952543
transform 1 0 4201 0 1 3870
box -10 -3 10 3
use M3_M2  M3_M2_423
timestamp 1682952543
transform 1 0 132 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_461
timestamp 1682952543
transform 1 0 116 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1682952543
transform 1 0 124 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_544
timestamp 1682952543
transform 1 0 124 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1682952543
transform 1 0 140 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1682952543
transform 1 0 164 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1682952543
transform 1 0 164 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_463
timestamp 1682952543
transform 1 0 148 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1682952543
transform 1 0 164 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1682952543
transform 1 0 180 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1682952543
transform 1 0 140 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1682952543
transform 1 0 148 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_545
timestamp 1682952543
transform 1 0 172 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1682952543
transform 1 0 204 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1682952543
transform 1 0 196 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_466
timestamp 1682952543
transform 1 0 204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1682952543
transform 1 0 196 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_502
timestamp 1682952543
transform 1 0 220 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_467
timestamp 1682952543
transform 1 0 228 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_503
timestamp 1682952543
transform 1 0 252 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_386
timestamp 1682952543
transform 1 0 284 0 1 3865
box -3 -3 3 3
use M2_M1  M2_M1_468
timestamp 1682952543
transform 1 0 284 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_504
timestamp 1682952543
transform 1 0 292 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_469
timestamp 1682952543
transform 1 0 300 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_409
timestamp 1682952543
transform 1 0 324 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_450
timestamp 1682952543
transform 1 0 324 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_470
timestamp 1682952543
transform 1 0 324 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_588
timestamp 1682952543
transform 1 0 284 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1682952543
transform 1 0 292 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1682952543
transform 1 0 308 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1682952543
transform 1 0 316 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_546
timestamp 1682952543
transform 1 0 316 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_471
timestamp 1682952543
transform 1 0 348 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_505
timestamp 1682952543
transform 1 0 356 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_472
timestamp 1682952543
transform 1 0 364 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1682952543
transform 1 0 332 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1682952543
transform 1 0 356 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1682952543
transform 1 0 364 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_425
timestamp 1682952543
transform 1 0 484 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1682952543
transform 1 0 380 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_452
timestamp 1682952543
transform 1 0 420 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_453
timestamp 1682952543
transform 1 0 436 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_473
timestamp 1682952543
transform 1 0 380 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1682952543
transform 1 0 420 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_506
timestamp 1682952543
transform 1 0 460 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1682952543
transform 1 0 492 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_475
timestamp 1682952543
transform 1 0 476 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1682952543
transform 1 0 492 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1682952543
transform 1 0 508 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1682952543
transform 1 0 396 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1682952543
transform 1 0 476 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_596
timestamp 1682952543
transform 1 0 484 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1682952543
transform 1 0 500 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1682952543
transform 1 0 508 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1682952543
transform 1 0 580 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1682952543
transform 1 0 668 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1682952543
transform 1 0 628 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_456
timestamp 1682952543
transform 1 0 668 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_478
timestamp 1682952543
transform 1 0 564 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_479
timestamp 1682952543
transform 1 0 620 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1682952543
transform 1 0 628 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_481
timestamp 1682952543
transform 1 0 668 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1682952543
transform 1 0 724 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1682952543
transform 1 0 516 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1682952543
transform 1 0 532 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1682952543
transform 1 0 620 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_586
timestamp 1682952543
transform 1 0 500 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1682952543
transform 1 0 532 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_601
timestamp 1682952543
transform 1 0 644 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_548
timestamp 1682952543
transform 1 0 644 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_602
timestamp 1682952543
transform 1 0 740 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_398
timestamp 1682952543
transform 1 0 828 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_411
timestamp 1682952543
transform 1 0 764 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_457
timestamp 1682952543
transform 1 0 756 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1682952543
transform 1 0 796 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_483
timestamp 1682952543
transform 1 0 756 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1682952543
transform 1 0 764 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1682952543
transform 1 0 796 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_507
timestamp 1682952543
transform 1 0 804 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1682952543
transform 1 0 940 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1682952543
transform 1 0 868 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_486
timestamp 1682952543
transform 1 0 860 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_487
timestamp 1682952543
transform 1 0 916 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_534
timestamp 1682952543
transform 1 0 764 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1682952543
transform 1 0 796 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_603
timestamp 1682952543
transform 1 0 844 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_549
timestamp 1682952543
transform 1 0 844 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_604
timestamp 1682952543
transform 1 0 940 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_536
timestamp 1682952543
transform 1 0 956 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1682952543
transform 1 0 876 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_551
timestamp 1682952543
transform 1 0 900 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_552
timestamp 1682952543
transform 1 0 940 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_703
timestamp 1682952543
transform 1 0 956 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_587
timestamp 1682952543
transform 1 0 956 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1682952543
transform 1 0 972 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_488
timestamp 1682952543
transform 1 0 972 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_412
timestamp 1682952543
transform 1 0 1108 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_426
timestamp 1682952543
transform 1 0 1012 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_427
timestamp 1682952543
transform 1 0 1052 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1682952543
transform 1 0 1092 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1682952543
transform 1 0 1060 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1682952543
transform 1 0 1108 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_489
timestamp 1682952543
transform 1 0 996 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_490
timestamp 1682952543
transform 1 0 1060 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1682952543
transform 1 0 1092 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_492
timestamp 1682952543
transform 1 0 1108 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1682952543
transform 1 0 972 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1682952543
transform 1 0 988 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_704
timestamp 1682952543
transform 1 0 980 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1682952543
transform 1 0 1012 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_553
timestamp 1682952543
transform 1 0 996 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1682952543
transform 1 0 1012 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1682952543
transform 1 0 1076 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1682952543
transform 1 0 1132 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_608
timestamp 1682952543
transform 1 0 1124 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1682952543
transform 1 0 1132 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1682952543
transform 1 0 1148 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1682952543
transform 1 0 1156 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_554
timestamp 1682952543
transform 1 0 1156 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_555
timestamp 1682952543
transform 1 0 1172 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1682952543
transform 1 0 1204 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_463
timestamp 1682952543
transform 1 0 1204 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_494
timestamp 1682952543
transform 1 0 1196 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1682952543
transform 1 0 1204 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1682952543
transform 1 0 1220 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_497
timestamp 1682952543
transform 1 0 1236 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_508
timestamp 1682952543
transform 1 0 1244 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1682952543
transform 1 0 1332 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1682952543
transform 1 0 1292 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1682952543
transform 1 0 1308 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_498
timestamp 1682952543
transform 1 0 1260 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_499
timestamp 1682952543
transform 1 0 1300 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_500
timestamp 1682952543
transform 1 0 1356 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1682952543
transform 1 0 1204 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1682952543
transform 1 0 1212 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1682952543
transform 1 0 1228 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1682952543
transform 1 0 1236 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_556
timestamp 1682952543
transform 1 0 1228 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_705
timestamp 1682952543
transform 1 0 1244 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_590
timestamp 1682952543
transform 1 0 1204 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_615
timestamp 1682952543
transform 1 0 1276 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_557
timestamp 1682952543
transform 1 0 1356 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_616
timestamp 1682952543
transform 1 0 1372 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_591
timestamp 1682952543
transform 1 0 1380 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1682952543
transform 1 0 1420 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_414
timestamp 1682952543
transform 1 0 1460 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_430
timestamp 1682952543
transform 1 0 1508 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1682952543
transform 1 0 1404 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1682952543
transform 1 0 1444 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1682952543
transform 1 0 1468 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_431
timestamp 1682952543
transform 1 0 1540 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_501
timestamp 1682952543
transform 1 0 1404 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_502
timestamp 1682952543
transform 1 0 1412 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_503
timestamp 1682952543
transform 1 0 1444 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_504
timestamp 1682952543
transform 1 0 1508 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1682952543
transform 1 0 1524 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1682952543
transform 1 0 1540 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1682952543
transform 1 0 1492 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_592
timestamp 1682952543
transform 1 0 1412 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_618
timestamp 1682952543
transform 1 0 1516 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1682952543
transform 1 0 1532 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1682952543
transform 1 0 1540 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_558
timestamp 1682952543
transform 1 0 1524 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_559
timestamp 1682952543
transform 1 0 1540 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1682952543
transform 1 0 1516 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1682952543
transform 1 0 1620 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1682952543
transform 1 0 1588 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1682952543
transform 1 0 1652 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1682952543
transform 1 0 1620 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_507
timestamp 1682952543
transform 1 0 1572 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1682952543
transform 1 0 1580 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1682952543
transform 1 0 1604 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_509
timestamp 1682952543
transform 1 0 1612 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_510
timestamp 1682952543
transform 1 0 1620 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1682952543
transform 1 0 1636 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_510
timestamp 1682952543
transform 1 0 1644 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_512
timestamp 1682952543
transform 1 0 1652 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1682952543
transform 1 0 1580 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_537
timestamp 1682952543
transform 1 0 1588 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_622
timestamp 1682952543
transform 1 0 1596 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1682952543
transform 1 0 1612 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1682952543
transform 1 0 1620 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_625
timestamp 1682952543
transform 1 0 1628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1682952543
transform 1 0 1644 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1682952543
transform 1 0 1652 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_560
timestamp 1682952543
transform 1 0 1580 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_594
timestamp 1682952543
transform 1 0 1596 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1682952543
transform 1 0 1620 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1682952543
transform 1 0 1684 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1682952543
transform 1 0 1724 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_513
timestamp 1682952543
transform 1 0 1684 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1682952543
transform 1 0 1692 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_511
timestamp 1682952543
transform 1 0 1700 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_515
timestamp 1682952543
transform 1 0 1724 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1682952543
transform 1 0 1772 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_471
timestamp 1682952543
transform 1 0 1796 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1682952543
transform 1 0 1828 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_516
timestamp 1682952543
transform 1 0 1796 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1682952543
transform 1 0 1812 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1682952543
transform 1 0 1788 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_561
timestamp 1682952543
transform 1 0 1740 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_562
timestamp 1682952543
transform 1 0 1788 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1682952543
transform 1 0 1820 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1682952543
transform 1 0 1836 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_518
timestamp 1682952543
transform 1 0 1828 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1682952543
transform 1 0 1836 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1682952543
transform 1 0 1820 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_596
timestamp 1682952543
transform 1 0 1820 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_631
timestamp 1682952543
transform 1 0 1844 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1682952543
transform 1 0 1868 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1682952543
transform 1 0 1876 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_521
timestamp 1682952543
transform 1 0 1884 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1682952543
transform 1 0 1876 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_633
timestamp 1682952543
transform 1 0 1884 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_597
timestamp 1682952543
transform 1 0 1868 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_522
timestamp 1682952543
transform 1 0 1908 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_415
timestamp 1682952543
transform 1 0 1924 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_523
timestamp 1682952543
transform 1 0 1924 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_416
timestamp 1682952543
transform 1 0 2052 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_435
timestamp 1682952543
transform 1 0 1996 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1682952543
transform 1 0 2044 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1682952543
transform 1 0 2012 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1682952543
transform 1 0 2036 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_524
timestamp 1682952543
transform 1 0 2012 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1682952543
transform 1 0 2036 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1682952543
transform 1 0 2124 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_476
timestamp 1682952543
transform 1 0 2140 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_525
timestamp 1682952543
transform 1 0 2140 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1682952543
transform 1 0 2092 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_563
timestamp 1682952543
transform 1 0 2140 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_390
timestamp 1682952543
transform 1 0 2188 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_391
timestamp 1682952543
transform 1 0 2252 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1682952543
transform 1 0 2244 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_526
timestamp 1682952543
transform 1 0 2228 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1682952543
transform 1 0 2244 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_402
timestamp 1682952543
transform 1 0 2276 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1682952543
transform 1 0 2268 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1682952543
transform 1 0 2260 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_528
timestamp 1682952543
transform 1 0 2268 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1682952543
transform 1 0 2220 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_637
timestamp 1682952543
transform 1 0 2236 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1682952543
transform 1 0 2252 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1682952543
transform 1 0 2260 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_564
timestamp 1682952543
transform 1 0 2236 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1682952543
transform 1 0 2252 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1682952543
transform 1 0 2220 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1682952543
transform 1 0 2260 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_417
timestamp 1682952543
transform 1 0 2300 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_529
timestamp 1682952543
transform 1 0 2300 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_515
timestamp 1682952543
transform 1 0 2316 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_640
timestamp 1682952543
transform 1 0 2292 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1682952543
transform 1 0 2308 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1682952543
transform 1 0 2316 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_566
timestamp 1682952543
transform 1 0 2308 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_438
timestamp 1682952543
transform 1 0 2364 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1682952543
transform 1 0 2420 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_478
timestamp 1682952543
transform 1 0 2404 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_530
timestamp 1682952543
transform 1 0 2364 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1682952543
transform 1 0 2372 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1682952543
transform 1 0 2388 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_516
timestamp 1682952543
transform 1 0 2396 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_533
timestamp 1682952543
transform 1 0 2412 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1682952543
transform 1 0 2428 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_517
timestamp 1682952543
transform 1 0 2436 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_643
timestamp 1682952543
transform 1 0 2364 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_644
timestamp 1682952543
transform 1 0 2380 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1682952543
transform 1 0 2396 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1682952543
transform 1 0 2404 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_647
timestamp 1682952543
transform 1 0 2420 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1682952543
transform 1 0 2436 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_567
timestamp 1682952543
transform 1 0 2356 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1682952543
transform 1 0 2364 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1682952543
transform 1 0 2396 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1682952543
transform 1 0 2404 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_403
timestamp 1682952543
transform 1 0 2460 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_535
timestamp 1682952543
transform 1 0 2508 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1682952543
transform 1 0 2460 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_569
timestamp 1682952543
transform 1 0 2508 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1682952543
transform 1 0 2476 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_536
timestamp 1682952543
transform 1 0 2564 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1682952543
transform 1 0 2596 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_518
timestamp 1682952543
transform 1 0 2604 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_650
timestamp 1682952543
transform 1 0 2572 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1682952543
transform 1 0 2588 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1682952543
transform 1 0 2604 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_570
timestamp 1682952543
transform 1 0 2588 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1682952543
transform 1 0 2572 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_392
timestamp 1682952543
transform 1 0 2636 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1682952543
transform 1 0 2628 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_419
timestamp 1682952543
transform 1 0 2652 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_439
timestamp 1682952543
transform 1 0 2676 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_538
timestamp 1682952543
transform 1 0 2676 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_519
timestamp 1682952543
transform 1 0 2692 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_539
timestamp 1682952543
transform 1 0 2708 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1682952543
transform 1 0 2716 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_653
timestamp 1682952543
transform 1 0 2628 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_571
timestamp 1682952543
transform 1 0 2676 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1682952543
transform 1 0 2668 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_420
timestamp 1682952543
transform 1 0 2740 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1682952543
transform 1 0 2748 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_541
timestamp 1682952543
transform 1 0 2748 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_520
timestamp 1682952543
transform 1 0 2756 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_654
timestamp 1682952543
transform 1 0 2724 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1682952543
transform 1 0 2740 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1682952543
transform 1 0 2756 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1682952543
transform 1 0 2764 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_572
timestamp 1682952543
transform 1 0 2740 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1682952543
transform 1 0 2724 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_393
timestamp 1682952543
transform 1 0 2788 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1682952543
transform 1 0 2772 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_481
timestamp 1682952543
transform 1 0 2836 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_542
timestamp 1682952543
transform 1 0 2772 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1682952543
transform 1 0 2836 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_606
timestamp 1682952543
transform 1 0 2764 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_658
timestamp 1682952543
transform 1 0 2788 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_482
timestamp 1682952543
transform 1 0 2908 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1682952543
transform 1 0 2988 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_544
timestamp 1682952543
transform 1 0 2884 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1682952543
transform 1 0 2892 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1682952543
transform 1 0 2924 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1682952543
transform 1 0 2988 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1682952543
transform 1 0 2972 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_607
timestamp 1682952543
transform 1 0 2980 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1682952543
transform 1 0 3028 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_394
timestamp 1682952543
transform 1 0 3140 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1682952543
transform 1 0 3052 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_406
timestamp 1682952543
transform 1 0 3076 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1682952543
transform 1 0 3116 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_548
timestamp 1682952543
transform 1 0 3012 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_549
timestamp 1682952543
transform 1 0 3028 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_521
timestamp 1682952543
transform 1 0 3036 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_486
timestamp 1682952543
transform 1 0 3148 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_550
timestamp 1682952543
transform 1 0 3100 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1682952543
transform 1 0 3132 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1682952543
transform 1 0 3148 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1682952543
transform 1 0 3164 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_522
timestamp 1682952543
transform 1 0 3172 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_487
timestamp 1682952543
transform 1 0 3276 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1682952543
transform 1 0 3372 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1682952543
transform 1 0 3388 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1682952543
transform 1 0 3300 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_554
timestamp 1682952543
transform 1 0 3236 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_555
timestamp 1682952543
transform 1 0 3268 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1682952543
transform 1 0 3276 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1682952543
transform 1 0 2996 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1682952543
transform 1 0 3004 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1682952543
transform 1 0 3020 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1682952543
transform 1 0 3036 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1682952543
transform 1 0 3052 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1682952543
transform 1 0 3140 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1682952543
transform 1 0 3156 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1682952543
transform 1 0 3172 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1682952543
transform 1 0 3188 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_573
timestamp 1682952543
transform 1 0 3004 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1682952543
transform 1 0 3140 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1682952543
transform 1 0 3188 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1682952543
transform 1 0 3292 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_557
timestamp 1682952543
transform 1 0 3324 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_489
timestamp 1682952543
transform 1 0 3412 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_558
timestamp 1682952543
transform 1 0 3396 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1682952543
transform 1 0 3412 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1682952543
transform 1 0 3428 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_490
timestamp 1682952543
transform 1 0 3436 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_669
timestamp 1682952543
transform 1 0 3372 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_670
timestamp 1682952543
transform 1 0 3388 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_575
timestamp 1682952543
transform 1 0 3340 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1682952543
transform 1 0 3324 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1682952543
transform 1 0 3340 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_538
timestamp 1682952543
transform 1 0 3396 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_671
timestamp 1682952543
transform 1 0 3404 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1682952543
transform 1 0 3420 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_539
timestamp 1682952543
transform 1 0 3428 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_673
timestamp 1682952543
transform 1 0 3436 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_576
timestamp 1682952543
transform 1 0 3420 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1682952543
transform 1 0 3460 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1682952543
transform 1 0 3492 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_441
timestamp 1682952543
transform 1 0 3508 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_524
timestamp 1682952543
transform 1 0 3500 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_561
timestamp 1682952543
transform 1 0 3508 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1682952543
transform 1 0 3460 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_421
timestamp 1682952543
transform 1 0 3580 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1682952543
transform 1 0 3572 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1682952543
transform 1 0 3596 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1682952543
transform 1 0 3564 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_492
timestamp 1682952543
transform 1 0 3612 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_493
timestamp 1682952543
transform 1 0 3636 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_562
timestamp 1682952543
transform 1 0 3564 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1682952543
transform 1 0 3580 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_525
timestamp 1682952543
transform 1 0 3588 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_564
timestamp 1682952543
transform 1 0 3596 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_526
timestamp 1682952543
transform 1 0 3604 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1682952543
transform 1 0 3716 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1682952543
transform 1 0 3692 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1682952543
transform 1 0 3716 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_494
timestamp 1682952543
transform 1 0 3676 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_495
timestamp 1682952543
transform 1 0 3692 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_565
timestamp 1682952543
transform 1 0 3620 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1682952543
transform 1 0 3636 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_527
timestamp 1682952543
transform 1 0 3644 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_567
timestamp 1682952543
transform 1 0 3660 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1682952543
transform 1 0 3676 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1682952543
transform 1 0 3692 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1682952543
transform 1 0 3588 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1682952543
transform 1 0 3604 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1682952543
transform 1 0 3612 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_540
timestamp 1682952543
transform 1 0 3620 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_678
timestamp 1682952543
transform 1 0 3628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1682952543
transform 1 0 3644 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1682952543
transform 1 0 3652 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_541
timestamp 1682952543
transform 1 0 3660 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1682952543
transform 1 0 3708 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_570
timestamp 1682952543
transform 1 0 3716 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_681
timestamp 1682952543
transform 1 0 3668 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1682952543
transform 1 0 3684 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1682952543
transform 1 0 3692 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1682952543
transform 1 0 3708 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_542
timestamp 1682952543
transform 1 0 3716 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1682952543
transform 1 0 3756 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_496
timestamp 1682952543
transform 1 0 3740 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_571
timestamp 1682952543
transform 1 0 3740 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_529
timestamp 1682952543
transform 1 0 3748 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_572
timestamp 1682952543
transform 1 0 3756 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_408
timestamp 1682952543
transform 1 0 3772 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_685
timestamp 1682952543
transform 1 0 3724 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1682952543
transform 1 0 3732 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1682952543
transform 1 0 3748 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1682952543
transform 1 0 3764 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1682952543
transform 1 0 3772 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_577
timestamp 1682952543
transform 1 0 3652 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1682952543
transform 1 0 3692 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1682952543
transform 1 0 3636 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_612
timestamp 1682952543
transform 1 0 3684 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1682952543
transform 1 0 3756 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1682952543
transform 1 0 3724 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_497
timestamp 1682952543
transform 1 0 3796 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_573
timestamp 1682952543
transform 1 0 3796 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_574
timestamp 1682952543
transform 1 0 3812 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1682952543
transform 1 0 3804 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1682952543
transform 1 0 3820 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_580
timestamp 1682952543
transform 1 0 3828 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_575
timestamp 1682952543
transform 1 0 3844 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1682952543
transform 1 0 3868 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1682952543
transform 1 0 3884 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1682952543
transform 1 0 3876 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1682952543
transform 1 0 3892 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_581
timestamp 1682952543
transform 1 0 3876 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_498
timestamp 1682952543
transform 1 0 3924 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_499
timestamp 1682952543
transform 1 0 3940 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_530
timestamp 1682952543
transform 1 0 3916 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_578
timestamp 1682952543
transform 1 0 3924 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1682952543
transform 1 0 3940 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1682952543
transform 1 0 3916 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1682952543
transform 1 0 3932 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_696
timestamp 1682952543
transform 1 0 3948 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_582
timestamp 1682952543
transform 1 0 3916 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1682952543
transform 1 0 3932 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_500
timestamp 1682952543
transform 1 0 4060 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_580
timestamp 1682952543
transform 1 0 3996 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_531
timestamp 1682952543
transform 1 0 4012 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_581
timestamp 1682952543
transform 1 0 4052 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1682952543
transform 1 0 4060 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1682952543
transform 1 0 3972 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_543
timestamp 1682952543
transform 1 0 3996 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1682952543
transform 1 0 4012 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1682952543
transform 1 0 4036 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1682952543
transform 1 0 4084 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_583
timestamp 1682952543
transform 1 0 4084 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1682952543
transform 1 0 4100 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1682952543
transform 1 0 4068 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1682952543
transform 1 0 4076 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_700
timestamp 1682952543
transform 1 0 4092 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1682952543
transform 1 0 4108 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_585
timestamp 1682952543
transform 1 0 4108 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_702
timestamp 1682952543
transform 1 0 4148 0 1 3805
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_6
timestamp 1682952543
transform 1 0 48 0 1 3770
box -10 -3 10 3
use FILL  FILL_127
timestamp 1682952543
transform 1 0 72 0 1 3770
box -8 -3 16 105
use FILL  FILL_128
timestamp 1682952543
transform 1 0 80 0 1 3770
box -8 -3 16 105
use FILL  FILL_129
timestamp 1682952543
transform 1 0 88 0 1 3770
box -8 -3 16 105
use FILL  FILL_130
timestamp 1682952543
transform 1 0 96 0 1 3770
box -8 -3 16 105
use FILL  FILL_131
timestamp 1682952543
transform 1 0 104 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_40
timestamp 1682952543
transform -1 0 128 0 1 3770
box -9 -3 26 105
use FILL  FILL_132
timestamp 1682952543
transform 1 0 128 0 1 3770
box -8 -3 16 105
use FILL  FILL_133
timestamp 1682952543
transform 1 0 136 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_18
timestamp 1682952543
transform -1 0 184 0 1 3770
box -8 -3 46 105
use FILL  FILL_134
timestamp 1682952543
transform 1 0 184 0 1 3770
box -8 -3 16 105
use FILL  FILL_135
timestamp 1682952543
transform 1 0 192 0 1 3770
box -8 -3 16 105
use FILL  FILL_136
timestamp 1682952543
transform 1 0 200 0 1 3770
box -8 -3 16 105
use FILL  FILL_137
timestamp 1682952543
transform 1 0 208 0 1 3770
box -8 -3 16 105
use FILL  FILL_138
timestamp 1682952543
transform 1 0 216 0 1 3770
box -8 -3 16 105
use FILL  FILL_139
timestamp 1682952543
transform 1 0 224 0 1 3770
box -8 -3 16 105
use FILL  FILL_140
timestamp 1682952543
transform 1 0 232 0 1 3770
box -8 -3 16 105
use FILL  FILL_141
timestamp 1682952543
transform 1 0 240 0 1 3770
box -8 -3 16 105
use FILL  FILL_142
timestamp 1682952543
transform 1 0 248 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_41
timestamp 1682952543
transform -1 0 272 0 1 3770
box -9 -3 26 105
use FILL  FILL_143
timestamp 1682952543
transform 1 0 272 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_19
timestamp 1682952543
transform 1 0 280 0 1 3770
box -8 -3 46 105
use FILL  FILL_144
timestamp 1682952543
transform 1 0 320 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_20
timestamp 1682952543
transform 1 0 328 0 1 3770
box -8 -3 46 105
use INVX2  INVX2_42
timestamp 1682952543
transform 1 0 368 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1682952543
transform 1 0 384 0 1 3770
box -8 -3 104 105
use OAI22X1  OAI22X1_30
timestamp 1682952543
transform 1 0 480 0 1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1682952543
transform 1 0 520 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_43
timestamp 1682952543
transform 1 0 616 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1682952543
transform 1 0 632 0 1 3770
box -8 -3 104 105
use FILL  FILL_145
timestamp 1682952543
transform 1 0 728 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_44
timestamp 1682952543
transform 1 0 736 0 1 3770
box -9 -3 26 105
use FILL  FILL_146
timestamp 1682952543
transform 1 0 752 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1682952543
transform -1 0 856 0 1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1682952543
transform -1 0 952 0 1 3770
box -8 -3 104 105
use NOR2X1  NOR2X1_3
timestamp 1682952543
transform 1 0 952 0 1 3770
box -8 -3 32 105
use NOR2X1  NOR2X1_4
timestamp 1682952543
transform 1 0 976 0 1 3770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1682952543
transform 1 0 1000 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_45
timestamp 1682952543
transform -1 0 1112 0 1 3770
box -9 -3 26 105
use FILL  FILL_147
timestamp 1682952543
transform 1 0 1112 0 1 3770
box -8 -3 16 105
use FILL  FILL_148
timestamp 1682952543
transform 1 0 1120 0 1 3770
box -8 -3 16 105
use FILL  FILL_149
timestamp 1682952543
transform 1 0 1128 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_31
timestamp 1682952543
transform -1 0 1176 0 1 3770
box -8 -3 46 105
use FILL  FILL_150
timestamp 1682952543
transform 1 0 1176 0 1 3770
box -8 -3 16 105
use FILL  FILL_151
timestamp 1682952543
transform 1 0 1184 0 1 3770
box -8 -3 16 105
use FILL  FILL_152
timestamp 1682952543
transform 1 0 1192 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_21
timestamp 1682952543
transform 1 0 1200 0 1 3770
box -8 -3 46 105
use NOR2X1  NOR2X1_5
timestamp 1682952543
transform 1 0 1240 0 1 3770
box -8 -3 32 105
use M3_M2  M3_M2_615
timestamp 1682952543
transform 1 0 1276 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_53
timestamp 1682952543
transform 1 0 1264 0 1 3770
box -8 -3 104 105
use FILL  FILL_153
timestamp 1682952543
transform 1 0 1360 0 1 3770
box -8 -3 16 105
use FILL  FILL_154
timestamp 1682952543
transform 1 0 1368 0 1 3770
box -8 -3 16 105
use FILL  FILL_155
timestamp 1682952543
transform 1 0 1376 0 1 3770
box -8 -3 16 105
use FILL  FILL_156
timestamp 1682952543
transform 1 0 1384 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_46
timestamp 1682952543
transform 1 0 1392 0 1 3770
box -9 -3 26 105
use M3_M2  M3_M2_616
timestamp 1682952543
transform 1 0 1452 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_59
timestamp 1682952543
transform -1 0 1504 0 1 3770
box -8 -3 104 105
use AOI22X1  AOI22X1_31
timestamp 1682952543
transform 1 0 1504 0 1 3770
box -8 -3 46 105
use INVX2  INVX2_56
timestamp 1682952543
transform 1 0 1544 0 1 3770
box -9 -3 26 105
use FILL  FILL_178
timestamp 1682952543
transform 1 0 1560 0 1 3770
box -8 -3 16 105
use FILL  FILL_179
timestamp 1682952543
transform 1 0 1568 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_36
timestamp 1682952543
transform 1 0 1576 0 1 3770
box -8 -3 46 105
use AOI22X1  AOI22X1_32
timestamp 1682952543
transform 1 0 1616 0 1 3770
box -8 -3 46 105
use FILL  FILL_180
timestamp 1682952543
transform 1 0 1656 0 1 3770
box -8 -3 16 105
use FILL  FILL_181
timestamp 1682952543
transform 1 0 1664 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_57
timestamp 1682952543
transform 1 0 1672 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1682952543
transform -1 0 1784 0 1 3770
box -8 -3 104 105
use FILL  FILL_182
timestamp 1682952543
transform 1 0 1784 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_33
timestamp 1682952543
transform -1 0 1832 0 1 3770
box -8 -3 46 105
use FILL  FILL_183
timestamp 1682952543
transform 1 0 1832 0 1 3770
box -8 -3 16 105
use FILL  FILL_184
timestamp 1682952543
transform 1 0 1840 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_34
timestamp 1682952543
transform -1 0 1888 0 1 3770
box -8 -3 46 105
use INVX2  INVX2_58
timestamp 1682952543
transform 1 0 1888 0 1 3770
box -9 -3 26 105
use FILL  FILL_185
timestamp 1682952543
transform 1 0 1904 0 1 3770
box -8 -3 16 105
use FILL  FILL_186
timestamp 1682952543
transform 1 0 1912 0 1 3770
box -8 -3 16 105
use FILL  FILL_187
timestamp 1682952543
transform 1 0 1920 0 1 3770
box -8 -3 16 105
use FILL  FILL_188
timestamp 1682952543
transform 1 0 1928 0 1 3770
box -8 -3 16 105
use FILL  FILL_189
timestamp 1682952543
transform 1 0 1936 0 1 3770
box -8 -3 16 105
use FILL  FILL_190
timestamp 1682952543
transform 1 0 1944 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1682952543
transform -1 0 2048 0 1 3770
box -8 -3 104 105
use FILL  FILL_191
timestamp 1682952543
transform 1 0 2048 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_617
timestamp 1682952543
transform 1 0 2068 0 1 3775
box -3 -3 3 3
use FILL  FILL_192
timestamp 1682952543
transform 1 0 2056 0 1 3770
box -8 -3 16 105
use FILL  FILL_193
timestamp 1682952543
transform 1 0 2064 0 1 3770
box -8 -3 16 105
use FILL  FILL_194
timestamp 1682952543
transform 1 0 2072 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_618
timestamp 1682952543
transform 1 0 2092 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_62
timestamp 1682952543
transform 1 0 2080 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_59
timestamp 1682952543
transform 1 0 2176 0 1 3770
box -9 -3 26 105
use FILL  FILL_195
timestamp 1682952543
transform 1 0 2192 0 1 3770
box -8 -3 16 105
use FILL  FILL_196
timestamp 1682952543
transform 1 0 2200 0 1 3770
box -8 -3 16 105
use FILL  FILL_197
timestamp 1682952543
transform 1 0 2208 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_37
timestamp 1682952543
transform 1 0 2216 0 1 3770
box -8 -3 46 105
use FILL  FILL_198
timestamp 1682952543
transform 1 0 2256 0 1 3770
box -8 -3 16 105
use FILL  FILL_207
timestamp 1682952543
transform 1 0 2264 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_39
timestamp 1682952543
transform 1 0 2272 0 1 3770
box -8 -3 46 105
use FILL  FILL_209
timestamp 1682952543
transform 1 0 2312 0 1 3770
box -8 -3 16 105
use FILL  FILL_210
timestamp 1682952543
transform 1 0 2320 0 1 3770
box -8 -3 16 105
use FILL  FILL_215
timestamp 1682952543
transform 1 0 2328 0 1 3770
box -8 -3 16 105
use FILL  FILL_217
timestamp 1682952543
transform 1 0 2336 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_62
timestamp 1682952543
transform 1 0 2344 0 1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_40
timestamp 1682952543
transform 1 0 2360 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_42
timestamp 1682952543
transform 1 0 2400 0 1 3770
box -8 -3 46 105
use FILL  FILL_221
timestamp 1682952543
transform 1 0 2440 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1682952543
transform 1 0 2448 0 1 3770
box -8 -3 104 105
use M3_M2  M3_M2_619
timestamp 1682952543
transform 1 0 2556 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1682952543
transform 1 0 2572 0 1 3775
box -3 -3 3 3
use INVX2  INVX2_63
timestamp 1682952543
transform 1 0 2544 0 1 3770
box -9 -3 26 105
use FILL  FILL_222
timestamp 1682952543
transform 1 0 2560 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_43
timestamp 1682952543
transform 1 0 2568 0 1 3770
box -8 -3 46 105
use FILL  FILL_223
timestamp 1682952543
transform 1 0 2608 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_621
timestamp 1682952543
transform 1 0 2652 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_622
timestamp 1682952543
transform 1 0 2684 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_71
timestamp 1682952543
transform 1 0 2616 0 1 3770
box -8 -3 104 105
use FILL  FILL_224
timestamp 1682952543
transform 1 0 2712 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_623
timestamp 1682952543
transform 1 0 2756 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_44
timestamp 1682952543
transform 1 0 2720 0 1 3770
box -8 -3 46 105
use M3_M2  M3_M2_624
timestamp 1682952543
transform 1 0 2772 0 1 3775
box -3 -3 3 3
use INVX2  INVX2_64
timestamp 1682952543
transform 1 0 2760 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1682952543
transform 1 0 2776 0 1 3770
box -8 -3 104 105
use M3_M2  M3_M2_625
timestamp 1682952543
transform 1 0 2900 0 1 3775
box -3 -3 3 3
use INVX2  INVX2_65
timestamp 1682952543
transform 1 0 2872 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1682952543
transform -1 0 2984 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_66
timestamp 1682952543
transform -1 0 3000 0 1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_45
timestamp 1682952543
transform -1 0 3040 0 1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1682952543
transform 1 0 3040 0 1 3770
box -8 -3 104 105
use OAI22X1  OAI22X1_46
timestamp 1682952543
transform -1 0 3176 0 1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_75
timestamp 1682952543
transform 1 0 3176 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_67
timestamp 1682952543
transform -1 0 3288 0 1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1682952543
transform -1 0 3384 0 1 3770
box -8 -3 104 105
use M3_M2  M3_M2_626
timestamp 1682952543
transform 1 0 3412 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_47
timestamp 1682952543
transform 1 0 3384 0 1 3770
box -8 -3 46 105
use INVX2  INVX2_68
timestamp 1682952543
transform -1 0 3440 0 1 3770
box -9 -3 26 105
use M3_M2  M3_M2_627
timestamp 1682952543
transform 1 0 3452 0 1 3775
box -3 -3 3 3
use FILL  FILL_225
timestamp 1682952543
transform 1 0 3440 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_628
timestamp 1682952543
transform 1 0 3516 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_77
timestamp 1682952543
transform 1 0 3448 0 1 3770
box -8 -3 104 105
use FILL  FILL_226
timestamp 1682952543
transform 1 0 3544 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_69
timestamp 1682952543
transform 1 0 3552 0 1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_48
timestamp 1682952543
transform 1 0 3568 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_49
timestamp 1682952543
transform 1 0 3608 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_50
timestamp 1682952543
transform 1 0 3648 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_51
timestamp 1682952543
transform 1 0 3688 0 1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_69
timestamp 1682952543
transform 1 0 3728 0 1 3770
box -8 -3 46 105
use FILL  FILL_256
timestamp 1682952543
transform 1 0 3768 0 1 3770
box -8 -3 16 105
use FILL  FILL_257
timestamp 1682952543
transform 1 0 3776 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_71
timestamp 1682952543
transform -1 0 3824 0 1 3770
box -8 -3 46 105
use FILL  FILL_258
timestamp 1682952543
transform 1 0 3824 0 1 3770
box -8 -3 16 105
use FILL  FILL_259
timestamp 1682952543
transform 1 0 3832 0 1 3770
box -8 -3 16 105
use FILL  FILL_260
timestamp 1682952543
transform 1 0 3840 0 1 3770
box -8 -3 16 105
use FILL  FILL_261
timestamp 1682952543
transform 1 0 3848 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_72
timestamp 1682952543
transform 1 0 3856 0 1 3770
box -8 -3 46 105
use FILL  FILL_262
timestamp 1682952543
transform 1 0 3896 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_629
timestamp 1682952543
transform 1 0 3916 0 1 3775
box -3 -3 3 3
use FILL  FILL_263
timestamp 1682952543
transform 1 0 3904 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_73
timestamp 1682952543
transform -1 0 3952 0 1 3770
box -8 -3 46 105
use M3_M2  M3_M2_630
timestamp 1682952543
transform 1 0 3972 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1682952543
transform 1 0 4004 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_632
timestamp 1682952543
transform 1 0 4028 0 1 3775
box -3 -3 3 3
use FILL  FILL_264
timestamp 1682952543
transform 1 0 3952 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1682952543
transform 1 0 3960 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_78
timestamp 1682952543
transform -1 0 4072 0 1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_74
timestamp 1682952543
transform -1 0 4112 0 1 3770
box -8 -3 46 105
use FILL  FILL_265
timestamp 1682952543
transform 1 0 4112 0 1 3770
box -8 -3 16 105
use FILL  FILL_266
timestamp 1682952543
transform 1 0 4120 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_79
timestamp 1682952543
transform -1 0 4144 0 1 3770
box -9 -3 26 105
use FILL  FILL_267
timestamp 1682952543
transform 1 0 4144 0 1 3770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_7
timestamp 1682952543
transform 1 0 4177 0 1 3770
box -10 -3 10 3
use M3_M2  M3_M2_633
timestamp 1682952543
transform 1 0 108 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1682952543
transform 1 0 180 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1682952543
transform 1 0 164 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_664
timestamp 1682952543
transform 1 0 180 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1682952543
transform 1 0 156 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_707
timestamp 1682952543
transform 1 0 84 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1682952543
transform 1 0 172 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1682952543
transform 1 0 180 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1682952543
transform 1 0 196 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1682952543
transform 1 0 132 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_853
timestamp 1682952543
transform 1 0 164 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_785
timestamp 1682952543
transform 1 0 172 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1682952543
transform 1 0 220 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1682952543
transform 1 0 244 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1682952543
transform 1 0 268 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1682952543
transform 1 0 236 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_711
timestamp 1682952543
transform 1 0 220 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_704
timestamp 1682952543
transform 1 0 348 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_712
timestamp 1682952543
transform 1 0 324 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1682952543
transform 1 0 332 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1682952543
transform 1 0 348 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1682952543
transform 1 0 364 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_854
timestamp 1682952543
transform 1 0 188 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_855
timestamp 1682952543
transform 1 0 204 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1682952543
transform 1 0 132 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1682952543
transform 1 0 172 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1682952543
transform 1 0 196 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1682952543
transform 1 0 220 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_856
timestamp 1682952543
transform 1 0 260 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_787
timestamp 1682952543
transform 1 0 292 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_857
timestamp 1682952543
transform 1 0 300 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1682952543
transform 1 0 308 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1682952543
transform 1 0 316 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1682952543
transform 1 0 340 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_788
timestamp 1682952543
transform 1 0 348 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_861
timestamp 1682952543
transform 1 0 356 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_811
timestamp 1682952543
transform 1 0 244 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1682952543
transform 1 0 260 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_813
timestamp 1682952543
transform 1 0 308 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1682952543
transform 1 0 324 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1682952543
transform 1 0 340 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1682952543
transform 1 0 204 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_859
timestamp 1682952543
transform 1 0 316 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1682952543
transform 1 0 388 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_665
timestamp 1682952543
transform 1 0 476 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_705
timestamp 1682952543
transform 1 0 508 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_716
timestamp 1682952543
transform 1 0 388 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1682952543
transform 1 0 476 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1682952543
transform 1 0 492 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1682952543
transform 1 0 508 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1682952543
transform 1 0 516 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1682952543
transform 1 0 372 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1682952543
transform 1 0 412 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1682952543
transform 1 0 476 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1682952543
transform 1 0 484 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_816
timestamp 1682952543
transform 1 0 372 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1682952543
transform 1 0 412 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1682952543
transform 1 0 492 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_866
timestamp 1682952543
transform 1 0 500 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_706
timestamp 1682952543
transform 1 0 540 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1682952543
transform 1 0 532 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_721
timestamp 1682952543
transform 1 0 540 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1682952543
transform 1 0 524 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1682952543
transform 1 0 532 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1682952543
transform 1 0 548 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_818
timestamp 1682952543
transform 1 0 516 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1682952543
transform 1 0 548 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_870
timestamp 1682952543
transform 1 0 572 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_707
timestamp 1682952543
transform 1 0 588 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_708
timestamp 1682952543
transform 1 0 620 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1682952543
transform 1 0 740 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1682952543
transform 1 0 740 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_709
timestamp 1682952543
transform 1 0 724 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_722
timestamp 1682952543
transform 1 0 580 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1682952543
transform 1 0 588 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1682952543
transform 1 0 596 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1682952543
transform 1 0 620 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1682952543
transform 1 0 636 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_727
timestamp 1682952543
transform 1 0 724 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1682952543
transform 1 0 740 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_820
timestamp 1682952543
transform 1 0 572 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_871
timestamp 1682952543
transform 1 0 588 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1682952543
transform 1 0 604 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1682952543
transform 1 0 620 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1682952543
transform 1 0 660 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_875
timestamp 1682952543
transform 1 0 716 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1682952543
transform 1 0 732 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1682952543
transform 1 0 748 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_860
timestamp 1682952543
transform 1 0 588 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1682952543
transform 1 0 620 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1682952543
transform 1 0 620 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_880
timestamp 1682952543
transform 1 0 652 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_878
timestamp 1682952543
transform 1 0 764 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1682952543
transform 1 0 772 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_822
timestamp 1682952543
transform 1 0 764 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1682952543
transform 1 0 804 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1682952543
transform 1 0 788 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_729
timestamp 1682952543
transform 1 0 788 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1682952543
transform 1 0 796 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1682952543
transform 1 0 812 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_765
timestamp 1682952543
transform 1 0 820 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_880
timestamp 1682952543
transform 1 0 804 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1682952543
transform 1 0 820 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1682952543
transform 1 0 828 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_823
timestamp 1682952543
transform 1 0 828 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1682952543
transform 1 0 812 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_896
timestamp 1682952543
transform 1 0 820 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_711
timestamp 1682952543
transform 1 0 844 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_732
timestamp 1682952543
transform 1 0 844 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_733
timestamp 1682952543
transform 1 0 860 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_734
timestamp 1682952543
transform 1 0 884 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1682952543
transform 1 0 892 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1682952543
transform 1 0 876 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1682952543
transform 1 0 892 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_862
timestamp 1682952543
transform 1 0 884 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1682952543
transform 1 0 892 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_667
timestamp 1682952543
transform 1 0 924 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_706
timestamp 1682952543
transform 1 0 924 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1682952543
transform 1 0 916 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_790
timestamp 1682952543
transform 1 0 924 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_736
timestamp 1682952543
transform 1 0 932 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_641
timestamp 1682952543
transform 1 0 988 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1682952543
transform 1 0 1076 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_668
timestamp 1682952543
transform 1 0 972 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_669
timestamp 1682952543
transform 1 0 1044 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1682952543
transform 1 0 1060 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1682952543
transform 1 0 980 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1682952543
transform 1 0 1012 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_737
timestamp 1682952543
transform 1 0 980 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_671
timestamp 1682952543
transform 1 0 1108 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1682952543
transform 1 0 1084 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_738
timestamp 1682952543
transform 1 0 1084 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1682952543
transform 1 0 1092 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_740
timestamp 1682952543
transform 1 0 1108 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1682952543
transform 1 0 964 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1682952543
transform 1 0 1020 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1682952543
transform 1 0 1060 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1682952543
transform 1 0 1068 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1682952543
transform 1 0 1084 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1682952543
transform 1 0 1100 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_824
timestamp 1682952543
transform 1 0 1020 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1682952543
transform 1 0 1068 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_863
timestamp 1682952543
transform 1 0 964 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1682952543
transform 1 0 1108 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_897
timestamp 1682952543
transform 1 0 1084 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_892
timestamp 1682952543
transform 1 0 1124 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_643
timestamp 1682952543
transform 1 0 1164 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1682952543
transform 1 0 1156 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1682952543
transform 1 0 1140 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1682952543
transform 1 0 1204 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1682952543
transform 1 0 1196 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_741
timestamp 1682952543
transform 1 0 1148 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_742
timestamp 1682952543
transform 1 0 1164 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1682952543
transform 1 0 1172 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1682952543
transform 1 0 1188 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1682952543
transform 1 0 1140 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1682952543
transform 1 0 1164 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_792
timestamp 1682952543
transform 1 0 1172 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_895
timestamp 1682952543
transform 1 0 1180 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1682952543
transform 1 0 1196 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_826
timestamp 1682952543
transform 1 0 1164 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_827
timestamp 1682952543
transform 1 0 1196 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_864
timestamp 1682952543
transform 1 0 1188 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_745
timestamp 1682952543
transform 1 0 1212 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_793
timestamp 1682952543
transform 1 0 1212 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_716
timestamp 1682952543
transform 1 0 1228 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_746
timestamp 1682952543
transform 1 0 1220 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_767
timestamp 1682952543
transform 1 0 1244 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_747
timestamp 1682952543
transform 1 0 1252 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1682952543
transform 1 0 1244 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_717
timestamp 1682952543
transform 1 0 1292 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_748
timestamp 1682952543
transform 1 0 1276 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_749
timestamp 1682952543
transform 1 0 1292 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_768
timestamp 1682952543
transform 1 0 1300 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_750
timestamp 1682952543
transform 1 0 1308 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1682952543
transform 1 0 1260 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_899
timestamp 1682952543
transform 1 0 1268 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1682952543
transform 1 0 1284 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_828
timestamp 1682952543
transform 1 0 1252 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1682952543
transform 1 0 1284 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_865
timestamp 1682952543
transform 1 0 1268 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_898
timestamp 1682952543
transform 1 0 1276 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1682952543
transform 1 0 1308 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_901
timestamp 1682952543
transform 1 0 1324 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1682952543
transform 1 0 1332 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1682952543
transform 1 0 1340 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_866
timestamp 1682952543
transform 1 0 1332 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_751
timestamp 1682952543
transform 1 0 1380 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1682952543
transform 1 0 1388 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1682952543
transform 1 0 1372 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_794
timestamp 1682952543
transform 1 0 1380 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_905
timestamp 1682952543
transform 1 0 1388 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1682952543
transform 1 0 1492 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1682952543
transform 1 0 1404 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1682952543
transform 1 0 1412 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_795
timestamp 1682952543
transform 1 0 1420 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_908
timestamp 1682952543
transform 1 0 1444 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1682952543
transform 1 0 1508 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_830
timestamp 1682952543
transform 1 0 1404 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1682952543
transform 1 0 1444 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1682952543
transform 1 0 1524 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_754
timestamp 1682952543
transform 1 0 1524 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_883
timestamp 1682952543
transform 1 0 1516 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_718
timestamp 1682952543
transform 1 0 1620 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_755
timestamp 1682952543
transform 1 0 1620 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1682952543
transform 1 0 1532 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1682952543
transform 1 0 1572 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_899
timestamp 1682952543
transform 1 0 1524 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_884
timestamp 1682952543
transform 1 0 1548 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_900
timestamp 1682952543
transform 1 0 1548 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_912
timestamp 1682952543
transform 1 0 1636 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1682952543
transform 1 0 1724 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_756
timestamp 1682952543
transform 1 0 1724 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_645
timestamp 1682952543
transform 1 0 1812 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1682952543
transform 1 0 1836 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_674
timestamp 1682952543
transform 1 0 1780 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_720
timestamp 1682952543
transform 1 0 1772 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_757
timestamp 1682952543
transform 1 0 1820 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_758
timestamp 1682952543
transform 1 0 1836 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1682952543
transform 1 0 1676 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1682952543
transform 1 0 1740 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1682952543
transform 1 0 1796 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1682952543
transform 1 0 1836 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_832
timestamp 1682952543
transform 1 0 1796 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1682952543
transform 1 0 1836 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_675
timestamp 1682952543
transform 1 0 1852 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_721
timestamp 1682952543
transform 1 0 1876 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1682952543
transform 1 0 1924 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1682952543
transform 1 0 1940 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_759
timestamp 1682952543
transform 1 0 1940 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_676
timestamp 1682952543
transform 1 0 2052 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1682952543
transform 1 0 1972 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1682952543
transform 1 0 2036 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_760
timestamp 1682952543
transform 1 0 2036 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1682952543
transform 1 0 1860 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1682952543
transform 1 0 1916 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_919
timestamp 1682952543
transform 1 0 1956 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1682952543
transform 1 0 2004 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_677
timestamp 1682952543
transform 1 0 2140 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_726
timestamp 1682952543
transform 1 0 2108 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_761
timestamp 1682952543
transform 1 0 2060 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1682952543
transform 1 0 2108 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1682952543
transform 1 0 2204 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_728
timestamp 1682952543
transform 1 0 2228 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_762
timestamp 1682952543
transform 1 0 2188 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1682952543
transform 1 0 2204 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1682952543
transform 1 0 2220 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_922
timestamp 1682952543
transform 1 0 2196 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1682952543
transform 1 0 2212 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1682952543
transform 1 0 2228 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_834
timestamp 1682952543
transform 1 0 2212 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1682952543
transform 1 0 2196 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1682952543
transform 1 0 2244 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1682952543
transform 1 0 2252 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1682952543
transform 1 0 2276 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_678
timestamp 1682952543
transform 1 0 2332 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1682952543
transform 1 0 2348 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_766
timestamp 1682952543
transform 1 0 2340 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1682952543
transform 1 0 2348 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_679
timestamp 1682952543
transform 1 0 2380 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_680
timestamp 1682952543
transform 1 0 2396 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_770
timestamp 1682952543
transform 1 0 2372 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1682952543
transform 1 0 2404 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_768
timestamp 1682952543
transform 1 0 2380 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1682952543
transform 1 0 2396 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1682952543
transform 1 0 2404 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1682952543
transform 1 0 2372 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1682952543
transform 1 0 2388 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_885
timestamp 1682952543
transform 1 0 2388 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1682952543
transform 1 0 2412 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_928
timestamp 1682952543
transform 1 0 2412 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_647
timestamp 1682952543
transform 1 0 2460 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1682952543
transform 1 0 2452 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_771
timestamp 1682952543
transform 1 0 2436 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_772
timestamp 1682952543
transform 1 0 2452 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_773
timestamp 1682952543
transform 1 0 2460 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1682952543
transform 1 0 2444 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_835
timestamp 1682952543
transform 1 0 2444 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_772
timestamp 1682952543
transform 1 0 2468 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_774
timestamp 1682952543
transform 1 0 2484 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_648
timestamp 1682952543
transform 1 0 2516 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_649
timestamp 1682952543
transform 1 0 2540 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_731
timestamp 1682952543
transform 1 0 2508 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_732
timestamp 1682952543
transform 1 0 2548 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1682952543
transform 1 0 2580 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1682952543
transform 1 0 2596 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_733
timestamp 1682952543
transform 1 0 2564 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_775
timestamp 1682952543
transform 1 0 2508 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1682952543
transform 1 0 2516 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1682952543
transform 1 0 2532 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_778
timestamp 1682952543
transform 1 0 2548 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1682952543
transform 1 0 2468 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1682952543
transform 1 0 2492 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_796
timestamp 1682952543
transform 1 0 2500 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_932
timestamp 1682952543
transform 1 0 2508 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_836
timestamp 1682952543
transform 1 0 2492 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_868
timestamp 1682952543
transform 1 0 2460 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_933
timestamp 1682952543
transform 1 0 2524 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1682952543
transform 1 0 2540 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_869
timestamp 1682952543
transform 1 0 2524 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1682952543
transform 1 0 2540 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_901
timestamp 1682952543
transform 1 0 2540 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1682952543
transform 1 0 2556 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1682952543
transform 1 0 2636 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1682952543
transform 1 0 2604 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_779
timestamp 1682952543
transform 1 0 2564 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1682952543
transform 1 0 2580 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_781
timestamp 1682952543
transform 1 0 2596 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1682952543
transform 1 0 2604 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1682952543
transform 1 0 2556 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1682952543
transform 1 0 2588 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_837
timestamp 1682952543
transform 1 0 2588 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_937
timestamp 1682952543
transform 1 0 2604 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_870
timestamp 1682952543
transform 1 0 2596 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_902
timestamp 1682952543
transform 1 0 2572 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1682952543
transform 1 0 2644 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1682952543
transform 1 0 2652 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1682952543
transform 1 0 2620 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_783
timestamp 1682952543
transform 1 0 2628 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1682952543
transform 1 0 2644 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_785
timestamp 1682952543
transform 1 0 2652 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1682952543
transform 1 0 2668 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1682952543
transform 1 0 2636 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_797
timestamp 1682952543
transform 1 0 2644 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_939
timestamp 1682952543
transform 1 0 2652 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1682952543
transform 1 0 2676 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_838
timestamp 1682952543
transform 1 0 2636 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1682952543
transform 1 0 2676 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1682952543
transform 1 0 2724 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_787
timestamp 1682952543
transform 1 0 2708 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1682952543
transform 1 0 2716 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_839
timestamp 1682952543
transform 1 0 2692 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1682952543
transform 1 0 2732 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1682952543
transform 1 0 2756 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_789
timestamp 1682952543
transform 1 0 2740 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1682952543
transform 1 0 2756 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1682952543
transform 1 0 2732 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1682952543
transform 1 0 2748 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_887
timestamp 1682952543
transform 1 0 2748 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1682952543
transform 1 0 2764 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_652
timestamp 1682952543
transform 1 0 2812 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1682952543
transform 1 0 2788 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1682952543
transform 1 0 2788 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1682952543
transform 1 0 2804 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1682952543
transform 1 0 2796 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_944
timestamp 1682952543
transform 1 0 2812 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_653
timestamp 1682952543
transform 1 0 2844 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1682952543
transform 1 0 2852 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1682952543
transform 1 0 2828 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_793
timestamp 1682952543
transform 1 0 2828 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1682952543
transform 1 0 2892 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1682952543
transform 1 0 2884 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1682952543
transform 1 0 2900 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1682952543
transform 1 0 2924 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_690
timestamp 1682952543
transform 1 0 2964 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_739
timestamp 1682952543
transform 1 0 2884 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1682952543
transform 1 0 2900 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_741
timestamp 1682952543
transform 1 0 2932 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_742
timestamp 1682952543
transform 1 0 2948 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_794
timestamp 1682952543
transform 1 0 2844 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1682952543
transform 1 0 2852 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1682952543
transform 1 0 2868 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1682952543
transform 1 0 2884 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1682952543
transform 1 0 2892 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1682952543
transform 1 0 2908 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1682952543
transform 1 0 2924 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1682952543
transform 1 0 2932 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1682952543
transform 1 0 2948 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1682952543
transform 1 0 2844 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1682952543
transform 1 0 2876 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1682952543
transform 1 0 2892 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_840
timestamp 1682952543
transform 1 0 2844 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_903
timestamp 1682952543
transform 1 0 2828 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_872
timestamp 1682952543
transform 1 0 2876 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1682952543
transform 1 0 2908 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_775
timestamp 1682952543
transform 1 0 2956 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_743
timestamp 1682952543
transform 1 0 3004 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_803
timestamp 1682952543
transform 1 0 2964 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1682952543
transform 1 0 2980 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1682952543
transform 1 0 2916 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1682952543
transform 1 0 2932 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_799
timestamp 1682952543
transform 1 0 2940 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_950
timestamp 1682952543
transform 1 0 2956 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_841
timestamp 1682952543
transform 1 0 2932 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1682952543
transform 1 0 2900 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_873
timestamp 1682952543
transform 1 0 2948 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1682952543
transform 1 0 3012 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_805
timestamp 1682952543
transform 1 0 3076 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1682952543
transform 1 0 3084 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_951
timestamp 1682952543
transform 1 0 3004 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1682952543
transform 1 0 3060 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1682952543
transform 1 0 3068 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_842
timestamp 1682952543
transform 1 0 3068 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1682952543
transform 1 0 2980 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1682952543
transform 1 0 3084 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_890
timestamp 1682952543
transform 1 0 3084 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_691
timestamp 1682952543
transform 1 0 3140 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_744
timestamp 1682952543
transform 1 0 3132 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_807
timestamp 1682952543
transform 1 0 3116 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1682952543
transform 1 0 3108 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1682952543
transform 1 0 3124 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1682952543
transform 1 0 3140 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1682952543
transform 1 0 3148 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_745
timestamp 1682952543
transform 1 0 3172 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_809
timestamp 1682952543
transform 1 0 3172 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1682952543
transform 1 0 3180 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_801
timestamp 1682952543
transform 1 0 3180 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1682952543
transform 1 0 3220 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1682952543
transform 1 0 3252 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_811
timestamp 1682952543
transform 1 0 3220 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1682952543
transform 1 0 3236 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_777
timestamp 1682952543
transform 1 0 3244 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_813
timestamp 1682952543
transform 1 0 3252 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1682952543
transform 1 0 3228 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1682952543
transform 1 0 3244 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_746
timestamp 1682952543
transform 1 0 3268 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_959
timestamp 1682952543
transform 1 0 3268 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_747
timestamp 1682952543
transform 1 0 3292 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1682952543
transform 1 0 3284 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_814
timestamp 1682952543
transform 1 0 3292 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_843
timestamp 1682952543
transform 1 0 3292 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1682952543
transform 1 0 3316 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_815
timestamp 1682952543
transform 1 0 3316 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1682952543
transform 1 0 3332 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1682952543
transform 1 0 3348 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1682952543
transform 1 0 3316 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_802
timestamp 1682952543
transform 1 0 3324 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_961
timestamp 1682952543
transform 1 0 3340 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_874
timestamp 1682952543
transform 1 0 3316 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1682952543
transform 1 0 3396 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_818
timestamp 1682952543
transform 1 0 3380 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1682952543
transform 1 0 3396 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1682952543
transform 1 0 3372 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1682952543
transform 1 0 3388 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_844
timestamp 1682952543
transform 1 0 3388 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_891
timestamp 1682952543
transform 1 0 3388 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1682952543
transform 1 0 3468 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_820
timestamp 1682952543
transform 1 0 3420 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1682952543
transform 1 0 3420 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_964
timestamp 1682952543
transform 1 0 3468 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_693
timestamp 1682952543
transform 1 0 3516 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_656
timestamp 1682952543
transform 1 0 3556 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_751
timestamp 1682952543
transform 1 0 3540 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_657
timestamp 1682952543
transform 1 0 3676 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_694
timestamp 1682952543
transform 1 0 3676 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1682952543
transform 1 0 3588 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1682952543
transform 1 0 3636 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_821
timestamp 1682952543
transform 1 0 3524 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1682952543
transform 1 0 3540 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1682952543
transform 1 0 3556 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1682952543
transform 1 0 3516 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1682952543
transform 1 0 3532 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_804
timestamp 1682952543
transform 1 0 3540 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_824
timestamp 1682952543
transform 1 0 3588 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_779
timestamp 1682952543
transform 1 0 3660 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_967
timestamp 1682952543
transform 1 0 3548 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1682952543
transform 1 0 3556 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1682952543
transform 1 0 3572 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1682952543
transform 1 0 3636 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_845
timestamp 1682952543
transform 1 0 3516 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1682952543
transform 1 0 3548 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_875
timestamp 1682952543
transform 1 0 3620 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_892
timestamp 1682952543
transform 1 0 3572 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1682952543
transform 1 0 3708 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1682952543
transform 1 0 3756 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_696
timestamp 1682952543
transform 1 0 3756 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1682952543
transform 1 0 3708 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1682952543
transform 1 0 3724 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_756
timestamp 1682952543
transform 1 0 3748 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_825
timestamp 1682952543
transform 1 0 3692 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1682952543
transform 1 0 3708 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1682952543
transform 1 0 3724 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1682952543
transform 1 0 3732 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_780
timestamp 1682952543
transform 1 0 3740 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1682952543
transform 1 0 3780 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_829
timestamp 1682952543
transform 1 0 3748 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1682952543
transform 1 0 3764 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1682952543
transform 1 0 3772 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_971
timestamp 1682952543
transform 1 0 3700 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1682952543
transform 1 0 3716 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_805
timestamp 1682952543
transform 1 0 3724 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_973
timestamp 1682952543
transform 1 0 3732 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1682952543
transform 1 0 3756 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_847
timestamp 1682952543
transform 1 0 3684 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_848
timestamp 1682952543
transform 1 0 3700 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_849
timestamp 1682952543
transform 1 0 3740 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_876
timestamp 1682952543
transform 1 0 3732 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1682952543
transform 1 0 3844 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1682952543
transform 1 0 3836 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_832
timestamp 1682952543
transform 1 0 3804 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_781
timestamp 1682952543
transform 1 0 3812 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1682952543
transform 1 0 3892 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1682952543
transform 1 0 3916 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_660
timestamp 1682952543
transform 1 0 3964 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_700
timestamp 1682952543
transform 1 0 3956 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_758
timestamp 1682952543
transform 1 0 3868 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1682952543
transform 1 0 3884 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_760
timestamp 1682952543
transform 1 0 3924 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1682952543
transform 1 0 3940 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_833
timestamp 1682952543
transform 1 0 3820 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1682952543
transform 1 0 3836 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_835
timestamp 1682952543
transform 1 0 3844 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1682952543
transform 1 0 3860 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1682952543
transform 1 0 3780 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_806
timestamp 1682952543
transform 1 0 3796 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_782
timestamp 1682952543
transform 1 0 3868 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_837
timestamp 1682952543
transform 1 0 3876 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1682952543
transform 1 0 3884 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1682952543
transform 1 0 3900 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_783
timestamp 1682952543
transform 1 0 3908 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_840
timestamp 1682952543
transform 1 0 3916 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1682952543
transform 1 0 3924 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1682952543
transform 1 0 3940 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1682952543
transform 1 0 3956 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1682952543
transform 1 0 3964 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1682952543
transform 1 0 3980 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1682952543
transform 1 0 3804 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_977
timestamp 1682952543
transform 1 0 3812 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1682952543
transform 1 0 3828 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1682952543
transform 1 0 3844 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1682952543
transform 1 0 3852 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_981
timestamp 1682952543
transform 1 0 3868 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_993
timestamp 1682952543
transform 1 0 3796 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_807
timestamp 1682952543
transform 1 0 3876 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_982
timestamp 1682952543
transform 1 0 3884 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1682952543
transform 1 0 3908 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_784
timestamp 1682952543
transform 1 0 3988 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1682952543
transform 1 0 4036 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_662
timestamp 1682952543
transform 1 0 4076 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1682952543
transform 1 0 4020 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1682952543
transform 1 0 4092 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_763
timestamp 1682952543
transform 1 0 4076 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_846
timestamp 1682952543
transform 1 0 3996 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1682952543
transform 1 0 4004 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1682952543
transform 1 0 4020 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1682952543
transform 1 0 4036 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1682952543
transform 1 0 4052 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_984
timestamp 1682952543
transform 1 0 3932 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1682952543
transform 1 0 3948 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1682952543
transform 1 0 3964 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_987
timestamp 1682952543
transform 1 0 3988 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1682952543
transform 1 0 4004 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1682952543
transform 1 0 4028 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_850
timestamp 1682952543
transform 1 0 3844 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1682952543
transform 1 0 3884 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_852
timestamp 1682952543
transform 1 0 3900 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_853
timestamp 1682952543
transform 1 0 3924 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1682952543
transform 1 0 3948 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1682952543
transform 1 0 3804 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_893
timestamp 1682952543
transform 1 0 3812 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_905
timestamp 1682952543
transform 1 0 3796 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_906
timestamp 1682952543
transform 1 0 3852 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_907
timestamp 1682952543
transform 1 0 3900 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1682952543
transform 1 0 3988 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_856
timestamp 1682952543
transform 1 0 4004 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1682952543
transform 1 0 3996 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_894
timestamp 1682952543
transform 1 0 3932 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_895
timestamp 1682952543
transform 1 0 3964 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1682952543
transform 1 0 3972 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_851
timestamp 1682952543
transform 1 0 4148 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1682952543
transform 1 0 4076 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_991
timestamp 1682952543
transform 1 0 4132 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_992
timestamp 1682952543
transform 1 0 4140 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_857
timestamp 1682952543
transform 1 0 4140 0 1 3715
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_8
timestamp 1682952543
transform 1 0 24 0 1 3670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_54
timestamp 1682952543
transform 1 0 72 0 -1 3770
box -8 -3 104 105
use AOI22X1  AOI22X1_22
timestamp 1682952543
transform -1 0 208 0 -1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1682952543
transform 1 0 208 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_47
timestamp 1682952543
transform -1 0 320 0 -1 3770
box -9 -3 26 105
use AOI22X1  AOI22X1_23
timestamp 1682952543
transform 1 0 320 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_48
timestamp 1682952543
transform 1 0 360 0 -1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1682952543
transform 1 0 376 0 -1 3770
box -8 -3 104 105
use OAI22X1  OAI22X1_32
timestamp 1682952543
transform 1 0 472 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_49
timestamp 1682952543
transform 1 0 512 0 -1 3770
box -9 -3 26 105
use AOI22X1  AOI22X1_24
timestamp 1682952543
transform 1 0 528 0 -1 3770
box -8 -3 46 105
use FILL  FILL_157
timestamp 1682952543
transform 1 0 568 0 -1 3770
box -8 -3 16 105
use FILL  FILL_158
timestamp 1682952543
transform 1 0 576 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_25
timestamp 1682952543
transform 1 0 584 0 -1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1682952543
transform 1 0 624 0 -1 3770
box -8 -3 104 105
use OAI22X1  OAI22X1_33
timestamp 1682952543
transform 1 0 720 0 -1 3770
box -8 -3 46 105
use FILL  FILL_159
timestamp 1682952543
transform 1 0 760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_160
timestamp 1682952543
transform 1 0 768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_161
timestamp 1682952543
transform 1 0 776 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_26
timestamp 1682952543
transform -1 0 824 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_50
timestamp 1682952543
transform 1 0 824 0 -1 3770
box -9 -3 26 105
use FILL  FILL_162
timestamp 1682952543
transform 1 0 840 0 -1 3770
box -8 -3 16 105
use FILL  FILL_163
timestamp 1682952543
transform 1 0 848 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_27
timestamp 1682952543
transform -1 0 896 0 -1 3770
box -8 -3 46 105
use FILL  FILL_164
timestamp 1682952543
transform 1 0 896 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_51
timestamp 1682952543
transform 1 0 904 0 -1 3770
box -9 -3 26 105
use FILL  FILL_165
timestamp 1682952543
transform 1 0 920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_166
timestamp 1682952543
transform 1 0 928 0 -1 3770
box -8 -3 16 105
use FILL  FILL_167
timestamp 1682952543
transform 1 0 936 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1682952543
transform 1 0 944 0 -1 3770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1682952543
transform 1 0 968 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_52
timestamp 1682952543
transform -1 0 1080 0 -1 3770
box -9 -3 26 105
use AOI22X1  AOI22X1_28
timestamp 1682952543
transform 1 0 1080 0 -1 3770
box -8 -3 46 105
use FILL  FILL_168
timestamp 1682952543
transform 1 0 1120 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_34
timestamp 1682952543
transform -1 0 1168 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_35
timestamp 1682952543
transform -1 0 1208 0 -1 3770
box -8 -3 46 105
use FILL  FILL_169
timestamp 1682952543
transform 1 0 1208 0 -1 3770
box -8 -3 16 105
use FILL  FILL_170
timestamp 1682952543
transform 1 0 1216 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_53
timestamp 1682952543
transform 1 0 1224 0 -1 3770
box -9 -3 26 105
use FILL  FILL_171
timestamp 1682952543
transform 1 0 1240 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_54
timestamp 1682952543
transform 1 0 1248 0 -1 3770
box -9 -3 26 105
use AOI22X1  AOI22X1_29
timestamp 1682952543
transform 1 0 1264 0 -1 3770
box -8 -3 46 105
use FILL  FILL_172
timestamp 1682952543
transform 1 0 1304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_173
timestamp 1682952543
transform 1 0 1312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_174
timestamp 1682952543
transform 1 0 1320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_175
timestamp 1682952543
transform 1 0 1328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_176
timestamp 1682952543
transform 1 0 1336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_177
timestamp 1682952543
transform 1 0 1344 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_30
timestamp 1682952543
transform 1 0 1352 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_55
timestamp 1682952543
transform 1 0 1392 0 -1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_63
timestamp 1682952543
transform -1 0 1504 0 -1 3770
box -8 -3 104 105
use BUFX2  BUFX2_0
timestamp 1682952543
transform 1 0 1504 0 -1 3770
box -5 -3 28 105
use FILL  FILL_199
timestamp 1682952543
transform 1 0 1528 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1682952543
transform -1 0 1632 0 -1 3770
box -8 -3 104 105
use FILL  FILL_200
timestamp 1682952543
transform 1 0 1632 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1682952543
transform -1 0 1736 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1682952543
transform -1 0 1832 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_60
timestamp 1682952543
transform 1 0 1832 0 -1 3770
box -9 -3 26 105
use FILL  FILL_201
timestamp 1682952543
transform 1 0 1848 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1682952543
transform -1 0 1952 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1682952543
transform -1 0 2048 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_69
timestamp 1682952543
transform 1 0 2048 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_61
timestamp 1682952543
transform 1 0 2144 0 -1 3770
box -9 -3 26 105
use FILL  FILL_202
timestamp 1682952543
transform 1 0 2160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_203
timestamp 1682952543
transform 1 0 2168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_204
timestamp 1682952543
transform 1 0 2176 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_38
timestamp 1682952543
transform 1 0 2184 0 -1 3770
box -8 -3 46 105
use BUFX2  BUFX2_1
timestamp 1682952543
transform 1 0 2224 0 -1 3770
box -5 -3 28 105
use FILL  FILL_205
timestamp 1682952543
transform 1 0 2248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_206
timestamp 1682952543
transform 1 0 2256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_208
timestamp 1682952543
transform 1 0 2264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_211
timestamp 1682952543
transform 1 0 2272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_212
timestamp 1682952543
transform 1 0 2280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_213
timestamp 1682952543
transform 1 0 2288 0 -1 3770
box -8 -3 16 105
use BUFX2  BUFX2_2
timestamp 1682952543
transform 1 0 2296 0 -1 3770
box -5 -3 28 105
use FILL  FILL_214
timestamp 1682952543
transform 1 0 2320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_216
timestamp 1682952543
transform 1 0 2328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_218
timestamp 1682952543
transform 1 0 2336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_219
timestamp 1682952543
transform 1 0 2344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_220
timestamp 1682952543
transform 1 0 2352 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_41
timestamp 1682952543
transform 1 0 2360 0 -1 3770
box -8 -3 46 105
use FILL  FILL_227
timestamp 1682952543
transform 1 0 2400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_228
timestamp 1682952543
transform 1 0 2408 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_52
timestamp 1682952543
transform 1 0 2416 0 -1 3770
box -8 -3 46 105
use FILL  FILL_229
timestamp 1682952543
transform 1 0 2456 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_53
timestamp 1682952543
transform 1 0 2464 0 -1 3770
box -8 -3 46 105
use FILL  FILL_230
timestamp 1682952543
transform 1 0 2504 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_54
timestamp 1682952543
transform 1 0 2512 0 -1 3770
box -8 -3 46 105
use FILL  FILL_231
timestamp 1682952543
transform 1 0 2552 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_55
timestamp 1682952543
transform 1 0 2560 0 -1 3770
box -8 -3 46 105
use FILL  FILL_232
timestamp 1682952543
transform 1 0 2600 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_56
timestamp 1682952543
transform 1 0 2608 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_57
timestamp 1682952543
transform 1 0 2648 0 -1 3770
box -8 -3 46 105
use FILL  FILL_233
timestamp 1682952543
transform 1 0 2688 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_70
timestamp 1682952543
transform -1 0 2712 0 -1 3770
box -9 -3 26 105
use FILL  FILL_234
timestamp 1682952543
transform 1 0 2712 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_58
timestamp 1682952543
transform -1 0 2760 0 -1 3770
box -8 -3 46 105
use FILL  FILL_235
timestamp 1682952543
transform 1 0 2760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_236
timestamp 1682952543
transform 1 0 2768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_237
timestamp 1682952543
transform 1 0 2776 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_59
timestamp 1682952543
transform 1 0 2784 0 -1 3770
box -8 -3 46 105
use FILL  FILL_238
timestamp 1682952543
transform 1 0 2824 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_71
timestamp 1682952543
transform -1 0 2848 0 -1 3770
box -9 -3 26 105
use M3_M2  M3_M2_909
timestamp 1682952543
transform 1 0 2876 0 1 3675
box -3 -3 3 3
use OAI22X1  OAI22X1_60
timestamp 1682952543
transform 1 0 2848 0 -1 3770
box -8 -3 46 105
use M3_M2  M3_M2_910
timestamp 1682952543
transform 1 0 2932 0 1 3675
box -3 -3 3 3
use OAI22X1  OAI22X1_61
timestamp 1682952543
transform 1 0 2888 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_62
timestamp 1682952543
transform 1 0 2928 0 -1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1682952543
transform 1 0 2968 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_72
timestamp 1682952543
transform -1 0 3080 0 -1 3770
box -9 -3 26 105
use FILL  FILL_239
timestamp 1682952543
transform 1 0 3080 0 -1 3770
box -8 -3 16 105
use FILL  FILL_240
timestamp 1682952543
transform 1 0 3088 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_63
timestamp 1682952543
transform 1 0 3096 0 -1 3770
box -8 -3 46 105
use FILL  FILL_241
timestamp 1682952543
transform 1 0 3136 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_911
timestamp 1682952543
transform 1 0 3156 0 1 3675
box -3 -3 3 3
use FILL  FILL_242
timestamp 1682952543
transform 1 0 3144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_243
timestamp 1682952543
transform 1 0 3152 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_73
timestamp 1682952543
transform -1 0 3176 0 -1 3770
box -9 -3 26 105
use FILL  FILL_244
timestamp 1682952543
transform 1 0 3176 0 -1 3770
box -8 -3 16 105
use FILL  FILL_245
timestamp 1682952543
transform 1 0 3184 0 -1 3770
box -8 -3 16 105
use FILL  FILL_246
timestamp 1682952543
transform 1 0 3192 0 -1 3770
box -8 -3 16 105
use FILL  FILL_247
timestamp 1682952543
transform 1 0 3200 0 -1 3770
box -8 -3 16 105
use FILL  FILL_248
timestamp 1682952543
transform 1 0 3208 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_64
timestamp 1682952543
transform 1 0 3216 0 -1 3770
box -8 -3 46 105
use FILL  FILL_249
timestamp 1682952543
transform 1 0 3256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_250
timestamp 1682952543
transform 1 0 3264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_251
timestamp 1682952543
transform 1 0 3272 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_74
timestamp 1682952543
transform -1 0 3296 0 -1 3770
box -9 -3 26 105
use FILL  FILL_252
timestamp 1682952543
transform 1 0 3296 0 -1 3770
box -8 -3 16 105
use FILL  FILL_253
timestamp 1682952543
transform 1 0 3304 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_65
timestamp 1682952543
transform 1 0 3312 0 -1 3770
box -8 -3 46 105
use FILL  FILL_254
timestamp 1682952543
transform 1 0 3352 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_66
timestamp 1682952543
transform -1 0 3400 0 -1 3770
box -8 -3 46 105
use FILL  FILL_255
timestamp 1682952543
transform 1 0 3400 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1682952543
transform 1 0 3408 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_75
timestamp 1682952543
transform 1 0 3504 0 -1 3770
box -9 -3 26 105
use M3_M2  M3_M2_912
timestamp 1682952543
transform 1 0 3564 0 1 3675
box -3 -3 3 3
use OAI22X1  OAI22X1_67
timestamp 1682952543
transform -1 0 3560 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_76
timestamp 1682952543
transform 1 0 3560 0 -1 3770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_80
timestamp 1682952543
transform 1 0 3576 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_77
timestamp 1682952543
transform 1 0 3672 0 -1 3770
box -9 -3 26 105
use OAI22X1  OAI22X1_68
timestamp 1682952543
transform 1 0 3688 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_70
timestamp 1682952543
transform 1 0 3728 0 -1 3770
box -8 -3 46 105
use OAI21X1  OAI21X1_0
timestamp 1682952543
transform 1 0 3768 0 -1 3770
box -8 -3 34 105
use OAI22X1  OAI22X1_75
timestamp 1682952543
transform 1 0 3800 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_76
timestamp 1682952543
transform 1 0 3840 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_77
timestamp 1682952543
transform 1 0 3880 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_78
timestamp 1682952543
transform 1 0 3920 0 -1 3770
box -8 -3 46 105
use OAI22X1  OAI22X1_79
timestamp 1682952543
transform 1 0 3960 0 -1 3770
box -8 -3 46 105
use M3_M2  M3_M2_913
timestamp 1682952543
transform 1 0 4012 0 1 3675
box -3 -3 3 3
use OAI22X1  OAI22X1_80
timestamp 1682952543
transform 1 0 4000 0 -1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1682952543
transform 1 0 4040 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_80
timestamp 1682952543
transform -1 0 4152 0 -1 3770
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_9
timestamp 1682952543
transform 1 0 4201 0 1 3670
box -10 -3 10 3
use M2_M1  M2_M1_1007
timestamp 1682952543
transform 1 0 132 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1682952543
transform 1 0 164 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1009
timestamp 1682952543
transform 1 0 172 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1682952543
transform 1 0 84 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1080
timestamp 1682952543
transform 1 0 132 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1081
timestamp 1682952543
transform 1 0 172 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1682952543
transform 1 0 244 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1682952543
transform 1 0 284 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1010
timestamp 1682952543
transform 1 0 244 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1041
timestamp 1682952543
transform 1 0 268 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1682952543
transform 1 0 276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1682952543
transform 1 0 284 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1682952543
transform 1 0 292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1682952543
transform 1 0 180 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1682952543
transform 1 0 196 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1101
timestamp 1682952543
transform 1 0 84 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1102
timestamp 1682952543
transform 1 0 148 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1082
timestamp 1682952543
transform 1 0 292 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1103
timestamp 1682952543
transform 1 0 276 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1042
timestamp 1682952543
transform 1 0 316 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1014
timestamp 1682952543
transform 1 0 324 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1043
timestamp 1682952543
transform 1 0 332 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1145
timestamp 1682952543
transform 1 0 308 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1682952543
transform 1 0 316 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1682952543
transform 1 0 332 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1682952543
transform 1 0 340 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1104
timestamp 1682952543
transform 1 0 332 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_1015
timestamp 1682952543
transform 1 0 356 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1682952543
transform 1 0 388 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1044
timestamp 1682952543
transform 1 0 396 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_914
timestamp 1682952543
transform 1 0 412 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_1017
timestamp 1682952543
transform 1 0 412 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1682952543
transform 1 0 380 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1682952543
transform 1 0 396 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1151
timestamp 1682952543
transform 1 0 404 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1105
timestamp 1682952543
transform 1 0 380 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1106
timestamp 1682952543
transform 1 0 404 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1001
timestamp 1682952543
transform 1 0 444 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1018
timestamp 1682952543
transform 1 0 444 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1682952543
transform 1 0 460 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1152
timestamp 1682952543
transform 1 0 452 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_931
timestamp 1682952543
transform 1 0 484 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_1020
timestamp 1682952543
transform 1 0 484 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1682952543
transform 1 0 484 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1107
timestamp 1682952543
transform 1 0 476 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1153
timestamp 1682952543
transform 1 0 468 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_915
timestamp 1682952543
transform 1 0 532 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1682952543
transform 1 0 532 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1682952543
transform 1 0 500 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1682952543
transform 1 0 580 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1021
timestamp 1682952543
transform 1 0 524 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1022
timestamp 1682952543
transform 1 0 580 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1682952543
transform 1 0 500 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1108
timestamp 1682952543
transform 1 0 500 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1682952543
transform 1 0 532 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1682952543
transform 1 0 604 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1682952543
transform 1 0 604 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1682952543
transform 1 0 596 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_948
timestamp 1682952543
transform 1 0 636 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_1024
timestamp 1682952543
transform 1 0 636 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1045
timestamp 1682952543
transform 1 0 644 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1025
timestamp 1682952543
transform 1 0 652 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1682952543
transform 1 0 660 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1083
timestamp 1682952543
transform 1 0 620 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1156
timestamp 1682952543
transform 1 0 628 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1682952543
transform 1 0 644 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1158
timestamp 1682952543
transform 1 0 652 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_932
timestamp 1682952543
transform 1 0 684 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1682952543
transform 1 0 676 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1682952543
transform 1 0 724 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1682952543
transform 1 0 708 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1027
timestamp 1682952543
transform 1 0 684 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1682952543
transform 1 0 700 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1046
timestamp 1682952543
transform 1 0 716 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_949
timestamp 1682952543
transform 1 0 780 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_950
timestamp 1682952543
transform 1 0 812 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_951
timestamp 1682952543
transform 1 0 828 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1682952543
transform 1 0 796 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1682952543
transform 1 0 788 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1682952543
transform 1 0 804 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1682952543
transform 1 0 844 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1029
timestamp 1682952543
transform 1 0 724 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1682952543
transform 1 0 740 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1682952543
transform 1 0 756 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1682952543
transform 1 0 772 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1033
timestamp 1682952543
transform 1 0 788 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1682952543
transform 1 0 804 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1682952543
transform 1 0 812 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1682952543
transform 1 0 844 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1682952543
transform 1 0 676 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1160
timestamp 1682952543
transform 1 0 692 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1084
timestamp 1682952543
transform 1 0 700 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1161
timestamp 1682952543
transform 1 0 708 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1682952543
transform 1 0 716 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1682952543
transform 1 0 732 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1154
timestamp 1682952543
transform 1 0 692 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1085
timestamp 1682952543
transform 1 0 740 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1164
timestamp 1682952543
transform 1 0 764 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1165
timestamp 1682952543
transform 1 0 780 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1682952543
transform 1 0 788 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1110
timestamp 1682952543
transform 1 0 764 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_1167
timestamp 1682952543
transform 1 0 892 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1111
timestamp 1682952543
transform 1 0 812 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_1168
timestamp 1682952543
transform 1 0 916 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1284
timestamp 1682952543
transform 1 0 908 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_1155
timestamp 1682952543
transform 1 0 908 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_1285
timestamp 1682952543
transform 1 0 924 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_1156
timestamp 1682952543
transform 1 0 924 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1682952543
transform 1 0 948 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1037
timestamp 1682952543
transform 1 0 948 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1008
timestamp 1682952543
transform 1 0 1028 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1009
timestamp 1682952543
transform 1 0 1068 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1038
timestamp 1682952543
transform 1 0 964 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1682952543
transform 1 0 1028 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1682952543
transform 1 0 1060 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1682952543
transform 1 0 1068 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1086
timestamp 1682952543
transform 1 0 964 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1169
timestamp 1682952543
transform 1 0 980 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1286
timestamp 1682952543
transform 1 0 964 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_1112
timestamp 1682952543
transform 1 0 1060 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_952
timestamp 1682952543
transform 1 0 1092 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1010
timestamp 1682952543
transform 1 0 1092 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1042
timestamp 1682952543
transform 1 0 1092 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1047
timestamp 1682952543
transform 1 0 1116 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1682952543
transform 1 0 1148 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1043
timestamp 1682952543
transform 1 0 1124 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1682952543
transform 1 0 1140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1170
timestamp 1682952543
transform 1 0 1108 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1171
timestamp 1682952543
transform 1 0 1116 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1682952543
transform 1 0 1132 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1113
timestamp 1682952543
transform 1 0 1132 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1682952543
transform 1 0 1156 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1045
timestamp 1682952543
transform 1 0 1180 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1682952543
transform 1 0 1196 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1682952543
transform 1 0 1188 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1114
timestamp 1682952543
transform 1 0 1180 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1115
timestamp 1682952543
transform 1 0 1196 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1682952543
transform 1 0 1220 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_916
timestamp 1682952543
transform 1 0 1276 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1682952543
transform 1 0 1308 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1011
timestamp 1682952543
transform 1 0 1324 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1047
timestamp 1682952543
transform 1 0 1228 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1682952543
transform 1 0 1260 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1682952543
transform 1 0 1324 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1174
timestamp 1682952543
transform 1 0 1220 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1682952543
transform 1 0 1308 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1682952543
transform 1 0 1324 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_953
timestamp 1682952543
transform 1 0 1348 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_1050
timestamp 1682952543
transform 1 0 1340 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1012
timestamp 1682952543
transform 1 0 1380 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1051
timestamp 1682952543
transform 1 0 1364 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1050
timestamp 1682952543
transform 1 0 1372 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1052
timestamp 1682952543
transform 1 0 1380 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1177
timestamp 1682952543
transform 1 0 1348 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1682952543
transform 1 0 1372 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1682952543
transform 1 0 1380 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_978
timestamp 1682952543
transform 1 0 1484 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1682952543
transform 1 0 1396 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1682952543
transform 1 0 1436 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1053
timestamp 1682952543
transform 1 0 1396 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1682952543
transform 1 0 1404 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1051
timestamp 1682952543
transform 1 0 1412 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1055
timestamp 1682952543
transform 1 0 1436 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1682952543
transform 1 0 1500 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1180
timestamp 1682952543
transform 1 0 1484 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_979
timestamp 1682952543
transform 1 0 1556 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1682952543
transform 1 0 1564 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1057
timestamp 1682952543
transform 1 0 1532 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1052
timestamp 1682952543
transform 1 0 1540 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1058
timestamp 1682952543
transform 1 0 1548 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_917
timestamp 1682952543
transform 1 0 1604 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_1059
timestamp 1682952543
transform 1 0 1572 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1053
timestamp 1682952543
transform 1 0 1580 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1060
timestamp 1682952543
transform 1 0 1588 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1054
timestamp 1682952543
transform 1 0 1596 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1061
timestamp 1682952543
transform 1 0 1604 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1062
timestamp 1682952543
transform 1 0 1620 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1055
timestamp 1682952543
transform 1 0 1628 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1063
timestamp 1682952543
transform 1 0 1644 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1682952543
transform 1 0 1516 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1182
timestamp 1682952543
transform 1 0 1524 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1682952543
transform 1 0 1540 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1682952543
transform 1 0 1556 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1682952543
transform 1 0 1564 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1682952543
transform 1 0 1580 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1682952543
transform 1 0 1596 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1682952543
transform 1 0 1612 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1682952543
transform 1 0 1628 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1682952543
transform 1 0 1636 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1116
timestamp 1682952543
transform 1 0 1540 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1682952543
transform 1 0 1580 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_1064
timestamp 1682952543
transform 1 0 1660 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1682952543
transform 1 0 1660 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_918
timestamp 1682952543
transform 1 0 1700 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1682952543
transform 1 0 1780 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1682952543
transform 1 0 1748 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_955
timestamp 1682952543
transform 1 0 1764 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1016
timestamp 1682952543
transform 1 0 1684 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1682952543
transform 1 0 1780 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1065
timestamp 1682952543
transform 1 0 1676 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1682952543
transform 1 0 1684 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1682952543
transform 1 0 1740 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1087
timestamp 1682952543
transform 1 0 1740 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1192
timestamp 1682952543
transform 1 0 1764 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_919
timestamp 1682952543
transform 1 0 1812 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_935
timestamp 1682952543
transform 1 0 1796 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1682952543
transform 1 0 1820 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1682952543
transform 1 0 1804 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1068
timestamp 1682952543
transform 1 0 1788 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1682952543
transform 1 0 1804 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1682952543
transform 1 0 1820 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1682952543
transform 1 0 1828 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1193
timestamp 1682952543
transform 1 0 1780 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1682952543
transform 1 0 1812 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1117
timestamp 1682952543
transform 1 0 1812 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1088
timestamp 1682952543
transform 1 0 1828 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1019
timestamp 1682952543
transform 1 0 1844 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1072
timestamp 1682952543
transform 1 0 1852 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1682952543
transform 1 0 1844 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1056
timestamp 1682952543
transform 1 0 1860 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_957
timestamp 1682952543
transform 1 0 1884 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_958
timestamp 1682952543
transform 1 0 1900 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1682952543
transform 1 0 1900 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1682952543
transform 1 0 1892 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1073
timestamp 1682952543
transform 1 0 1876 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1057
timestamp 1682952543
transform 1 0 1884 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1074
timestamp 1682952543
transform 1 0 1892 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1682952543
transform 1 0 1860 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1682952543
transform 1 0 1868 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1118
timestamp 1682952543
transform 1 0 1860 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1089
timestamp 1682952543
transform 1 0 1876 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1682952543
transform 1 0 1924 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_1075
timestamp 1682952543
transform 1 0 1916 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1682952543
transform 1 0 1900 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1682952543
transform 1 0 1908 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1158
timestamp 1682952543
transform 1 0 1876 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1682952543
transform 1 0 1932 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1682952543
transform 1 0 1956 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1682952543
transform 1 0 1988 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_983
timestamp 1682952543
transform 1 0 2004 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1682952543
transform 1 0 1948 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1159
timestamp 1682952543
transform 1 0 1940 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1023
timestamp 1682952543
transform 1 0 1988 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1076
timestamp 1682952543
transform 1 0 1948 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1682952543
transform 1 0 1956 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1682952543
transform 1 0 1988 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1058
timestamp 1682952543
transform 1 0 2036 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1682952543
transform 1 0 2036 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1119
timestamp 1682952543
transform 1 0 1964 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1682952543
transform 1 0 2148 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_1079
timestamp 1682952543
transform 1 0 2116 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1682952543
transform 1 0 2068 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1120
timestamp 1682952543
transform 1 0 2116 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1090
timestamp 1682952543
transform 1 0 2156 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_984
timestamp 1682952543
transform 1 0 2180 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1682952543
transform 1 0 2228 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1682952543
transform 1 0 2180 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1682952543
transform 1 0 2212 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1059
timestamp 1682952543
transform 1 0 2172 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1080
timestamp 1682952543
transform 1 0 2196 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1060
timestamp 1682952543
transform 1 0 2204 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1081
timestamp 1682952543
transform 1 0 2212 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1682952543
transform 1 0 2228 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1202
timestamp 1682952543
transform 1 0 2188 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1682952543
transform 1 0 2204 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1682952543
transform 1 0 2220 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1205
timestamp 1682952543
transform 1 0 2228 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1121
timestamp 1682952543
transform 1 0 2204 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1160
timestamp 1682952543
transform 1 0 2188 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_985
timestamp 1682952543
transform 1 0 2236 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1083
timestamp 1682952543
transform 1 0 2284 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1061
timestamp 1682952543
transform 1 0 2324 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1682952543
transform 1 0 2380 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_960
timestamp 1682952543
transform 1 0 2412 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_1084
timestamp 1682952543
transform 1 0 2348 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1682952543
transform 1 0 2364 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1682952543
transform 1 0 2380 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1062
timestamp 1682952543
transform 1 0 2388 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1087
timestamp 1682952543
transform 1 0 2396 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1206
timestamp 1682952543
transform 1 0 2252 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1091
timestamp 1682952543
transform 1 0 2340 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1207
timestamp 1682952543
transform 1 0 2356 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1092
timestamp 1682952543
transform 1 0 2364 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1208
timestamp 1682952543
transform 1 0 2372 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1209
timestamp 1682952543
transform 1 0 2388 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1210
timestamp 1682952543
transform 1 0 2396 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1122
timestamp 1682952543
transform 1 0 2252 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1682952543
transform 1 0 2228 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1162
timestamp 1682952543
transform 1 0 2268 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1682952543
transform 1 0 2332 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_994
timestamp 1682952543
transform 1 0 2420 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1123
timestamp 1682952543
transform 1 0 2372 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1124
timestamp 1682952543
transform 1 0 2396 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1682952543
transform 1 0 2388 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_1088
timestamp 1682952543
transform 1 0 2444 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1093
timestamp 1682952543
transform 1 0 2444 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1682952543
transform 1 0 2476 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1682952543
transform 1 0 2484 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1089
timestamp 1682952543
transform 1 0 2484 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1682952543
transform 1 0 2452 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1682952543
transform 1 0 2460 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1682952543
transform 1 0 2476 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1165
timestamp 1682952543
transform 1 0 2444 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1094
timestamp 1682952543
transform 1 0 2484 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1682952543
transform 1 0 2532 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_961
timestamp 1682952543
transform 1 0 2524 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1063
timestamp 1682952543
transform 1 0 2508 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_988
timestamp 1682952543
transform 1 0 2532 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_995
timestamp 1682952543
transform 1 0 2532 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1682952543
transform 1 0 2516 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1682952543
transform 1 0 2532 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1214
timestamp 1682952543
transform 1 0 2492 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1215
timestamp 1682952543
transform 1 0 2500 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1125
timestamp 1682952543
transform 1 0 2476 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1126
timestamp 1682952543
transform 1 0 2500 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1166
timestamp 1682952543
transform 1 0 2532 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_989
timestamp 1682952543
transform 1 0 2548 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1027
timestamp 1682952543
transform 1 0 2580 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1064
timestamp 1682952543
transform 1 0 2572 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1092
timestamp 1682952543
transform 1 0 2580 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1216
timestamp 1682952543
transform 1 0 2548 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1682952543
transform 1 0 2556 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1218
timestamp 1682952543
transform 1 0 2572 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1219
timestamp 1682952543
transform 1 0 2588 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1220
timestamp 1682952543
transform 1 0 2596 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1127
timestamp 1682952543
transform 1 0 2572 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1682952543
transform 1 0 2604 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1682952543
transform 1 0 2596 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1682952543
transform 1 0 2644 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_996
timestamp 1682952543
transform 1 0 2644 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1682952543
transform 1 0 2628 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1682952543
transform 1 0 2644 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1167
timestamp 1682952543
transform 1 0 2644 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1682952543
transform 1 0 2660 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_1221
timestamp 1682952543
transform 1 0 2660 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1682952543
transform 1 0 2652 0 1 3595
box -2 -2 2 2
use M3_M2  M3_M2_1129
timestamp 1682952543
transform 1 0 2660 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1682952543
transform 1 0 2660 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1029
timestamp 1682952543
transform 1 0 2700 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1065
timestamp 1682952543
transform 1 0 2692 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1095
timestamp 1682952543
transform 1 0 2700 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1682952543
transform 1 0 2732 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1682952543
transform 1 0 2724 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1682952543
transform 1 0 2692 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1223
timestamp 1682952543
transform 1 0 2708 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1224
timestamp 1682952543
transform 1 0 2716 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1130
timestamp 1682952543
transform 1 0 2692 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1169
timestamp 1682952543
transform 1 0 2684 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1066
timestamp 1682952543
transform 1 0 2732 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1097
timestamp 1682952543
transform 1 0 2740 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1682952543
transform 1 0 2732 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1131
timestamp 1682952543
transform 1 0 2732 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1682952543
transform 1 0 2740 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_938
timestamp 1682952543
transform 1 0 2772 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_939
timestamp 1682952543
transform 1 0 2796 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1682952543
transform 1 0 2764 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1226
timestamp 1682952543
transform 1 0 2764 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_963
timestamp 1682952543
transform 1 0 2780 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_998
timestamp 1682952543
transform 1 0 2780 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1068
timestamp 1682952543
transform 1 0 2780 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1227
timestamp 1682952543
transform 1 0 2780 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1132
timestamp 1682952543
transform 1 0 2772 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1682952543
transform 1 0 2812 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_990
timestamp 1682952543
transform 1 0 2812 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1098
timestamp 1682952543
transform 1 0 2804 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1030
timestamp 1682952543
transform 1 0 2820 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1228
timestamp 1682952543
transform 1 0 2804 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1229
timestamp 1682952543
transform 1 0 2812 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1682952543
transform 1 0 2852 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1069
timestamp 1682952543
transform 1 0 2852 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1099
timestamp 1682952543
transform 1 0 2860 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1682952543
transform 1 0 2868 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1171
timestamp 1682952543
transform 1 0 2844 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_1230
timestamp 1682952543
transform 1 0 2868 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1000
timestamp 1682952543
transform 1 0 2892 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1682952543
transform 1 0 2900 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1682952543
transform 1 0 2916 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_991
timestamp 1682952543
transform 1 0 2948 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1103
timestamp 1682952543
transform 1 0 2932 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1682952543
transform 1 0 2948 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_923
timestamp 1682952543
transform 1 0 2972 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_940
timestamp 1682952543
transform 1 0 2988 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1031
timestamp 1682952543
transform 1 0 2980 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1032
timestamp 1682952543
transform 1 0 2996 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1105
timestamp 1682952543
transform 1 0 2972 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1682952543
transform 1 0 2988 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1682952543
transform 1 0 2996 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_964
timestamp 1682952543
transform 1 0 3036 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1682952543
transform 1 0 3052 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_1231
timestamp 1682952543
transform 1 0 2916 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1232
timestamp 1682952543
transform 1 0 2924 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1682952543
transform 1 0 2940 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1682952543
transform 1 0 2956 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1235
timestamp 1682952543
transform 1 0 2964 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1236
timestamp 1682952543
transform 1 0 2980 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1237
timestamp 1682952543
transform 1 0 2996 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1682952543
transform 1 0 3004 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1133
timestamp 1682952543
transform 1 0 2924 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1134
timestamp 1682952543
transform 1 0 2964 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1095
timestamp 1682952543
transform 1 0 3012 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1239
timestamp 1682952543
transform 1 0 3028 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1001
timestamp 1682952543
transform 1 0 3036 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1033
timestamp 1682952543
transform 1 0 3060 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1108
timestamp 1682952543
transform 1 0 3060 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1682952543
transform 1 0 3076 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1110
timestamp 1682952543
transform 1 0 3092 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_924
timestamp 1682952543
transform 1 0 3116 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_941
timestamp 1682952543
transform 1 0 3132 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_966
timestamp 1682952543
transform 1 0 3124 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_967
timestamp 1682952543
transform 1 0 3188 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1682952543
transform 1 0 3172 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1034
timestamp 1682952543
transform 1 0 3156 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1682952543
transform 1 0 3188 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1111
timestamp 1682952543
transform 1 0 3116 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1070
timestamp 1682952543
transform 1 0 3124 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1112
timestamp 1682952543
transform 1 0 3132 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1071
timestamp 1682952543
transform 1 0 3140 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1113
timestamp 1682952543
transform 1 0 3156 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1072
timestamp 1682952543
transform 1 0 3164 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1114
timestamp 1682952543
transform 1 0 3172 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1073
timestamp 1682952543
transform 1 0 3180 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1115
timestamp 1682952543
transform 1 0 3188 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1240
timestamp 1682952543
transform 1 0 3036 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1241
timestamp 1682952543
transform 1 0 3060 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1682952543
transform 1 0 3068 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1243
timestamp 1682952543
transform 1 0 3084 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1244
timestamp 1682952543
transform 1 0 3100 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1245
timestamp 1682952543
transform 1 0 3108 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1246
timestamp 1682952543
transform 1 0 3124 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1247
timestamp 1682952543
transform 1 0 3140 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1682952543
transform 1 0 3148 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1249
timestamp 1682952543
transform 1 0 3164 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1682952543
transform 1 0 3180 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1682952543
transform 1 0 3188 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1135
timestamp 1682952543
transform 1 0 3060 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1682952543
transform 1 0 3084 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1137
timestamp 1682952543
transform 1 0 3108 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1682952543
transform 1 0 3148 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1172
timestamp 1682952543
transform 1 0 3148 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_993
timestamp 1682952543
transform 1 0 3212 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1116
timestamp 1682952543
transform 1 0 3212 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1682952543
transform 1 0 3204 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_968
timestamp 1682952543
transform 1 0 3236 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1682952543
transform 1 0 3252 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1682952543
transform 1 0 3276 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_942
timestamp 1682952543
transform 1 0 3292 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1036
timestamp 1682952543
transform 1 0 3260 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1117
timestamp 1682952543
transform 1 0 3236 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1682952543
transform 1 0 3252 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1074
timestamp 1682952543
transform 1 0 3260 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1119
timestamp 1682952543
transform 1 0 3276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1682952543
transform 1 0 3292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1253
timestamp 1682952543
transform 1 0 3228 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1096
timestamp 1682952543
transform 1 0 3236 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1075
timestamp 1682952543
transform 1 0 3300 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1254
timestamp 1682952543
transform 1 0 3244 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1255
timestamp 1682952543
transform 1 0 3260 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1682952543
transform 1 0 3268 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1257
timestamp 1682952543
transform 1 0 3284 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1258
timestamp 1682952543
transform 1 0 3300 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1139
timestamp 1682952543
transform 1 0 3228 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1140
timestamp 1682952543
transform 1 0 3268 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1682952543
transform 1 0 3372 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_943
timestamp 1682952543
transform 1 0 3332 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_944
timestamp 1682952543
transform 1 0 3364 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1682952543
transform 1 0 3340 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_995
timestamp 1682952543
transform 1 0 3316 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1682952543
transform 1 0 3348 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1121
timestamp 1682952543
transform 1 0 3372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1259
timestamp 1682952543
transform 1 0 3324 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1141
timestamp 1682952543
transform 1 0 3372 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_945
timestamp 1682952543
transform 1 0 3420 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1682952543
transform 1 0 3444 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1682952543
transform 1 0 3452 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1122
timestamp 1682952543
transform 1 0 3420 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1076
timestamp 1682952543
transform 1 0 3428 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1123
timestamp 1682952543
transform 1 0 3452 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1682952543
transform 1 0 3428 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1682952543
transform 1 0 3444 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1097
timestamp 1682952543
transform 1 0 3452 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1682952543
transform 1 0 3564 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1682952543
transform 1 0 3476 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1039
timestamp 1682952543
transform 1 0 3500 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1124
timestamp 1682952543
transform 1 0 3500 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1125
timestamp 1682952543
transform 1 0 3556 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1682952543
transform 1 0 3564 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1682952543
transform 1 0 3460 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1263
timestamp 1682952543
transform 1 0 3476 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1142
timestamp 1682952543
transform 1 0 3444 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1098
timestamp 1682952543
transform 1 0 3500 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1264
timestamp 1682952543
transform 1 0 3564 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1143
timestamp 1682952543
transform 1 0 3476 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1682952543
transform 1 0 3468 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1682952543
transform 1 0 3612 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_996
timestamp 1682952543
transform 1 0 3652 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1127
timestamp 1682952543
transform 1 0 3636 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1682952543
transform 1 0 3588 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1144
timestamp 1682952543
transform 1 0 3588 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1145
timestamp 1682952543
transform 1 0 3636 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1682952543
transform 1 0 3660 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1077
timestamp 1682952543
transform 1 0 3700 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1128
timestamp 1682952543
transform 1 0 3708 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1682952543
transform 1 0 3724 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1682952543
transform 1 0 3700 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1682952543
transform 1 0 3716 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1268
timestamp 1682952543
transform 1 0 3732 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1269
timestamp 1682952543
transform 1 0 3740 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1146
timestamp 1682952543
transform 1 0 3716 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1682952543
transform 1 0 3732 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_1130
timestamp 1682952543
transform 1 0 3756 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1682952543
transform 1 0 3780 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1270
timestamp 1682952543
transform 1 0 3772 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1271
timestamp 1682952543
transform 1 0 3788 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1147
timestamp 1682952543
transform 1 0 3780 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1148
timestamp 1682952543
transform 1 0 3804 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1176
timestamp 1682952543
transform 1 0 3796 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1682952543
transform 1 0 3828 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1682952543
transform 1 0 3820 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1682952543
transform 1 0 3828 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1002
timestamp 1682952543
transform 1 0 3852 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1099
timestamp 1682952543
transform 1 0 3860 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_1133
timestamp 1682952543
transform 1 0 3884 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1273
timestamp 1682952543
transform 1 0 3868 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1682952543
transform 1 0 3876 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1149
timestamp 1682952543
transform 1 0 3868 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_1275
timestamp 1682952543
transform 1 0 3892 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1150
timestamp 1682952543
transform 1 0 3892 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_1003
timestamp 1682952543
transform 1 0 3908 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_930
timestamp 1682952543
transform 1 0 3948 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1682952543
transform 1 0 3932 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1004
timestamp 1682952543
transform 1 0 3932 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1682952543
transform 1 0 3916 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_998
timestamp 1682952543
transform 1 0 3964 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_1005
timestamp 1682952543
transform 1 0 3964 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1682952543
transform 1 0 3948 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1100
timestamp 1682952543
transform 1 0 3932 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1078
timestamp 1682952543
transform 1 0 3964 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_1136
timestamp 1682952543
transform 1 0 3980 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1276
timestamp 1682952543
transform 1 0 3956 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1682952543
transform 1 0 3964 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1682952543
transform 1 0 4012 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1682952543
transform 1 0 4004 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1278
timestamp 1682952543
transform 1 0 3988 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1682952543
transform 1 0 3996 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1079
timestamp 1682952543
transform 1 0 4012 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1682952543
transform 1 0 4068 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1682952543
transform 1 0 4052 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_1138
timestamp 1682952543
transform 1 0 4028 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1682952543
transform 1 0 4044 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1682952543
transform 1 0 4092 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1682952543
transform 1 0 4148 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1682952543
transform 1 0 4012 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1682952543
transform 1 0 4036 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1682952543
transform 1 0 4052 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1682952543
transform 1 0 4068 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1151
timestamp 1682952543
transform 1 0 4036 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1682952543
transform 1 0 4012 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1152
timestamp 1682952543
transform 1 0 4092 0 1 3595
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_10
timestamp 1682952543
transform 1 0 48 0 1 3570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_83
timestamp 1682952543
transform 1 0 72 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_81
timestamp 1682952543
transform -1 0 184 0 1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1682952543
transform 1 0 184 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_82
timestamp 1682952543
transform -1 0 296 0 1 3570
box -9 -3 26 105
use FILL  FILL_268
timestamp 1682952543
transform 1 0 296 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_35
timestamp 1682952543
transform 1 0 304 0 1 3570
box -8 -3 46 105
use FILL  FILL_269
timestamp 1682952543
transform 1 0 344 0 1 3570
box -8 -3 16 105
use FILL  FILL_270
timestamp 1682952543
transform 1 0 352 0 1 3570
box -8 -3 16 105
use FILL  FILL_271
timestamp 1682952543
transform 1 0 360 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1178
timestamp 1682952543
transform 1 0 380 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1682952543
transform 1 0 412 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_36
timestamp 1682952543
transform -1 0 408 0 1 3570
box -8 -3 46 105
use FILL  FILL_272
timestamp 1682952543
transform 1 0 408 0 1 3570
box -8 -3 16 105
use FILL  FILL_273
timestamp 1682952543
transform 1 0 416 0 1 3570
box -8 -3 16 105
use FILL  FILL_275
timestamp 1682952543
transform 1 0 424 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1180
timestamp 1682952543
transform 1 0 452 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_82
timestamp 1682952543
transform -1 0 472 0 1 3570
box -8 -3 46 105
use FILL  FILL_276
timestamp 1682952543
transform 1 0 472 0 1 3570
box -8 -3 16 105
use FILL  FILL_279
timestamp 1682952543
transform 1 0 480 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1682952543
transform 1 0 488 0 1 3570
box -8 -3 104 105
use FILL  FILL_281
timestamp 1682952543
transform 1 0 584 0 1 3570
box -8 -3 16 105
use FILL  FILL_282
timestamp 1682952543
transform 1 0 592 0 1 3570
box -8 -3 16 105
use FILL  FILL_283
timestamp 1682952543
transform 1 0 600 0 1 3570
box -8 -3 16 105
use FILL  FILL_284
timestamp 1682952543
transform 1 0 608 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_39
timestamp 1682952543
transform 1 0 616 0 1 3570
box -8 -3 46 105
use INVX2  INVX2_86
timestamp 1682952543
transform 1 0 656 0 1 3570
box -9 -3 26 105
use OAI22X1  OAI22X1_84
timestamp 1682952543
transform 1 0 672 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_85
timestamp 1682952543
transform 1 0 712 0 1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_41
timestamp 1682952543
transform -1 0 792 0 1 3570
box -8 -3 46 105
use INVX2  INVX2_87
timestamp 1682952543
transform 1 0 792 0 1 3570
box -9 -3 26 105
use M3_M2  M3_M2_1181
timestamp 1682952543
transform 1 0 876 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1682952543
transform 1 0 900 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_89
timestamp 1682952543
transform -1 0 904 0 1 3570
box -8 -3 104 105
use M3_M2  M3_M2_1183
timestamp 1682952543
transform 1 0 932 0 1 3575
box -3 -3 3 3
use NOR2X1  NOR2X1_7
timestamp 1682952543
transform 1 0 904 0 1 3570
box -8 -3 32 105
use FILL  FILL_287
timestamp 1682952543
transform 1 0 928 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1184
timestamp 1682952543
transform 1 0 948 0 1 3575
box -3 -3 3 3
use FILL  FILL_288
timestamp 1682952543
transform 1 0 936 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1682952543
transform 1 0 944 0 1 3570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1682952543
transform 1 0 968 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_88
timestamp 1682952543
transform -1 0 1080 0 1 3570
box -9 -3 26 105
use FILL  FILL_289
timestamp 1682952543
transform 1 0 1080 0 1 3570
box -8 -3 16 105
use FILL  FILL_290
timestamp 1682952543
transform 1 0 1088 0 1 3570
box -8 -3 16 105
use FILL  FILL_291
timestamp 1682952543
transform 1 0 1096 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_42
timestamp 1682952543
transform 1 0 1104 0 1 3570
box -8 -3 46 105
use FILL  FILL_292
timestamp 1682952543
transform 1 0 1144 0 1 3570
box -8 -3 16 105
use FILL  FILL_293
timestamp 1682952543
transform 1 0 1152 0 1 3570
box -8 -3 16 105
use FILL  FILL_294
timestamp 1682952543
transform 1 0 1160 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1185
timestamp 1682952543
transform 1 0 1188 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_86
timestamp 1682952543
transform -1 0 1208 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_1186
timestamp 1682952543
transform 1 0 1220 0 1 3575
box -3 -3 3 3
use FILL  FILL_295
timestamp 1682952543
transform 1 0 1208 0 1 3570
box -8 -3 16 105
use FILL  FILL_296
timestamp 1682952543
transform 1 0 1216 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1187
timestamp 1682952543
transform 1 0 1324 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_91
timestamp 1682952543
transform -1 0 1320 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_89
timestamp 1682952543
transform 1 0 1320 0 1 3570
box -9 -3 26 105
use FILL  FILL_297
timestamp 1682952543
transform 1 0 1336 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_43
timestamp 1682952543
transform 1 0 1344 0 1 3570
box -8 -3 46 105
use INVX2  INVX2_93
timestamp 1682952543
transform 1 0 1384 0 1 3570
box -9 -3 26 105
use M3_M2  M3_M2_1188
timestamp 1682952543
transform 1 0 1452 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1682952543
transform 1 0 1484 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_94
timestamp 1682952543
transform -1 0 1496 0 1 3570
box -8 -3 104 105
use BUFX2  BUFX2_5
timestamp 1682952543
transform 1 0 1496 0 1 3570
box -5 -3 28 105
use OAI22X1  OAI22X1_89
timestamp 1682952543
transform -1 0 1560 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_90
timestamp 1682952543
transform 1 0 1560 0 1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_47
timestamp 1682952543
transform 1 0 1600 0 1 3570
box -8 -3 46 105
use INVX2  INVX2_95
timestamp 1682952543
transform 1 0 1640 0 1 3570
box -9 -3 26 105
use INVX2  INVX2_96
timestamp 1682952543
transform 1 0 1656 0 1 3570
box -9 -3 26 105
use FILL  FILL_316
timestamp 1682952543
transform 1 0 1672 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1190
timestamp 1682952543
transform 1 0 1756 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_95
timestamp 1682952543
transform -1 0 1776 0 1 3570
box -8 -3 104 105
use M3_M2  M3_M2_1191
timestamp 1682952543
transform 1 0 1788 0 1 3575
box -3 -3 3 3
use FILL  FILL_317
timestamp 1682952543
transform 1 0 1776 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_48
timestamp 1682952543
transform -1 0 1824 0 1 3570
box -8 -3 46 105
use FILL  FILL_318
timestamp 1682952543
transform 1 0 1824 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_97
timestamp 1682952543
transform -1 0 1848 0 1 3570
box -9 -3 26 105
use FILL  FILL_319
timestamp 1682952543
transform 1 0 1848 0 1 3570
box -8 -3 16 105
use FILL  FILL_320
timestamp 1682952543
transform 1 0 1856 0 1 3570
box -8 -3 16 105
use FILL  FILL_321
timestamp 1682952543
transform 1 0 1864 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1192
timestamp 1682952543
transform 1 0 1916 0 1 3575
box -3 -3 3 3
use AOI22X1  AOI22X1_49
timestamp 1682952543
transform 1 0 1872 0 1 3570
box -8 -3 46 105
use FILL  FILL_322
timestamp 1682952543
transform 1 0 1912 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1193
timestamp 1682952543
transform 1 0 1940 0 1 3575
box -3 -3 3 3
use INVX2  INVX2_99
timestamp 1682952543
transform 1 0 1920 0 1 3570
box -9 -3 26 105
use FILL  FILL_330
timestamp 1682952543
transform 1 0 1936 0 1 3570
box -8 -3 16 105
use FILL  FILL_331
timestamp 1682952543
transform 1 0 1944 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1682952543
transform -1 0 2048 0 1 3570
box -8 -3 104 105
use FILL  FILL_332
timestamp 1682952543
transform 1 0 2048 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1194
timestamp 1682952543
transform 1 0 2068 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_1195
timestamp 1682952543
transform 1 0 2124 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_100
timestamp 1682952543
transform 1 0 2056 0 1 3570
box -8 -3 104 105
use FILL  FILL_333
timestamp 1682952543
transform 1 0 2152 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1196
timestamp 1682952543
transform 1 0 2196 0 1 3575
box -3 -3 3 3
use FILL  FILL_334
timestamp 1682952543
transform 1 0 2160 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_100
timestamp 1682952543
transform 1 0 2168 0 1 3570
box -9 -3 26 105
use OAI22X1  OAI22X1_93
timestamp 1682952543
transform 1 0 2184 0 1 3570
box -8 -3 46 105
use INVX2  INVX2_101
timestamp 1682952543
transform 1 0 2224 0 1 3570
box -9 -3 26 105
use M3_M2  M3_M2_1197
timestamp 1682952543
transform 1 0 2332 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_101
timestamp 1682952543
transform 1 0 2240 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_102
timestamp 1682952543
transform 1 0 2336 0 1 3570
box -9 -3 26 105
use OAI22X1  OAI22X1_94
timestamp 1682952543
transform 1 0 2352 0 1 3570
box -8 -3 46 105
use OAI21X1  OAI21X1_1
timestamp 1682952543
transform 1 0 2392 0 1 3570
box -8 -3 34 105
use FILL  FILL_335
timestamp 1682952543
transform 1 0 2424 0 1 3570
box -8 -3 16 105
use FILL  FILL_336
timestamp 1682952543
transform 1 0 2432 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1198
timestamp 1682952543
transform 1 0 2452 0 1 3575
box -3 -3 3 3
use FILL  FILL_337
timestamp 1682952543
transform 1 0 2440 0 1 3570
box -8 -3 16 105
use FILL  FILL_338
timestamp 1682952543
transform 1 0 2448 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_95
timestamp 1682952543
transform 1 0 2456 0 1 3570
box -8 -3 46 105
use FILL  FILL_339
timestamp 1682952543
transform 1 0 2496 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1682952543
transform 1 0 2504 0 1 3570
box -8 -3 34 105
use FILL  FILL_340
timestamp 1682952543
transform 1 0 2536 0 1 3570
box -8 -3 16 105
use FILL  FILL_341
timestamp 1682952543
transform 1 0 2544 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_96
timestamp 1682952543
transform 1 0 2552 0 1 3570
box -8 -3 46 105
use FILL  FILL_342
timestamp 1682952543
transform 1 0 2592 0 1 3570
box -8 -3 16 105
use FILL  FILL_364
timestamp 1682952543
transform 1 0 2600 0 1 3570
box -8 -3 16 105
use FILL  FILL_365
timestamp 1682952543
transform 1 0 2608 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1682952543
transform 1 0 2616 0 1 3570
box -8 -3 34 105
use FILL  FILL_366
timestamp 1682952543
transform 1 0 2648 0 1 3570
box -8 -3 16 105
use FILL  FILL_370
timestamp 1682952543
transform 1 0 2656 0 1 3570
box -8 -3 16 105
use FILL  FILL_371
timestamp 1682952543
transform 1 0 2664 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1199
timestamp 1682952543
transform 1 0 2716 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_102
timestamp 1682952543
transform 1 0 2672 0 1 3570
box -8 -3 46 105
use NAND2X1  NAND2X1_0
timestamp 1682952543
transform 1 0 2712 0 1 3570
box -8 -3 32 105
use OAI21X1  OAI21X1_7
timestamp 1682952543
transform 1 0 2736 0 1 3570
box -8 -3 34 105
use M3_M2  M3_M2_1200
timestamp 1682952543
transform 1 0 2780 0 1 3575
box -3 -3 3 3
use FILL  FILL_372
timestamp 1682952543
transform 1 0 2768 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_8
timestamp 1682952543
transform -1 0 2808 0 1 3570
box -8 -3 34 105
use FILL  FILL_373
timestamp 1682952543
transform 1 0 2808 0 1 3570
box -8 -3 16 105
use FILL  FILL_374
timestamp 1682952543
transform 1 0 2816 0 1 3570
box -8 -3 16 105
use FILL  FILL_375
timestamp 1682952543
transform 1 0 2824 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1682952543
transform 1 0 2832 0 1 3570
box -8 -3 32 105
use FILL  FILL_384
timestamp 1682952543
transform 1 0 2856 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1201
timestamp 1682952543
transform 1 0 2892 0 1 3575
box -3 -3 3 3
use OAI21X1  OAI21X1_10
timestamp 1682952543
transform 1 0 2864 0 1 3570
box -8 -3 34 105
use FILL  FILL_385
timestamp 1682952543
transform 1 0 2896 0 1 3570
box -8 -3 16 105
use FILL  FILL_390
timestamp 1682952543
transform 1 0 2904 0 1 3570
box -8 -3 16 105
use FILL  FILL_391
timestamp 1682952543
transform 1 0 2912 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1202
timestamp 1682952543
transform 1 0 2932 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_1203
timestamp 1682952543
transform 1 0 2956 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_106
timestamp 1682952543
transform -1 0 2960 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_1204
timestamp 1682952543
transform 1 0 2996 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_107
timestamp 1682952543
transform -1 0 3000 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_1205
timestamp 1682952543
transform 1 0 3020 0 1 3575
box -3 -3 3 3
use OAI21X1  OAI21X1_11
timestamp 1682952543
transform 1 0 3000 0 1 3570
box -8 -3 34 105
use M3_M2  M3_M2_1206
timestamp 1682952543
transform 1 0 3068 0 1 3575
box -3 -3 3 3
use OAI21X1  OAI21X1_12
timestamp 1682952543
transform -1 0 3064 0 1 3570
box -8 -3 34 105
use OAI22X1  OAI22X1_108
timestamp 1682952543
transform 1 0 3064 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_1207
timestamp 1682952543
transform 1 0 3140 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_109
timestamp 1682952543
transform -1 0 3144 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_110
timestamp 1682952543
transform -1 0 3184 0 1 3570
box -8 -3 46 105
use INVX2  INVX2_104
timestamp 1682952543
transform 1 0 3184 0 1 3570
box -9 -3 26 105
use FILL  FILL_408
timestamp 1682952543
transform 1 0 3200 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_106
timestamp 1682952543
transform 1 0 3208 0 1 3570
box -9 -3 26 105
use OAI22X1  OAI22X1_113
timestamp 1682952543
transform -1 0 3264 0 1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_114
timestamp 1682952543
transform -1 0 3304 0 1 3570
box -8 -3 46 105
use FILL  FILL_409
timestamp 1682952543
transform 1 0 3304 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1682952543
transform 1 0 3312 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_107
timestamp 1682952543
transform 1 0 3408 0 1 3570
box -9 -3 26 105
use M3_M2  M3_M2_1208
timestamp 1682952543
transform 1 0 3460 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_115
timestamp 1682952543
transform 1 0 3424 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_1209
timestamp 1682952543
transform 1 0 3524 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_105
timestamp 1682952543
transform 1 0 3464 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_108
timestamp 1682952543
transform 1 0 3560 0 1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1682952543
transform 1 0 3576 0 1 3570
box -8 -3 104 105
use INVX2  INVX2_109
timestamp 1682952543
transform 1 0 3672 0 1 3570
box -9 -3 26 105
use FILL  FILL_410
timestamp 1682952543
transform 1 0 3688 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1210
timestamp 1682952543
transform 1 0 3716 0 1 3575
box -3 -3 3 3
use OAI22X1  OAI22X1_120
timestamp 1682952543
transform 1 0 3696 0 1 3570
box -8 -3 46 105
use FILL  FILL_425
timestamp 1682952543
transform 1 0 3736 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1211
timestamp 1682952543
transform 1 0 3756 0 1 3575
box -3 -3 3 3
use FILL  FILL_426
timestamp 1682952543
transform 1 0 3744 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_121
timestamp 1682952543
transform 1 0 3752 0 1 3570
box -8 -3 46 105
use FILL  FILL_427
timestamp 1682952543
transform 1 0 3792 0 1 3570
box -8 -3 16 105
use FILL  FILL_428
timestamp 1682952543
transform 1 0 3800 0 1 3570
box -8 -3 16 105
use FILL  FILL_429
timestamp 1682952543
transform 1 0 3808 0 1 3570
box -8 -3 16 105
use FILL  FILL_430
timestamp 1682952543
transform 1 0 3816 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_19
timestamp 1682952543
transform 1 0 3824 0 1 3570
box -8 -3 34 105
use FILL  FILL_438
timestamp 1682952543
transform 1 0 3856 0 1 3570
box -8 -3 16 105
use FILL  FILL_439
timestamp 1682952543
transform 1 0 3864 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_7
timestamp 1682952543
transform 1 0 3872 0 1 3570
box -8 -3 32 105
use FILL  FILL_440
timestamp 1682952543
transform 1 0 3896 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_8
timestamp 1682952543
transform 1 0 3904 0 1 3570
box -8 -3 32 105
use OAI21X1  OAI21X1_21
timestamp 1682952543
transform -1 0 3960 0 1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_22
timestamp 1682952543
transform -1 0 3992 0 1 3570
box -8 -3 34 105
use M3_M2  M3_M2_1212
timestamp 1682952543
transform 1 0 4004 0 1 3575
box -3 -3 3 3
use NAND2X1  NAND2X1_9
timestamp 1682952543
transform 1 0 3992 0 1 3570
box -8 -3 32 105
use OAI22X1  OAI22X1_123
timestamp 1682952543
transform 1 0 4016 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_1213
timestamp 1682952543
transform 1 0 4140 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_107
timestamp 1682952543
transform 1 0 4056 0 1 3570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_11
timestamp 1682952543
transform 1 0 4177 0 1 3570
box -10 -3 10 3
use M3_M2  M3_M2_1246
timestamp 1682952543
transform 1 0 84 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1682952543
transform 1 0 180 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1294
timestamp 1682952543
transform 1 0 164 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1294
timestamp 1682952543
transform 1 0 84 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1247
timestamp 1682952543
transform 1 0 196 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1682952543
transform 1 0 212 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1295
timestamp 1682952543
transform 1 0 188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1296
timestamp 1682952543
transform 1 0 196 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1682952543
transform 1 0 212 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1437
timestamp 1682952543
transform 1 0 116 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1682952543
transform 1 0 164 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1682952543
transform 1 0 172 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1682952543
transform 1 0 180 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1399
timestamp 1682952543
transform 1 0 148 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1442
timestamp 1682952543
transform 1 0 164 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1358
timestamp 1682952543
transform 1 0 196 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1298
timestamp 1682952543
transform 1 0 236 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1299
timestamp 1682952543
transform 1 0 252 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1682952543
transform 1 0 260 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1682952543
transform 1 0 204 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1682952543
transform 1 0 220 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1682952543
transform 1 0 228 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1359
timestamp 1682952543
transform 1 0 236 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1444
timestamp 1682952543
transform 1 0 244 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1360
timestamp 1682952543
transform 1 0 252 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1445
timestamp 1682952543
transform 1 0 260 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1400
timestamp 1682952543
transform 1 0 204 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1682952543
transform 1 0 220 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1682952543
transform 1 0 260 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1682952543
transform 1 0 228 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1490
timestamp 1682952543
transform 1 0 260 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1682952543
transform 1 0 292 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1301
timestamp 1682952543
transform 1 0 292 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1682952543
transform 1 0 276 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1447
timestamp 1682952543
transform 1 0 316 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1361
timestamp 1682952543
transform 1 0 364 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1682952543
transform 1 0 396 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1248
timestamp 1682952543
transform 1 0 404 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1324
timestamp 1682952543
transform 1 0 388 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1296
timestamp 1682952543
transform 1 0 420 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1302
timestamp 1682952543
transform 1 0 396 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1682952543
transform 1 0 412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1682952543
transform 1 0 420 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1448
timestamp 1682952543
transform 1 0 372 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1682952543
transform 1 0 388 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1450
timestamp 1682952543
transform 1 0 404 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1403
timestamp 1682952543
transform 1 0 276 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1682952543
transform 1 0 316 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1682952543
transform 1 0 300 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1682952543
transform 1 0 412 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1362
timestamp 1682952543
transform 1 0 428 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1682952543
transform 1 0 444 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1297
timestamp 1682952543
transform 1 0 452 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1305
timestamp 1682952543
transform 1 0 452 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1325
timestamp 1682952543
transform 1 0 460 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1306
timestamp 1682952543
transform 1 0 468 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1682952543
transform 1 0 436 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1363
timestamp 1682952543
transform 1 0 452 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1452
timestamp 1682952543
transform 1 0 460 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1405
timestamp 1682952543
transform 1 0 436 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1250
timestamp 1682952543
transform 1 0 500 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1307
timestamp 1682952543
transform 1 0 508 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1326
timestamp 1682952543
transform 1 0 516 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1308
timestamp 1682952543
transform 1 0 532 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1327
timestamp 1682952543
transform 1 0 556 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1309
timestamp 1682952543
transform 1 0 620 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1682952543
transform 1 0 628 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1682952543
transform 1 0 644 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1312
timestamp 1682952543
transform 1 0 652 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1453
timestamp 1682952543
transform 1 0 516 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1454
timestamp 1682952543
transform 1 0 556 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1455
timestamp 1682952543
transform 1 0 612 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1682952543
transform 1 0 636 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1444
timestamp 1682952543
transform 1 0 508 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1682952543
transform 1 0 644 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1457
timestamp 1682952543
transform 1 0 652 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1445
timestamp 1682952543
transform 1 0 556 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1446
timestamp 1682952543
transform 1 0 620 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1474
timestamp 1682952543
transform 1 0 604 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1682952543
transform 1 0 572 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1493
timestamp 1682952543
transform 1 0 588 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1682952543
transform 1 0 652 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_1458
timestamp 1682952543
transform 1 0 668 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1251
timestamp 1682952543
transform 1 0 700 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1682952543
transform 1 0 700 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1252
timestamp 1682952543
transform 1 0 732 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1313
timestamp 1682952543
transform 1 0 724 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1459
timestamp 1682952543
transform 1 0 748 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1682952543
transform 1 0 780 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1315
timestamp 1682952543
transform 1 0 788 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1366
timestamp 1682952543
transform 1 0 788 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1460
timestamp 1682952543
transform 1 0 796 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1406
timestamp 1682952543
transform 1 0 780 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_1316
timestamp 1682952543
transform 1 0 820 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1461
timestamp 1682952543
transform 1 0 828 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1447
timestamp 1682952543
transform 1 0 804 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1217
timestamp 1682952543
transform 1 0 844 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1288
timestamp 1682952543
transform 1 0 844 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1682952543
transform 1 0 844 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1682952543
transform 1 0 876 0 1 3545
box -2 -2 2 2
use M3_M2  M3_M2_1218
timestamp 1682952543
transform 1 0 892 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1298
timestamp 1682952543
transform 1 0 892 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1318
timestamp 1682952543
transform 1 0 884 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1462
timestamp 1682952543
transform 1 0 892 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1253
timestamp 1682952543
transform 1 0 908 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1290
timestamp 1682952543
transform 1 0 908 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1682952543
transform 1 0 908 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1682952543
transform 1 0 940 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1682952543
transform 1 0 932 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1682952543
transform 1 0 924 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1328
timestamp 1682952543
transform 1 0 940 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1682952543
transform 1 0 956 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1464
timestamp 1682952543
transform 1 0 948 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1682952543
transform 1 0 980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1682952543
transform 1 0 988 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1254
timestamp 1682952543
transform 1 0 1084 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1322
timestamp 1682952543
transform 1 0 1004 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1329
timestamp 1682952543
transform 1 0 1036 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1330
timestamp 1682952543
transform 1 0 1092 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1331
timestamp 1682952543
transform 1 0 1108 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1255
timestamp 1682952543
transform 1 0 1140 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1682952543
transform 1 0 1180 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1682952543
transform 1 0 1188 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1257
timestamp 1682952543
transform 1 0 1236 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1323
timestamp 1682952543
transform 1 0 1116 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1682952543
transform 1 0 1124 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1682952543
transform 1 0 1140 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1682952543
transform 1 0 1148 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1682952543
transform 1 0 1156 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1682952543
transform 1 0 1180 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1329
timestamp 1682952543
transform 1 0 1188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1330
timestamp 1682952543
transform 1 0 1212 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1682952543
transform 1 0 1036 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1682952543
transform 1 0 1084 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1468
timestamp 1682952543
transform 1 0 1092 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1682952543
transform 1 0 1100 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1682952543
transform 1 0 1108 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1407
timestamp 1682952543
transform 1 0 1100 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1682952543
transform 1 0 1124 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1471
timestamp 1682952543
transform 1 0 1132 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1682952543
transform 1 0 1156 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1368
timestamp 1682952543
transform 1 0 1164 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1473
timestamp 1682952543
transform 1 0 1172 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1369
timestamp 1682952543
transform 1 0 1180 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1332
timestamp 1682952543
transform 1 0 1220 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1682952543
transform 1 0 1340 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1682952543
transform 1 0 1356 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1258
timestamp 1682952543
transform 1 0 1292 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1259
timestamp 1682952543
transform 1 0 1324 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1331
timestamp 1682952543
transform 1 0 1228 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1332
timestamp 1682952543
transform 1 0 1236 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1333
timestamp 1682952543
transform 1 0 1244 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1333
timestamp 1682952543
transform 1 0 1260 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1334
timestamp 1682952543
transform 1 0 1284 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1260
timestamp 1682952543
transform 1 0 1356 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1334
timestamp 1682952543
transform 1 0 1348 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1682952543
transform 1 0 1356 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1682952543
transform 1 0 1372 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1682952543
transform 1 0 1380 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1474
timestamp 1682952543
transform 1 0 1188 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1682952543
transform 1 0 1204 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1682952543
transform 1 0 1220 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1370
timestamp 1682952543
transform 1 0 1236 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1477
timestamp 1682952543
transform 1 0 1244 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1478
timestamp 1682952543
transform 1 0 1284 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1479
timestamp 1682952543
transform 1 0 1340 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1480
timestamp 1682952543
transform 1 0 1364 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1481
timestamp 1682952543
transform 1 0 1388 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1408
timestamp 1682952543
transform 1 0 1148 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1682952543
transform 1 0 1188 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1410
timestamp 1682952543
transform 1 0 1220 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1682952543
transform 1 0 1156 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1448
timestamp 1682952543
transform 1 0 1228 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1495
timestamp 1682952543
transform 1 0 1196 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1449
timestamp 1682952543
transform 1 0 1372 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1476
timestamp 1682952543
transform 1 0 1372 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1682952543
transform 1 0 1276 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1497
timestamp 1682952543
transform 1 0 1348 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1682952543
transform 1 0 1380 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1261
timestamp 1682952543
transform 1 0 1420 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1682952543
transform 1 0 1500 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1335
timestamp 1682952543
transform 1 0 1396 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1336
timestamp 1682952543
transform 1 0 1436 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1263
timestamp 1682952543
transform 1 0 1532 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1338
timestamp 1682952543
transform 1 0 1484 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1682952543
transform 1 0 1500 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1682952543
transform 1 0 1516 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1482
timestamp 1682952543
transform 1 0 1396 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1682952543
transform 1 0 1404 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1484
timestamp 1682952543
transform 1 0 1436 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1485
timestamp 1682952543
transform 1 0 1508 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1486
timestamp 1682952543
transform 1 0 1524 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1411
timestamp 1682952543
transform 1 0 1524 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1450
timestamp 1682952543
transform 1 0 1404 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1451
timestamp 1682952543
transform 1 0 1420 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1452
timestamp 1682952543
transform 1 0 1492 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1499
timestamp 1682952543
transform 1 0 1476 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1682952543
transform 1 0 1500 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1264
timestamp 1682952543
transform 1 0 1548 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1299
timestamp 1682952543
transform 1 0 1572 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1341
timestamp 1682952543
transform 1 0 1548 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1342
timestamp 1682952543
transform 1 0 1556 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1682952543
transform 1 0 1572 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1371
timestamp 1682952543
transform 1 0 1556 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1487
timestamp 1682952543
transform 1 0 1564 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1488
timestamp 1682952543
transform 1 0 1580 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1223
timestamp 1682952543
transform 1 0 1596 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1489
timestamp 1682952543
transform 1 0 1596 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1300
timestamp 1682952543
transform 1 0 1612 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1301
timestamp 1682952543
transform 1 0 1636 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1682952543
transform 1 0 1652 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1344
timestamp 1682952543
transform 1 0 1612 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1682952543
transform 1 0 1620 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1337
timestamp 1682952543
transform 1 0 1628 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1346
timestamp 1682952543
transform 1 0 1636 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1682952543
transform 1 0 1644 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1338
timestamp 1682952543
transform 1 0 1660 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1348
timestamp 1682952543
transform 1 0 1732 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1682952543
transform 1 0 1748 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1490
timestamp 1682952543
transform 1 0 1628 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1491
timestamp 1682952543
transform 1 0 1652 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1492
timestamp 1682952543
transform 1 0 1684 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1477
timestamp 1682952543
transform 1 0 1612 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1682952543
transform 1 0 1748 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1224
timestamp 1682952543
transform 1 0 1788 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1303
timestamp 1682952543
transform 1 0 1780 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1350
timestamp 1682952543
transform 1 0 1780 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1351
timestamp 1682952543
transform 1 0 1788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1352
timestamp 1682952543
transform 1 0 1796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1493
timestamp 1682952543
transform 1 0 1756 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1494
timestamp 1682952543
transform 1 0 1772 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1453
timestamp 1682952543
transform 1 0 1732 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1412
timestamp 1682952543
transform 1 0 1772 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1682952543
transform 1 0 1796 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1454
timestamp 1682952543
transform 1 0 1772 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1304
timestamp 1682952543
transform 1 0 1812 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1353
timestamp 1682952543
transform 1 0 1900 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1682952543
transform 1 0 1812 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1496
timestamp 1682952543
transform 1 0 1820 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1414
timestamp 1682952543
transform 1 0 1812 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1373
timestamp 1682952543
transform 1 0 1828 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1497
timestamp 1682952543
transform 1 0 1860 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1374
timestamp 1682952543
transform 1 0 1900 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1682952543
transform 1 0 1860 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1265
timestamp 1682952543
transform 1 0 1916 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1354
timestamp 1682952543
transform 1 0 1916 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1375
timestamp 1682952543
transform 1 0 1924 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1355
timestamp 1682952543
transform 1 0 1964 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1682952543
transform 1 0 1940 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1455
timestamp 1682952543
transform 1 0 1932 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1682952543
transform 1 0 1948 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1499
timestamp 1682952543
transform 1 0 1956 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1377
timestamp 1682952543
transform 1 0 1964 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1356
timestamp 1682952543
transform 1 0 1980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1500
timestamp 1682952543
transform 1 0 1972 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1416
timestamp 1682952543
transform 1 0 1956 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1682952543
transform 1 0 1948 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1682952543
transform 1 0 1980 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1456
timestamp 1682952543
transform 1 0 1980 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1225
timestamp 1682952543
transform 1 0 2076 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1682952543
transform 1 0 2132 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1227
timestamp 1682952543
transform 1 0 2172 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1266
timestamp 1682952543
transform 1 0 2020 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1682952543
transform 1 0 2068 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1682952543
transform 1 0 2108 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1682952543
transform 1 0 2140 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1270
timestamp 1682952543
transform 1 0 2188 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1682952543
transform 1 0 2036 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1306
timestamp 1682952543
transform 1 0 2100 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1357
timestamp 1682952543
transform 1 0 2100 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1501
timestamp 1682952543
transform 1 0 2012 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1502
timestamp 1682952543
transform 1 0 2020 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1503
timestamp 1682952543
transform 1 0 2052 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1418
timestamp 1682952543
transform 1 0 2012 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1682952543
transform 1 0 2052 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1457
timestamp 1682952543
transform 1 0 2004 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1682952543
transform 1 0 1996 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1458
timestamp 1682952543
transform 1 0 2052 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1502
timestamp 1682952543
transform 1 0 2044 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1682952543
transform 1 0 2172 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1358
timestamp 1682952543
transform 1 0 2124 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1378
timestamp 1682952543
transform 1 0 2124 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1682952543
transform 1 0 2156 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1228
timestamp 1682952543
transform 1 0 2212 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1504
timestamp 1682952543
transform 1 0 2172 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1682952543
transform 1 0 2204 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1271
timestamp 1682952543
transform 1 0 2220 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1682952543
transform 1 0 2276 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1308
timestamp 1682952543
transform 1 0 2244 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1682952543
transform 1 0 2260 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1310
timestamp 1682952543
transform 1 0 2300 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1359
timestamp 1682952543
transform 1 0 2228 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1682952543
transform 1 0 2244 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1682952543
transform 1 0 2260 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1682952543
transform 1 0 2268 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1363
timestamp 1682952543
transform 1 0 2284 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1682952543
transform 1 0 2300 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1365
timestamp 1682952543
transform 1 0 2308 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1682952543
transform 1 0 2220 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1420
timestamp 1682952543
transform 1 0 2220 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_1507
timestamp 1682952543
transform 1 0 2252 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1479
timestamp 1682952543
transform 1 0 2252 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_1508
timestamp 1682952543
transform 1 0 2276 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1682952543
transform 1 0 2292 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1421
timestamp 1682952543
transform 1 0 2308 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1230
timestamp 1682952543
transform 1 0 2348 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1272
timestamp 1682952543
transform 1 0 2332 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1682952543
transform 1 0 2356 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1459
timestamp 1682952543
transform 1 0 2324 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1682952543
transform 1 0 2324 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_1366
timestamp 1682952543
transform 1 0 2348 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1367
timestamp 1682952543
transform 1 0 2364 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1368
timestamp 1682952543
transform 1 0 2372 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1682952543
transform 1 0 2340 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1682952543
transform 1 0 2356 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1422
timestamp 1682952543
transform 1 0 2356 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_1512
timestamp 1682952543
transform 1 0 2388 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1423
timestamp 1682952543
transform 1 0 2380 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1460
timestamp 1682952543
transform 1 0 2388 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1274
timestamp 1682952543
transform 1 0 2428 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1369
timestamp 1682952543
transform 1 0 2412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1370
timestamp 1682952543
transform 1 0 2428 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1565
timestamp 1682952543
transform 1 0 2412 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1481
timestamp 1682952543
transform 1 0 2404 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1503
timestamp 1682952543
transform 1 0 2404 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1339
timestamp 1682952543
transform 1 0 2436 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1371
timestamp 1682952543
transform 1 0 2444 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1340
timestamp 1682952543
transform 1 0 2452 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1372
timestamp 1682952543
transform 1 0 2460 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1682952543
transform 1 0 2468 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1513
timestamp 1682952543
transform 1 0 2436 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1380
timestamp 1682952543
transform 1 0 2444 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1514
timestamp 1682952543
transform 1 0 2452 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1424
timestamp 1682952543
transform 1 0 2452 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1682952543
transform 1 0 2436 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1682952543
transform 1 0 2468 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1231
timestamp 1682952543
transform 1 0 2508 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1275
timestamp 1682952543
transform 1 0 2492 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1276
timestamp 1682952543
transform 1 0 2508 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1515
timestamp 1682952543
transform 1 0 2484 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1374
timestamp 1682952543
transform 1 0 2508 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1375
timestamp 1682952543
transform 1 0 2516 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1682952543
transform 1 0 2516 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1682952543
transform 1 0 2508 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1425
timestamp 1682952543
transform 1 0 2516 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1682952543
transform 1 0 2524 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1682952543
transform 1 0 2556 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1376
timestamp 1682952543
transform 1 0 2548 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1682952543
transform 1 0 2564 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1682952543
transform 1 0 2572 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1682952543
transform 1 0 2556 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1462
timestamp 1682952543
transform 1 0 2556 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_1518
timestamp 1682952543
transform 1 0 2604 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1341
timestamp 1682952543
transform 1 0 2628 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1519
timestamp 1682952543
transform 1 0 2628 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1682952543
transform 1 0 2628 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1233
timestamp 1682952543
transform 1 0 2644 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1379
timestamp 1682952543
transform 1 0 2644 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1380
timestamp 1682952543
transform 1 0 2652 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1463
timestamp 1682952543
transform 1 0 2644 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1342
timestamp 1682952543
transform 1 0 2668 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1381
timestamp 1682952543
transform 1 0 2676 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1682952543
transform 1 0 2692 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1682952543
transform 1 0 2700 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1682952543
transform 1 0 2668 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1382
timestamp 1682952543
transform 1 0 2676 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1521
timestamp 1682952543
transform 1 0 2684 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1426
timestamp 1682952543
transform 1 0 2676 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1427
timestamp 1682952543
transform 1 0 2692 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1505
timestamp 1682952543
transform 1 0 2684 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1343
timestamp 1682952543
transform 1 0 2708 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1522
timestamp 1682952543
transform 1 0 2708 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1428
timestamp 1682952543
transform 1 0 2716 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1682952543
transform 1 0 2756 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1523
timestamp 1682952543
transform 1 0 2756 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1429
timestamp 1682952543
transform 1 0 2740 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1430
timestamp 1682952543
transform 1 0 2756 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_1384
timestamp 1682952543
transform 1 0 2764 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1277
timestamp 1682952543
transform 1 0 2788 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1385
timestamp 1682952543
transform 1 0 2788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1386
timestamp 1682952543
transform 1 0 2804 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1568
timestamp 1682952543
transform 1 0 2780 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1682952543
transform 1 0 2796 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1682952543
transform 1 0 2812 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1383
timestamp 1682952543
transform 1 0 2820 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1278
timestamp 1682952543
transform 1 0 2844 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1387
timestamp 1682952543
transform 1 0 2836 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1235
timestamp 1682952543
transform 1 0 2892 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1279
timestamp 1682952543
transform 1 0 2884 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1682952543
transform 1 0 2860 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1388
timestamp 1682952543
transform 1 0 2868 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1389
timestamp 1682952543
transform 1 0 2884 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1682952543
transform 1 0 2892 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1682952543
transform 1 0 2860 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1682952543
transform 1 0 2876 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1431
timestamp 1682952543
transform 1 0 2876 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1682952543
transform 1 0 2860 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1236
timestamp 1682952543
transform 1 0 2908 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1432
timestamp 1682952543
transform 1 0 2916 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_1569
timestamp 1682952543
transform 1 0 2924 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1433
timestamp 1682952543
transform 1 0 2940 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1507
timestamp 1682952543
transform 1 0 2932 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1682952543
transform 1 0 2956 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1682952543
transform 1 0 2972 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1682952543
transform 1 0 2980 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1391
timestamp 1682952543
transform 1 0 2956 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1392
timestamp 1682952543
transform 1 0 2972 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1682952543
transform 1 0 2948 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1682952543
transform 1 0 2964 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1384
timestamp 1682952543
transform 1 0 2972 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1530
timestamp 1682952543
transform 1 0 2980 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1434
timestamp 1682952543
transform 1 0 2964 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1682952543
transform 1 0 3004 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_1393
timestamp 1682952543
transform 1 0 2996 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1508
timestamp 1682952543
transform 1 0 2988 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_1394
timestamp 1682952543
transform 1 0 3012 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1345
timestamp 1682952543
transform 1 0 3020 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1531
timestamp 1682952543
transform 1 0 3012 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1240
timestamp 1682952543
transform 1 0 3044 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1346
timestamp 1682952543
transform 1 0 3036 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1395
timestamp 1682952543
transform 1 0 3044 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1682952543
transform 1 0 3028 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1464
timestamp 1682952543
transform 1 0 3036 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1682952543
transform 1 0 3044 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1682952543
transform 1 0 3076 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1682952543
transform 1 0 3076 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1571
timestamp 1682952543
transform 1 0 3076 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1385
timestamp 1682952543
transform 1 0 3092 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1682952543
transform 1 0 3108 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1396
timestamp 1682952543
transform 1 0 3100 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1348
timestamp 1682952543
transform 1 0 3108 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1397
timestamp 1682952543
transform 1 0 3124 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1398
timestamp 1682952543
transform 1 0 3140 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1399
timestamp 1682952543
transform 1 0 3148 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1532
timestamp 1682952543
transform 1 0 3100 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1533
timestamp 1682952543
transform 1 0 3116 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1534
timestamp 1682952543
transform 1 0 3132 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1509
timestamp 1682952543
transform 1 0 3116 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1283
timestamp 1682952543
transform 1 0 3180 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1241
timestamp 1682952543
transform 1 0 3196 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1284
timestamp 1682952543
transform 1 0 3204 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1285
timestamp 1682952543
transform 1 0 3220 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1400
timestamp 1682952543
transform 1 0 3188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1401
timestamp 1682952543
transform 1 0 3204 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1349
timestamp 1682952543
transform 1 0 3212 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1402
timestamp 1682952543
transform 1 0 3220 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1403
timestamp 1682952543
transform 1 0 3236 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1404
timestamp 1682952543
transform 1 0 3244 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1286
timestamp 1682952543
transform 1 0 3276 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_1405
timestamp 1682952543
transform 1 0 3268 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1682952543
transform 1 0 3276 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1535
timestamp 1682952543
transform 1 0 3196 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1682952543
transform 1 0 3212 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1386
timestamp 1682952543
transform 1 0 3220 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1537
timestamp 1682952543
transform 1 0 3228 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1387
timestamp 1682952543
transform 1 0 3244 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1538
timestamp 1682952543
transform 1 0 3252 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1388
timestamp 1682952543
transform 1 0 3268 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1539
timestamp 1682952543
transform 1 0 3284 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1389
timestamp 1682952543
transform 1 0 3292 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1435
timestamp 1682952543
transform 1 0 3228 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1465
timestamp 1682952543
transform 1 0 3196 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1483
timestamp 1682952543
transform 1 0 3188 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_1572
timestamp 1682952543
transform 1 0 3268 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1510
timestamp 1682952543
transform 1 0 3252 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1511
timestamp 1682952543
transform 1 0 3268 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_1573
timestamp 1682952543
transform 1 0 3300 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1466
timestamp 1682952543
transform 1 0 3300 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_1540
timestamp 1682952543
transform 1 0 3324 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1682952543
transform 1 0 3332 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1484
timestamp 1682952543
transform 1 0 3332 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1682952543
transform 1 0 3372 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1407
timestamp 1682952543
transform 1 0 3388 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1408
timestamp 1682952543
transform 1 0 3396 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1682952543
transform 1 0 3380 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1682952543
transform 1 0 3388 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1351
timestamp 1682952543
transform 1 0 3404 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1409
timestamp 1682952543
transform 1 0 3412 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1352
timestamp 1682952543
transform 1 0 3420 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1311
timestamp 1682952543
transform 1 0 3468 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1312
timestamp 1682952543
transform 1 0 3492 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1410
timestamp 1682952543
transform 1 0 3428 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1411
timestamp 1682952543
transform 1 0 3436 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1682952543
transform 1 0 3452 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1413
timestamp 1682952543
transform 1 0 3468 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1682952543
transform 1 0 3476 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1682952543
transform 1 0 3492 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1416
timestamp 1682952543
transform 1 0 3508 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1543
timestamp 1682952543
transform 1 0 3404 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1390
timestamp 1682952543
transform 1 0 3412 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1544
timestamp 1682952543
transform 1 0 3420 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1436
timestamp 1682952543
transform 1 0 3420 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1485
timestamp 1682952543
transform 1 0 3420 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_1545
timestamp 1682952543
transform 1 0 3444 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1546
timestamp 1682952543
transform 1 0 3460 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1682952543
transform 1 0 3484 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1391
timestamp 1682952543
transform 1 0 3492 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1548
timestamp 1682952543
transform 1 0 3500 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1392
timestamp 1682952543
transform 1 0 3508 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1549
timestamp 1682952543
transform 1 0 3516 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1242
timestamp 1682952543
transform 1 0 3524 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1313
timestamp 1682952543
transform 1 0 3532 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1417
timestamp 1682952543
transform 1 0 3524 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1682952543
transform 1 0 3532 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1437
timestamp 1682952543
transform 1 0 3444 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1438
timestamp 1682952543
transform 1 0 3476 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1682952543
transform 1 0 3516 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1486
timestamp 1682952543
transform 1 0 3500 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_1550
timestamp 1682952543
transform 1 0 3540 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1243
timestamp 1682952543
transform 1 0 3556 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1287
timestamp 1682952543
transform 1 0 3580 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1467
timestamp 1682952543
transform 1 0 3572 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_1575
timestamp 1682952543
transform 1 0 3580 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1512
timestamp 1682952543
transform 1 0 3580 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_1393
timestamp 1682952543
transform 1 0 3604 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1551
timestamp 1682952543
transform 1 0 3612 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1682952543
transform 1 0 3636 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1487
timestamp 1682952543
transform 1 0 3636 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_1577
timestamp 1682952543
transform 1 0 3652 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1488
timestamp 1682952543
transform 1 0 3652 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_1552
timestamp 1682952543
transform 1 0 3676 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1682952543
transform 1 0 3708 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_1419
timestamp 1682952543
transform 1 0 3708 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1682952543
transform 1 0 3732 0 1 3545
box -2 -2 2 2
use M3_M2  M3_M2_1314
timestamp 1682952543
transform 1 0 3756 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1420
timestamp 1682952543
transform 1 0 3740 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1353
timestamp 1682952543
transform 1 0 3748 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1315
timestamp 1682952543
transform 1 0 3780 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1421
timestamp 1682952543
transform 1 0 3756 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1422
timestamp 1682952543
transform 1 0 3772 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1682952543
transform 1 0 3780 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1553
timestamp 1682952543
transform 1 0 3748 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1682952543
transform 1 0 3764 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1394
timestamp 1682952543
transform 1 0 3772 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_1440
timestamp 1682952543
transform 1 0 3764 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1468
timestamp 1682952543
transform 1 0 3748 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1682952543
transform 1 0 3788 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1555
timestamp 1682952543
transform 1 0 3788 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1578
timestamp 1682952543
transform 1 0 3812 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1489
timestamp 1682952543
transform 1 0 3812 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_1288
timestamp 1682952543
transform 1 0 3852 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1682952543
transform 1 0 3868 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1682952543
transform 1 0 3844 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1424
timestamp 1682952543
transform 1 0 3844 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1682952543
transform 1 0 3852 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1317
timestamp 1682952543
transform 1 0 3876 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1426
timestamp 1682952543
transform 1 0 3876 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1395
timestamp 1682952543
transform 1 0 3876 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1427
timestamp 1682952543
transform 1 0 3908 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1556
timestamp 1682952543
transform 1 0 3900 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1290
timestamp 1682952543
transform 1 0 3948 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1291
timestamp 1682952543
transform 1 0 3988 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1682952543
transform 1 0 3940 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1682952543
transform 1 0 3964 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1682952543
transform 1 0 3980 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1428
timestamp 1682952543
transform 1 0 3940 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1682952543
transform 1 0 3948 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1355
timestamp 1682952543
transform 1 0 3956 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_1321
timestamp 1682952543
transform 1 0 4020 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1430
timestamp 1682952543
transform 1 0 3964 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1682952543
transform 1 0 3980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1432
timestamp 1682952543
transform 1 0 3988 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1356
timestamp 1682952543
transform 1 0 3996 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1433
timestamp 1682952543
transform 1 0 4004 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1357
timestamp 1682952543
transform 1 0 4012 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_1434
timestamp 1682952543
transform 1 0 4020 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1557
timestamp 1682952543
transform 1 0 3932 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1682952543
transform 1 0 3940 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1682952543
transform 1 0 3972 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1682952543
transform 1 0 3916 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_1396
timestamp 1682952543
transform 1 0 3980 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1560
timestamp 1682952543
transform 1 0 3988 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1682952543
transform 1 0 4012 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1682952543
transform 1 0 4028 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1441
timestamp 1682952543
transform 1 0 3972 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1682952543
transform 1 0 3924 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1470
timestamp 1682952543
transform 1 0 3940 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1682952543
transform 1 0 4052 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1245
timestamp 1682952543
transform 1 0 4084 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_1292
timestamp 1682952543
transform 1 0 4044 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1293
timestamp 1682952543
transform 1 0 4116 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_1322
timestamp 1682952543
transform 1 0 4036 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_1435
timestamp 1682952543
transform 1 0 4036 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1682952543
transform 1 0 4052 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_1397
timestamp 1682952543
transform 1 0 4052 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1563
timestamp 1682952543
transform 1 0 4076 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1398
timestamp 1682952543
transform 1 0 4092 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_1564
timestamp 1682952543
transform 1 0 4132 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_1471
timestamp 1682952543
transform 1 0 4044 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1472
timestamp 1682952543
transform 1 0 4076 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1682952543
transform 1 0 4148 0 1 3545
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_12
timestamp 1682952543
transform 1 0 24 0 1 3470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_84
timestamp 1682952543
transform 1 0 72 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_83
timestamp 1682952543
transform -1 0 184 0 -1 3570
box -9 -3 26 105
use AOI22X1  AOI22X1_37
timestamp 1682952543
transform 1 0 184 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_38
timestamp 1682952543
transform 1 0 224 0 -1 3570
box -8 -3 46 105
use INVX2  INVX2_84
timestamp 1682952543
transform 1 0 264 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1682952543
transform 1 0 280 0 -1 3570
box -8 -3 104 105
use OAI22X1  OAI22X1_81
timestamp 1682952543
transform 1 0 376 0 -1 3570
box -8 -3 46 105
use FILL  FILL_274
timestamp 1682952543
transform 1 0 416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_277
timestamp 1682952543
transform 1 0 424 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_83
timestamp 1682952543
transform 1 0 432 0 -1 3570
box -8 -3 46 105
use FILL  FILL_278
timestamp 1682952543
transform 1 0 472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_280
timestamp 1682952543
transform 1 0 480 0 -1 3570
box -8 -3 16 105
use FILL  FILL_285
timestamp 1682952543
transform 1 0 488 0 -1 3570
box -8 -3 16 105
use FILL  FILL_286
timestamp 1682952543
transform 1 0 496 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_85
timestamp 1682952543
transform 1 0 504 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1682952543
transform 1 0 520 0 -1 3570
box -8 -3 104 105
use AOI22X1  AOI22X1_40
timestamp 1682952543
transform 1 0 616 0 -1 3570
box -8 -3 46 105
use FILL  FILL_298
timestamp 1682952543
transform 1 0 656 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_90
timestamp 1682952543
transform 1 0 664 0 -1 3570
box -9 -3 26 105
use FILL  FILL_299
timestamp 1682952543
transform 1 0 680 0 -1 3570
box -8 -3 16 105
use FILL  FILL_300
timestamp 1682952543
transform 1 0 688 0 -1 3570
box -8 -3 16 105
use FILL  FILL_301
timestamp 1682952543
transform 1 0 696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_302
timestamp 1682952543
transform 1 0 704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_303
timestamp 1682952543
transform 1 0 712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_304
timestamp 1682952543
transform 1 0 720 0 -1 3570
box -8 -3 16 105
use BUFX2  BUFX2_3
timestamp 1682952543
transform -1 0 752 0 -1 3570
box -5 -3 28 105
use FILL  FILL_305
timestamp 1682952543
transform 1 0 752 0 -1 3570
box -8 -3 16 105
use BUFX2  BUFX2_4
timestamp 1682952543
transform 1 0 760 0 -1 3570
box -5 -3 28 105
use FILL  FILL_306
timestamp 1682952543
transform 1 0 784 0 -1 3570
box -8 -3 16 105
use FILL  FILL_307
timestamp 1682952543
transform 1 0 792 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_87
timestamp 1682952543
transform 1 0 800 0 -1 3570
box -8 -3 46 105
use FILL  FILL_308
timestamp 1682952543
transform 1 0 840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_309
timestamp 1682952543
transform 1 0 848 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_9
timestamp 1682952543
transform 1 0 856 0 -1 3570
box -8 -3 32 105
use FILL  FILL_310
timestamp 1682952543
transform 1 0 880 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1682952543
transform 1 0 888 0 -1 3570
box -8 -3 32 105
use FILL  FILL_311
timestamp 1682952543
transform 1 0 912 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_11
timestamp 1682952543
transform 1 0 920 0 -1 3570
box -8 -3 32 105
use FILL  FILL_312
timestamp 1682952543
transform 1 0 944 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1682952543
transform 1 0 952 0 -1 3570
box -8 -3 32 105
use M3_M2  M3_M2_1513
timestamp 1682952543
transform 1 0 988 0 1 3475
box -3 -3 3 3
use FILL  FILL_313
timestamp 1682952543
transform 1 0 976 0 -1 3570
box -8 -3 16 105
use FILL  FILL_314
timestamp 1682952543
transform 1 0 984 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1682952543
transform 1 0 992 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_91
timestamp 1682952543
transform -1 0 1104 0 -1 3570
box -9 -3 26 105
use FILL  FILL_315
timestamp 1682952543
transform 1 0 1104 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_44
timestamp 1682952543
transform 1 0 1112 0 -1 3570
box -8 -3 46 105
use AOI22X1  AOI22X1_45
timestamp 1682952543
transform 1 0 1152 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_88
timestamp 1682952543
transform -1 0 1232 0 -1 3570
box -8 -3 46 105
use INVX2  INVX2_92
timestamp 1682952543
transform 1 0 1232 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1682952543
transform 1 0 1248 0 -1 3570
box -8 -3 104 105
use AOI22X1  AOI22X1_46
timestamp 1682952543
transform 1 0 1344 0 -1 3570
box -8 -3 46 105
use INVX2  INVX2_94
timestamp 1682952543
transform 1 0 1384 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1682952543
transform -1 0 1496 0 -1 3570
box -8 -3 104 105
use M3_M2  M3_M2_1514
timestamp 1682952543
transform 1 0 1516 0 1 3475
box -3 -3 3 3
use OAI22X1  OAI22X1_91
timestamp 1682952543
transform -1 0 1536 0 -1 3570
box -8 -3 46 105
use FILL  FILL_323
timestamp 1682952543
transform 1 0 1536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_324
timestamp 1682952543
transform 1 0 1544 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_92
timestamp 1682952543
transform 1 0 1552 0 -1 3570
box -8 -3 46 105
use FILL  FILL_325
timestamp 1682952543
transform 1 0 1592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_326
timestamp 1682952543
transform 1 0 1600 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_50
timestamp 1682952543
transform 1 0 1608 0 -1 3570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_97
timestamp 1682952543
transform -1 0 1744 0 -1 3570
box -8 -3 104 105
use FILL  FILL_327
timestamp 1682952543
transform 1 0 1744 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_51
timestamp 1682952543
transform -1 0 1792 0 -1 3570
box -8 -3 46 105
use INVX2  INVX2_98
timestamp 1682952543
transform 1 0 1792 0 -1 3570
box -9 -3 26 105
use FILL  FILL_328
timestamp 1682952543
transform 1 0 1808 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1682952543
transform -1 0 1912 0 -1 3570
box -8 -3 104 105
use FILL  FILL_329
timestamp 1682952543
transform 1 0 1912 0 -1 3570
box -8 -3 16 105
use FILL  FILL_343
timestamp 1682952543
transform 1 0 1920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_344
timestamp 1682952543
transform 1 0 1928 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_52
timestamp 1682952543
transform -1 0 1976 0 -1 3570
box -8 -3 46 105
use FILL  FILL_345
timestamp 1682952543
transform 1 0 1976 0 -1 3570
box -8 -3 16 105
use FILL  FILL_346
timestamp 1682952543
transform 1 0 1984 0 -1 3570
box -8 -3 16 105
use FILL  FILL_347
timestamp 1682952543
transform 1 0 1992 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_103
timestamp 1682952543
transform 1 0 2000 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1682952543
transform -1 0 2112 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1682952543
transform 1 0 2112 0 -1 3570
box -8 -3 104 105
use FILL  FILL_348
timestamp 1682952543
transform 1 0 2208 0 -1 3570
box -8 -3 16 105
use FILL  FILL_349
timestamp 1682952543
transform 1 0 2216 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_97
timestamp 1682952543
transform 1 0 2224 0 -1 3570
box -8 -3 46 105
use M3_M2  M3_M2_1515
timestamp 1682952543
transform 1 0 2284 0 1 3475
box -3 -3 3 3
use OAI22X1  OAI22X1_98
timestamp 1682952543
transform 1 0 2264 0 -1 3570
box -8 -3 46 105
use FILL  FILL_350
timestamp 1682952543
transform 1 0 2304 0 -1 3570
box -8 -3 16 105
use FILL  FILL_351
timestamp 1682952543
transform 1 0 2312 0 -1 3570
box -8 -3 16 105
use FILL  FILL_352
timestamp 1682952543
transform 1 0 2320 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_99
timestamp 1682952543
transform 1 0 2328 0 -1 3570
box -8 -3 46 105
use FILL  FILL_353
timestamp 1682952543
transform 1 0 2368 0 -1 3570
box -8 -3 16 105
use FILL  FILL_354
timestamp 1682952543
transform 1 0 2376 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1682952543
transform 1 0 2384 0 -1 3570
box -8 -3 34 105
use M3_M2  M3_M2_1516
timestamp 1682952543
transform 1 0 2428 0 1 3475
box -3 -3 3 3
use FILL  FILL_355
timestamp 1682952543
transform 1 0 2416 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_100
timestamp 1682952543
transform -1 0 2464 0 -1 3570
box -8 -3 46 105
use FILL  FILL_356
timestamp 1682952543
transform 1 0 2464 0 -1 3570
box -8 -3 16 105
use FILL  FILL_357
timestamp 1682952543
transform 1 0 2472 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1682952543
transform 1 0 2480 0 -1 3570
box -8 -3 34 105
use FILL  FILL_358
timestamp 1682952543
transform 1 0 2512 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1517
timestamp 1682952543
transform 1 0 2532 0 1 3475
box -3 -3 3 3
use FILL  FILL_359
timestamp 1682952543
transform 1 0 2520 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_101
timestamp 1682952543
transform 1 0 2528 0 -1 3570
box -8 -3 46 105
use FILL  FILL_360
timestamp 1682952543
transform 1 0 2568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_361
timestamp 1682952543
transform 1 0 2576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_362
timestamp 1682952543
transform 1 0 2584 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1518
timestamp 1682952543
transform 1 0 2604 0 1 3475
box -3 -3 3 3
use FILL  FILL_363
timestamp 1682952543
transform 1 0 2592 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1519
timestamp 1682952543
transform 1 0 2628 0 1 3475
box -3 -3 3 3
use OAI21X1  OAI21X1_6
timestamp 1682952543
transform 1 0 2600 0 -1 3570
box -8 -3 34 105
use FILL  FILL_367
timestamp 1682952543
transform 1 0 2632 0 -1 3570
box -8 -3 16 105
use FILL  FILL_368
timestamp 1682952543
transform 1 0 2640 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1520
timestamp 1682952543
transform 1 0 2660 0 1 3475
box -3 -3 3 3
use FILL  FILL_369
timestamp 1682952543
transform 1 0 2648 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_103
timestamp 1682952543
transform 1 0 2656 0 -1 3570
box -8 -3 46 105
use FILL  FILL_376
timestamp 1682952543
transform 1 0 2696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_377
timestamp 1682952543
transform 1 0 2704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_378
timestamp 1682952543
transform 1 0 2712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_379
timestamp 1682952543
transform 1 0 2720 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1682952543
transform 1 0 2728 0 -1 3570
box -8 -3 34 105
use FILL  FILL_380
timestamp 1682952543
transform 1 0 2760 0 -1 3570
box -8 -3 16 105
use FILL  FILL_381
timestamp 1682952543
transform 1 0 2768 0 -1 3570
box -8 -3 16 105
use FILL  FILL_382
timestamp 1682952543
transform 1 0 2776 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1521
timestamp 1682952543
transform 1 0 2796 0 1 3475
box -3 -3 3 3
use OAI22X1  OAI22X1_104
timestamp 1682952543
transform 1 0 2784 0 -1 3570
box -8 -3 46 105
use FILL  FILL_383
timestamp 1682952543
transform 1 0 2824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_386
timestamp 1682952543
transform 1 0 2832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_387
timestamp 1682952543
transform 1 0 2840 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_105
timestamp 1682952543
transform -1 0 2888 0 -1 3570
box -8 -3 46 105
use FILL  FILL_388
timestamp 1682952543
transform 1 0 2888 0 -1 3570
box -8 -3 16 105
use FILL  FILL_389
timestamp 1682952543
transform 1 0 2896 0 -1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_2
timestamp 1682952543
transform 1 0 2904 0 -1 3570
box -8 -3 32 105
use FILL  FILL_392
timestamp 1682952543
transform 1 0 2928 0 -1 3570
box -8 -3 16 105
use FILL  FILL_393
timestamp 1682952543
transform 1 0 2936 0 -1 3570
box -8 -3 16 105
use FILL  FILL_394
timestamp 1682952543
transform 1 0 2944 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1522
timestamp 1682952543
transform 1 0 2980 0 1 3475
box -3 -3 3 3
use OAI22X1  OAI22X1_111
timestamp 1682952543
transform -1 0 2992 0 -1 3570
box -8 -3 46 105
use FILL  FILL_395
timestamp 1682952543
transform 1 0 2992 0 -1 3570
box -8 -3 16 105
use FILL  FILL_396
timestamp 1682952543
transform 1 0 3000 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1523
timestamp 1682952543
transform 1 0 3028 0 1 3475
box -3 -3 3 3
use NAND2X1  NAND2X1_3
timestamp 1682952543
transform 1 0 3008 0 -1 3570
box -8 -3 32 105
use FILL  FILL_397
timestamp 1682952543
transform 1 0 3032 0 -1 3570
box -8 -3 16 105
use FILL  FILL_398
timestamp 1682952543
transform 1 0 3040 0 -1 3570
box -8 -3 16 105
use FILL  FILL_399
timestamp 1682952543
transform 1 0 3048 0 -1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1682952543
transform 1 0 3056 0 -1 3570
box -8 -3 32 105
use FILL  FILL_400
timestamp 1682952543
transform 1 0 3080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_401
timestamp 1682952543
transform 1 0 3088 0 -1 3570
box -8 -3 16 105
use FILL  FILL_402
timestamp 1682952543
transform 1 0 3096 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_112
timestamp 1682952543
transform -1 0 3144 0 -1 3570
box -8 -3 46 105
use FILL  FILL_403
timestamp 1682952543
transform 1 0 3144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_404
timestamp 1682952543
transform 1 0 3152 0 -1 3570
box -8 -3 16 105
use FILL  FILL_405
timestamp 1682952543
transform 1 0 3160 0 -1 3570
box -8 -3 16 105
use FILL  FILL_406
timestamp 1682952543
transform 1 0 3168 0 -1 3570
box -8 -3 16 105
use FILL  FILL_407
timestamp 1682952543
transform 1 0 3176 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_105
timestamp 1682952543
transform 1 0 3184 0 -1 3570
box -9 -3 26 105
use OAI22X1  OAI22X1_116
timestamp 1682952543
transform 1 0 3200 0 -1 3570
box -8 -3 46 105
use OAI21X1  OAI21X1_13
timestamp 1682952543
transform 1 0 3240 0 -1 3570
box -8 -3 34 105
use OAI21X1  OAI21X1_14
timestamp 1682952543
transform 1 0 3272 0 -1 3570
box -8 -3 34 105
use FILL  FILL_411
timestamp 1682952543
transform 1 0 3304 0 -1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1682952543
transform -1 0 3336 0 -1 3570
box -8 -3 32 105
use FILL  FILL_412
timestamp 1682952543
transform 1 0 3336 0 -1 3570
box -8 -3 16 105
use FILL  FILL_413
timestamp 1682952543
transform 1 0 3344 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_15
timestamp 1682952543
transform -1 0 3384 0 -1 3570
box -8 -3 34 105
use FILL  FILL_414
timestamp 1682952543
transform 1 0 3384 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_1524
timestamp 1682952543
transform 1 0 3436 0 1 3475
box -3 -3 3 3
use OAI22X1  OAI22X1_117
timestamp 1682952543
transform 1 0 3392 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_118
timestamp 1682952543
transform 1 0 3432 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_119
timestamp 1682952543
transform 1 0 3472 0 -1 3570
box -8 -3 46 105
use INVX2  INVX2_110
timestamp 1682952543
transform -1 0 3528 0 -1 3570
box -9 -3 26 105
use FILL  FILL_415
timestamp 1682952543
transform 1 0 3528 0 -1 3570
box -8 -3 16 105
use FILL  FILL_416
timestamp 1682952543
transform 1 0 3536 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_16
timestamp 1682952543
transform 1 0 3544 0 -1 3570
box -8 -3 34 105
use FILL  FILL_417
timestamp 1682952543
transform 1 0 3576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_418
timestamp 1682952543
transform 1 0 3584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_419
timestamp 1682952543
transform 1 0 3592 0 -1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_6
timestamp 1682952543
transform 1 0 3600 0 -1 3570
box -8 -3 32 105
use FILL  FILL_420
timestamp 1682952543
transform 1 0 3624 0 -1 3570
box -8 -3 16 105
use FILL  FILL_421
timestamp 1682952543
transform 1 0 3632 0 -1 3570
box -8 -3 16 105
use FILL  FILL_422
timestamp 1682952543
transform 1 0 3640 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_17
timestamp 1682952543
transform -1 0 3680 0 -1 3570
box -8 -3 34 105
use FILL  FILL_423
timestamp 1682952543
transform 1 0 3680 0 -1 3570
box -8 -3 16 105
use FILL  FILL_424
timestamp 1682952543
transform 1 0 3688 0 -1 3570
box -8 -3 16 105
use FILL  FILL_431
timestamp 1682952543
transform 1 0 3696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_432
timestamp 1682952543
transform 1 0 3704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_433
timestamp 1682952543
transform 1 0 3712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_434
timestamp 1682952543
transform 1 0 3720 0 -1 3570
box -8 -3 16 105
use FILL  FILL_435
timestamp 1682952543
transform 1 0 3728 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_122
timestamp 1682952543
transform 1 0 3736 0 -1 3570
box -8 -3 46 105
use FILL  FILL_436
timestamp 1682952543
transform 1 0 3776 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_18
timestamp 1682952543
transform 1 0 3784 0 -1 3570
box -8 -3 34 105
use FILL  FILL_437
timestamp 1682952543
transform 1 0 3816 0 -1 3570
box -8 -3 16 105
use FILL  FILL_441
timestamp 1682952543
transform 1 0 3824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_442
timestamp 1682952543
transform 1 0 3832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_443
timestamp 1682952543
transform 1 0 3840 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_20
timestamp 1682952543
transform -1 0 3880 0 -1 3570
box -8 -3 34 105
use FILL  FILL_444
timestamp 1682952543
transform 1 0 3880 0 -1 3570
box -8 -3 16 105
use FILL  FILL_445
timestamp 1682952543
transform 1 0 3888 0 -1 3570
box -8 -3 16 105
use FILL  FILL_446
timestamp 1682952543
transform 1 0 3896 0 -1 3570
box -8 -3 16 105
use FILL  FILL_447
timestamp 1682952543
transform 1 0 3904 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_23
timestamp 1682952543
transform -1 0 3944 0 -1 3570
box -8 -3 34 105
use OAI22X1  OAI22X1_124
timestamp 1682952543
transform 1 0 3944 0 -1 3570
box -8 -3 46 105
use OAI22X1  OAI22X1_125
timestamp 1682952543
transform 1 0 3984 0 -1 3570
box -8 -3 46 105
use INVX2  INVX2_111
timestamp 1682952543
transform -1 0 4040 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1682952543
transform 1 0 4040 0 -1 3570
box -8 -3 104 105
use FILL  FILL_448
timestamp 1682952543
transform 1 0 4136 0 -1 3570
box -8 -3 16 105
use FILL  FILL_449
timestamp 1682952543
transform 1 0 4144 0 -1 3570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_13
timestamp 1682952543
transform 1 0 4201 0 1 3470
box -10 -3 10 3
use M2_M1  M2_M1_1597
timestamp 1682952543
transform 1 0 116 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1750
timestamp 1682952543
transform 1 0 124 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1682952543
transform 1 0 140 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1682952543
transform 1 0 148 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1598
timestamp 1682952543
transform 1 0 140 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1727
timestamp 1682952543
transform 1 0 148 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1587
timestamp 1682952543
transform 1 0 268 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1613
timestamp 1682952543
transform 1 0 172 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1614
timestamp 1682952543
transform 1 0 188 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1615
timestamp 1682952543
transform 1 0 228 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1557
timestamp 1682952543
transform 1 0 300 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1588
timestamp 1682952543
transform 1 0 300 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1599
timestamp 1682952543
transform 1 0 172 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1682952543
transform 1 0 188 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1682952543
transform 1 0 228 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1602
timestamp 1682952543
transform 1 0 284 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1654
timestamp 1682952543
transform 1 0 292 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1603
timestamp 1682952543
transform 1 0 300 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1682952543
transform 1 0 164 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1682952543
transform 1 0 188 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1730
timestamp 1682952543
transform 1 0 204 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1731
timestamp 1682952543
transform 1 0 292 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1712
timestamp 1682952543
transform 1 0 164 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1682952543
transform 1 0 180 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1694
timestamp 1682952543
transform 1 0 300 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1682952543
transform 1 0 316 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1682952543
transform 1 0 340 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1682952543
transform 1 0 356 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1682952543
transform 1 0 332 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1682952543
transform 1 0 396 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1616
timestamp 1682952543
transform 1 0 388 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1617
timestamp 1682952543
transform 1 0 492 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1604
timestamp 1682952543
transform 1 0 324 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1682952543
transform 1 0 340 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1682952543
transform 1 0 356 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1682952543
transform 1 0 364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1682952543
transform 1 0 380 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1609
timestamp 1682952543
transform 1 0 396 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1682952543
transform 1 0 308 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1752
timestamp 1682952543
transform 1 0 236 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1753
timestamp 1682952543
transform 1 0 292 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1682952543
transform 1 0 308 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1695
timestamp 1682952543
transform 1 0 340 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1733
timestamp 1682952543
transform 1 0 364 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1682952543
transform 1 0 372 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1682952543
transform 1 0 388 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1755
timestamp 1682952543
transform 1 0 372 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1682952543
transform 1 0 412 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1682952543
transform 1 0 564 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1590
timestamp 1682952543
transform 1 0 532 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1610
timestamp 1682952543
transform 1 0 436 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1611
timestamp 1682952543
transform 1 0 492 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1682952543
transform 1 0 508 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1613
timestamp 1682952543
transform 1 0 524 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1614
timestamp 1682952543
transform 1 0 532 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1657
timestamp 1682952543
transform 1 0 548 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1615
timestamp 1682952543
transform 1 0 556 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1658
timestamp 1682952543
transform 1 0 580 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1616
timestamp 1682952543
transform 1 0 588 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1682952543
transform 1 0 412 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1737
timestamp 1682952543
transform 1 0 500 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1682952543
transform 1 0 516 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1739
timestamp 1682952543
transform 1 0 532 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1682952543
transform 1 0 548 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1741
timestamp 1682952543
transform 1 0 564 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1742
timestamp 1682952543
transform 1 0 572 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1682952543
transform 1 0 580 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1713
timestamp 1682952543
transform 1 0 500 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1714
timestamp 1682952543
transform 1 0 524 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1682952543
transform 1 0 524 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1682952543
transform 1 0 540 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1659
timestamp 1682952543
transform 1 0 596 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1682952543
transform 1 0 612 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1682952543
transform 1 0 708 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1682952543
transform 1 0 644 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1619
timestamp 1682952543
transform 1 0 748 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1682952543
transform 1 0 764 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1682952543
transform 1 0 796 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1591
timestamp 1682952543
transform 1 0 796 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1617
timestamp 1682952543
transform 1 0 668 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1682952543
transform 1 0 700 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1619
timestamp 1682952543
transform 1 0 716 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1620
timestamp 1682952543
transform 1 0 732 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1660
timestamp 1682952543
transform 1 0 740 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1621
timestamp 1682952543
transform 1 0 748 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1661
timestamp 1682952543
transform 1 0 756 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1622
timestamp 1682952543
transform 1 0 764 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1662
timestamp 1682952543
transform 1 0 772 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1623
timestamp 1682952543
transform 1 0 780 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1682952543
transform 1 0 796 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1682952543
transform 1 0 804 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1682952543
transform 1 0 620 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1682952543
transform 1 0 708 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1682952543
transform 1 0 724 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1747
timestamp 1682952543
transform 1 0 740 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1715
timestamp 1682952543
transform 1 0 636 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1682952543
transform 1 0 716 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1682952543
transform 1 0 724 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1748
timestamp 1682952543
transform 1 0 764 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1682952543
transform 1 0 772 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1541
timestamp 1682952543
transform 1 0 820 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1682952543
transform 1 0 844 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1682952543
transform 1 0 852 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1626
timestamp 1682952543
transform 1 0 836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1627
timestamp 1682952543
transform 1 0 852 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1682952543
transform 1 0 828 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1751
timestamp 1682952543
transform 1 0 844 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1682952543
transform 1 0 852 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1564
timestamp 1682952543
transform 1 0 876 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1542
timestamp 1682952543
transform 1 0 972 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1682952543
transform 1 0 964 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1682952543
transform 1 0 868 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1623
timestamp 1682952543
transform 1 0 916 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1628
timestamp 1682952543
transform 1 0 868 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1682952543
transform 1 0 876 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1682952543
transform 1 0 916 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1696
timestamp 1682952543
transform 1 0 876 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1697
timestamp 1682952543
transform 1 0 932 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1753
timestamp 1682952543
transform 1 0 956 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1663
timestamp 1682952543
transform 1 0 980 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1754
timestamp 1682952543
transform 1 0 980 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1682952543
transform 1 0 972 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_1848
timestamp 1682952543
transform 1 0 988 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_1543
timestamp 1682952543
transform 1 0 1004 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1682952543
transform 1 0 1052 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1624
timestamp 1682952543
transform 1 0 1068 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1631
timestamp 1682952543
transform 1 0 1068 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1592
timestamp 1682952543
transform 1 0 1092 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1682952543
transform 1 0 1092 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1755
timestamp 1682952543
transform 1 0 1100 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1682952543
transform 1 0 1092 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_1759
timestamp 1682952543
transform 1 0 1092 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1756
timestamp 1682952543
transform 1 0 1116 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1682952543
transform 1 0 1124 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1633
timestamp 1682952543
transform 1 0 1132 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1526
timestamp 1682952543
transform 1 0 1156 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_1634
timestamp 1682952543
transform 1 0 1148 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1635
timestamp 1682952543
transform 1 0 1156 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1698
timestamp 1682952543
transform 1 0 1140 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1717
timestamp 1682952543
transform 1 0 1132 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1527
timestamp 1682952543
transform 1 0 1204 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1544
timestamp 1682952543
transform 1 0 1252 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1625
timestamp 1682952543
transform 1 0 1212 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1682952543
transform 1 0 1276 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_1636
timestamp 1682952543
transform 1 0 1172 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1637
timestamp 1682952543
transform 1 0 1220 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1665
timestamp 1682952543
transform 1 0 1268 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1638
timestamp 1682952543
transform 1 0 1276 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1758
timestamp 1682952543
transform 1 0 1252 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1682952543
transform 1 0 1268 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1682952543
transform 1 0 1284 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1718
timestamp 1682952543
transform 1 0 1284 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1682952543
transform 1 0 1308 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1567
timestamp 1682952543
transform 1 0 1348 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_1639
timestamp 1682952543
transform 1 0 1332 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1666
timestamp 1682952543
transform 1 0 1340 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1528
timestamp 1682952543
transform 1 0 1492 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1529
timestamp 1682952543
transform 1 0 1508 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1682952543
transform 1 0 1388 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1569
timestamp 1682952543
transform 1 0 1468 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1570
timestamp 1682952543
transform 1 0 1484 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1682952543
transform 1 0 1444 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1627
timestamp 1682952543
transform 1 0 1484 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1640
timestamp 1682952543
transform 1 0 1348 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1682952543
transform 1 0 1364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1642
timestamp 1682952543
transform 1 0 1380 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1682952543
transform 1 0 1444 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1644
timestamp 1682952543
transform 1 0 1476 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1645
timestamp 1682952543
transform 1 0 1484 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1646
timestamp 1682952543
transform 1 0 1500 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1699
timestamp 1682952543
transform 1 0 1332 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1850
timestamp 1682952543
transform 1 0 1340 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_1761
timestamp 1682952543
transform 1 0 1372 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1762
timestamp 1682952543
transform 1 0 1396 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1667
timestamp 1682952543
transform 1 0 1508 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1647
timestamp 1682952543
transform 1 0 1516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1682952543
transform 1 0 1500 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1682952543
transform 1 0 1508 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1682952543
transform 1 0 1524 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1719
timestamp 1682952543
transform 1 0 1396 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1720
timestamp 1682952543
transform 1 0 1420 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1682952543
transform 1 0 1476 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1682952543
transform 1 0 1524 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1648
timestamp 1682952543
transform 1 0 1540 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1628
timestamp 1682952543
transform 1 0 1548 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1700
timestamp 1682952543
transform 1 0 1540 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1546
timestamp 1682952543
transform 1 0 1580 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1593
timestamp 1682952543
transform 1 0 1572 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1629
timestamp 1682952543
transform 1 0 1596 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1649
timestamp 1682952543
transform 1 0 1580 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1682952543
transform 1 0 1596 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1682952543
transform 1 0 1548 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1767
timestamp 1682952543
transform 1 0 1556 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1682952543
transform 1 0 1572 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1682952543
transform 1 0 1588 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1682952543
transform 1 0 1596 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1723
timestamp 1682952543
transform 1 0 1588 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1668
timestamp 1682952543
transform 1 0 1604 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1682952543
transform 1 0 1652 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1682952543
transform 1 0 1636 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1631
timestamp 1682952543
transform 1 0 1660 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1651
timestamp 1682952543
transform 1 0 1612 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1652
timestamp 1682952543
transform 1 0 1620 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1682952543
transform 1 0 1636 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1654
timestamp 1682952543
transform 1 0 1652 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1682952543
transform 1 0 1612 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1760
timestamp 1682952543
transform 1 0 1620 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1772
timestamp 1682952543
transform 1 0 1652 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1682952543
transform 1 0 1660 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1724
timestamp 1682952543
transform 1 0 1652 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1632
timestamp 1682952543
transform 1 0 1684 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1633
timestamp 1682952543
transform 1 0 1724 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1634
timestamp 1682952543
transform 1 0 1748 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1655
timestamp 1682952543
transform 1 0 1684 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1656
timestamp 1682952543
transform 1 0 1692 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1657
timestamp 1682952543
transform 1 0 1724 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1682952543
transform 1 0 1772 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1725
timestamp 1682952543
transform 1 0 1700 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1682952543
transform 1 0 1788 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1658
timestamp 1682952543
transform 1 0 1788 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1530
timestamp 1682952543
transform 1 0 1812 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1531
timestamp 1682952543
transform 1 0 1868 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1682952543
transform 1 0 1804 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1659
timestamp 1682952543
transform 1 0 1836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1682952543
transform 1 0 1876 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1726
timestamp 1682952543
transform 1 0 1876 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1682952543
transform 1 0 1804 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1670
timestamp 1682952543
transform 1 0 1892 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1776
timestamp 1682952543
transform 1 0 1892 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1636
timestamp 1682952543
transform 1 0 2004 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1660
timestamp 1682952543
transform 1 0 1924 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1661
timestamp 1682952543
transform 1 0 1980 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1682952543
transform 1 0 2020 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1682952543
transform 1 0 1940 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1727
timestamp 1682952543
transform 1 0 1940 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1637
timestamp 1682952543
transform 1 0 2036 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1663
timestamp 1682952543
transform 1 0 2036 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1682952543
transform 1 0 2076 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1665
timestamp 1682952543
transform 1 0 2132 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1666
timestamp 1682952543
transform 1 0 2140 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1778
timestamp 1682952543
transform 1 0 2116 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1547
timestamp 1682952543
transform 1 0 2156 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_1779
timestamp 1682952543
transform 1 0 2156 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1638
timestamp 1682952543
transform 1 0 2220 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1682952543
transform 1 0 2212 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1667
timestamp 1682952543
transform 1 0 2220 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1682952543
transform 1 0 2204 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1781
timestamp 1682952543
transform 1 0 2236 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1639
timestamp 1682952543
transform 1 0 2252 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1782
timestamp 1682952543
transform 1 0 2252 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1682952543
transform 1 0 2260 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1701
timestamp 1682952543
transform 1 0 2268 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1682952543
transform 1 0 2292 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1640
timestamp 1682952543
transform 1 0 2316 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1669
timestamp 1682952543
transform 1 0 2284 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1672
timestamp 1682952543
transform 1 0 2292 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1670
timestamp 1682952543
transform 1 0 2300 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1673
timestamp 1682952543
transform 1 0 2308 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1671
timestamp 1682952543
transform 1 0 2316 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1783
timestamp 1682952543
transform 1 0 2308 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1702
timestamp 1682952543
transform 1 0 2316 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1682952543
transform 1 0 2308 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1672
timestamp 1682952543
transform 1 0 2332 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1571
timestamp 1682952543
transform 1 0 2364 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1641
timestamp 1682952543
transform 1 0 2380 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1682952543
transform 1 0 2356 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1673
timestamp 1682952543
transform 1 0 2364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1682952543
transform 1 0 2380 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1682952543
transform 1 0 2348 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1595
timestamp 1682952543
transform 1 0 2396 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1785
timestamp 1682952543
transform 1 0 2372 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1682952543
transform 1 0 2388 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1682952543
transform 1 0 2396 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1728
timestamp 1682952543
transform 1 0 2372 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1763
timestamp 1682952543
transform 1 0 2396 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1682952543
transform 1 0 2412 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1572
timestamp 1682952543
transform 1 0 2452 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1597
timestamp 1682952543
transform 1 0 2436 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1580
timestamp 1682952543
transform 1 0 2436 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1675
timestamp 1682952543
transform 1 0 2420 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1675
timestamp 1682952543
transform 1 0 2436 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1581
timestamp 1682952543
transform 1 0 2468 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1676
timestamp 1682952543
transform 1 0 2444 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1703
timestamp 1682952543
transform 1 0 2428 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1676
timestamp 1682952543
transform 1 0 2468 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1533
timestamp 1682952543
transform 1 0 2516 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1573
timestamp 1682952543
transform 1 0 2508 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1598
timestamp 1682952543
transform 1 0 2492 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1599
timestamp 1682952543
transform 1 0 2524 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1582
timestamp 1682952543
transform 1 0 2492 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_1642
timestamp 1682952543
transform 1 0 2500 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1583
timestamp 1682952543
transform 1 0 2524 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1682952543
transform 1 0 2492 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1677
timestamp 1682952543
transform 1 0 2508 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1788
timestamp 1682952543
transform 1 0 2436 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1682952543
transform 1 0 2444 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1682952543
transform 1 0 2468 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1682952543
transform 1 0 2476 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1682952543
transform 1 0 2492 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1729
timestamp 1682952543
transform 1 0 2444 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1682952543
transform 1 0 2468 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1793
timestamp 1682952543
transform 1 0 2524 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1678
timestamp 1682952543
transform 1 0 2532 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1682952543
transform 1 0 2532 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1730
timestamp 1682952543
transform 1 0 2524 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1643
timestamp 1682952543
transform 1 0 2564 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1678
timestamp 1682952543
transform 1 0 2556 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1795
timestamp 1682952543
transform 1 0 2556 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1796
timestamp 1682952543
transform 1 0 2564 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1731
timestamp 1682952543
transform 1 0 2556 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1584
timestamp 1682952543
transform 1 0 2580 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_1534
timestamp 1682952543
transform 1 0 2612 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_1679
timestamp 1682952543
transform 1 0 2588 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1732
timestamp 1682952543
transform 1 0 2580 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1679
timestamp 1682952543
transform 1 0 2596 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1797
timestamp 1682952543
transform 1 0 2596 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1574
timestamp 1682952543
transform 1 0 2620 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1600
timestamp 1682952543
transform 1 0 2620 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1585
timestamp 1682952543
transform 1 0 2620 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1682952543
transform 1 0 2628 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1681
timestamp 1682952543
transform 1 0 2636 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1682952543
transform 1 0 2628 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1733
timestamp 1682952543
transform 1 0 2620 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1575
timestamp 1682952543
transform 1 0 2652 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1601
timestamp 1682952543
transform 1 0 2652 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1586
timestamp 1682952543
transform 1 0 2660 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1682952543
transform 1 0 2668 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_1734
timestamp 1682952543
transform 1 0 2668 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1680
timestamp 1682952543
transform 1 0 2700 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1682952543
transform 1 0 2724 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_1602
timestamp 1682952543
transform 1 0 2724 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1588
timestamp 1682952543
transform 1 0 2724 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1682952543
transform 1 0 2708 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1682952543
transform 1 0 2692 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1682952543
transform 1 0 2700 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1681
timestamp 1682952543
transform 1 0 2724 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1682952543
transform 1 0 2708 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1683
timestamp 1682952543
transform 1 0 2748 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1682952543
transform 1 0 2740 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1736
timestamp 1682952543
transform 1 0 2732 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1765
timestamp 1682952543
transform 1 0 2740 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1682952543
transform 1 0 2772 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_1589
timestamp 1682952543
transform 1 0 2764 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1684
timestamp 1682952543
transform 1 0 2764 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1685
timestamp 1682952543
transform 1 0 2772 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1548
timestamp 1682952543
transform 1 0 2828 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1549
timestamp 1682952543
transform 1 0 2884 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1682952543
transform 1 0 2820 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1603
timestamp 1682952543
transform 1 0 2804 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1686
timestamp 1682952543
transform 1 0 2836 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1682
timestamp 1682952543
transform 1 0 2860 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1802
timestamp 1682952543
transform 1 0 2884 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1550
timestamp 1682952543
transform 1 0 2916 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_1687
timestamp 1682952543
transform 1 0 2916 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1578
timestamp 1682952543
transform 1 0 2940 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1644
timestamp 1682952543
transform 1 0 2948 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1683
timestamp 1682952543
transform 1 0 2940 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1688
timestamp 1682952543
transform 1 0 2948 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1682952543
transform 1 0 2964 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1682952543
transform 1 0 2924 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1682952543
transform 1 0 2940 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1682952543
transform 1 0 2956 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1682952543
transform 1 0 2964 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1682952543
transform 1 0 2988 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1690
timestamp 1682952543
transform 1 0 2988 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1737
timestamp 1682952543
transform 1 0 2940 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1738
timestamp 1682952543
transform 1 0 2964 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1766
timestamp 1682952543
transform 1 0 2924 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1682952543
transform 1 0 2988 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1682952543
transform 1 0 3004 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1807
timestamp 1682952543
transform 1 0 3004 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1604
timestamp 1682952543
transform 1 0 3028 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_1591
timestamp 1682952543
transform 1 0 3052 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_1685
timestamp 1682952543
transform 1 0 3052 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1691
timestamp 1682952543
transform 1 0 3060 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1808
timestamp 1682952543
transform 1 0 3028 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1682952543
transform 1 0 3036 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1704
timestamp 1682952543
transform 1 0 3044 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1810
timestamp 1682952543
transform 1 0 3052 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1579
timestamp 1682952543
transform 1 0 3108 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1605
timestamp 1682952543
transform 1 0 3100 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1645
timestamp 1682952543
transform 1 0 3092 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1692
timestamp 1682952543
transform 1 0 3100 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1768
timestamp 1682952543
transform 1 0 3100 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1592
timestamp 1682952543
transform 1 0 3116 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_1551
timestamp 1682952543
transform 1 0 3132 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1682952543
transform 1 0 3124 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1693
timestamp 1682952543
transform 1 0 3156 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1687
timestamp 1682952543
transform 1 0 3164 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1811
timestamp 1682952543
transform 1 0 3164 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1552
timestamp 1682952543
transform 1 0 3212 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1682952543
transform 1 0 3228 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_1694
timestamp 1682952543
transform 1 0 3204 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1682952543
transform 1 0 3212 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1696
timestamp 1682952543
transform 1 0 3228 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1682952543
transform 1 0 3188 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1682952543
transform 1 0 3204 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1705
timestamp 1682952543
transform 1 0 3212 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1814
timestamp 1682952543
transform 1 0 3220 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1682952543
transform 1 0 3236 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1581
timestamp 1682952543
transform 1 0 3268 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_1697
timestamp 1682952543
transform 1 0 3268 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1593
timestamp 1682952543
transform 1 0 3292 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1698
timestamp 1682952543
transform 1 0 3284 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1682952543
transform 1 0 3292 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1706
timestamp 1682952543
transform 1 0 3308 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1594
timestamp 1682952543
transform 1 0 3332 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1699
timestamp 1682952543
transform 1 0 3364 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1536
timestamp 1682952543
transform 1 0 3404 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_1700
timestamp 1682952543
transform 1 0 3396 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1817
timestamp 1682952543
transform 1 0 3396 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1739
timestamp 1682952543
transform 1 0 3396 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1553
timestamp 1682952543
transform 1 0 3412 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1682952543
transform 1 0 3420 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_1701
timestamp 1682952543
transform 1 0 3412 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1682952543
transform 1 0 3428 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1707
timestamp 1682952543
transform 1 0 3412 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1818
timestamp 1682952543
transform 1 0 3420 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1682952543
transform 1 0 3436 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1740
timestamp 1682952543
transform 1 0 3420 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1820
timestamp 1682952543
transform 1 0 3468 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1537
timestamp 1682952543
transform 1 0 3484 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_1703
timestamp 1682952543
transform 1 0 3476 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1646
timestamp 1682952543
transform 1 0 3500 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1704
timestamp 1682952543
transform 1 0 3500 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1682952543
transform 1 0 3500 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1741
timestamp 1682952543
transform 1 0 3492 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1822
timestamp 1682952543
transform 1 0 3508 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1742
timestamp 1682952543
transform 1 0 3508 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1705
timestamp 1682952543
transform 1 0 3532 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1688
timestamp 1682952543
transform 1 0 3540 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1682952543
transform 1 0 3580 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1682952543
transform 1 0 3596 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_1706
timestamp 1682952543
transform 1 0 3548 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1682952543
transform 1 0 3564 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1708
timestamp 1682952543
transform 1 0 3580 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1682952543
transform 1 0 3596 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1823
timestamp 1682952543
transform 1 0 3540 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1708
timestamp 1682952543
transform 1 0 3564 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1824
timestamp 1682952543
transform 1 0 3572 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1825
timestamp 1682952543
transform 1 0 3588 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1826
timestamp 1682952543
transform 1 0 3604 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1682952543
transform 1 0 3612 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1743
timestamp 1682952543
transform 1 0 3548 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1682952543
transform 1 0 3588 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1682952543
transform 1 0 3572 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1682952543
transform 1 0 3644 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_1710
timestamp 1682952543
transform 1 0 3628 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1682952543
transform 1 0 3644 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1745
timestamp 1682952543
transform 1 0 3612 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1828
timestamp 1682952543
transform 1 0 3644 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1770
timestamp 1682952543
transform 1 0 3628 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1595
timestamp 1682952543
transform 1 0 3652 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_1606
timestamp 1682952543
transform 1 0 3676 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1682952543
transform 1 0 3700 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1682952543
transform 1 0 3692 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1682952543
transform 1 0 3716 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1682952543
transform 1 0 3716 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1712
timestamp 1682952543
transform 1 0 3692 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1682952543
transform 1 0 3716 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1829
timestamp 1682952543
transform 1 0 3684 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1689
timestamp 1682952543
transform 1 0 3724 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1830
timestamp 1682952543
transform 1 0 3708 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1831
timestamp 1682952543
transform 1 0 3724 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1832
timestamp 1682952543
transform 1 0 3732 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1556
timestamp 1682952543
transform 1 0 3748 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1682952543
transform 1 0 3740 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1682952543
transform 1 0 3732 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_1714
timestamp 1682952543
transform 1 0 3748 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1585
timestamp 1682952543
transform 1 0 3764 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1586
timestamp 1682952543
transform 1 0 3780 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_1690
timestamp 1682952543
transform 1 0 3764 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1715
timestamp 1682952543
transform 1 0 3780 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1682952543
transform 1 0 3772 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1709
timestamp 1682952543
transform 1 0 3780 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_1609
timestamp 1682952543
transform 1 0 3812 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1682952543
transform 1 0 3804 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1682952543
transform 1 0 3796 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1834
timestamp 1682952543
transform 1 0 3788 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1835
timestamp 1682952543
transform 1 0 3796 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1747
timestamp 1682952543
transform 1 0 3796 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1682952543
transform 1 0 3836 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1716
timestamp 1682952543
transform 1 0 3812 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1682952543
transform 1 0 3836 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1682952543
transform 1 0 3828 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1682952543
transform 1 0 3844 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1838
timestamp 1682952543
transform 1 0 3860 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1682952543
transform 1 0 3876 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1710
timestamp 1682952543
transform 1 0 3884 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1596
timestamp 1682952543
transform 1 0 3916 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1682952543
transform 1 0 3932 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1771
timestamp 1682952543
transform 1 0 3916 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_1720
timestamp 1682952543
transform 1 0 3948 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1839
timestamp 1682952543
transform 1 0 3956 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1610
timestamp 1682952543
transform 1 0 3972 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1611
timestamp 1682952543
transform 1 0 3988 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_1650
timestamp 1682952543
transform 1 0 3988 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1721
timestamp 1682952543
transform 1 0 3972 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1722
timestamp 1682952543
transform 1 0 3988 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1840
timestamp 1682952543
transform 1 0 3980 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1841
timestamp 1682952543
transform 1 0 3996 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1651
timestamp 1682952543
transform 1 0 4012 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1842
timestamp 1682952543
transform 1 0 4012 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1652
timestamp 1682952543
transform 1 0 4036 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1723
timestamp 1682952543
transform 1 0 4036 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1724
timestamp 1682952543
transform 1 0 4052 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1692
timestamp 1682952543
transform 1 0 4060 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1725
timestamp 1682952543
transform 1 0 4068 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1682952543
transform 1 0 4044 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1711
timestamp 1682952543
transform 1 0 4052 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_1844
timestamp 1682952543
transform 1 0 4060 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_1653
timestamp 1682952543
transform 1 0 4084 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_1726
timestamp 1682952543
transform 1 0 4084 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_1748
timestamp 1682952543
transform 1 0 4060 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1682952543
transform 1 0 4076 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_1693
timestamp 1682952543
transform 1 0 4100 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_1845
timestamp 1682952543
transform 1 0 4092 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1682952543
transform 1 0 4132 0 1 3405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_14
timestamp 1682952543
transform 1 0 48 0 1 3370
box -10 -3 10 3
use FILL  FILL_450
timestamp 1682952543
transform 1 0 72 0 1 3370
box -8 -3 16 105
use FILL  FILL_451
timestamp 1682952543
transform 1 0 80 0 1 3370
box -8 -3 16 105
use FILL  FILL_452
timestamp 1682952543
transform 1 0 88 0 1 3370
box -8 -3 16 105
use FILL  FILL_453
timestamp 1682952543
transform 1 0 96 0 1 3370
box -8 -3 16 105
use FILL  FILL_454
timestamp 1682952543
transform 1 0 104 0 1 3370
box -8 -3 16 105
use FILL  FILL_455
timestamp 1682952543
transform 1 0 112 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_112
timestamp 1682952543
transform -1 0 136 0 1 3370
box -9 -3 26 105
use FILL  FILL_456
timestamp 1682952543
transform 1 0 136 0 1 3370
box -8 -3 16 105
use FILL  FILL_457
timestamp 1682952543
transform 1 0 144 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1772
timestamp 1682952543
transform 1 0 188 0 1 3375
box -3 -3 3 3
use AOI22X1  AOI22X1_53
timestamp 1682952543
transform -1 0 192 0 1 3370
box -8 -3 46 105
use M3_M2  M3_M2_1773
timestamp 1682952543
transform 1 0 212 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1682952543
transform 1 0 252 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_109
timestamp 1682952543
transform 1 0 192 0 1 3370
box -8 -3 104 105
use INVX2  INVX2_113
timestamp 1682952543
transform 1 0 288 0 1 3370
box -9 -3 26 105
use FILL  FILL_458
timestamp 1682952543
transform 1 0 304 0 1 3370
box -8 -3 16 105
use FILL  FILL_459
timestamp 1682952543
transform 1 0 312 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1775
timestamp 1682952543
transform 1 0 380 0 1 3375
box -3 -3 3 3
use AOI22X1  AOI22X1_54
timestamp 1682952543
transform 1 0 320 0 1 3370
box -8 -3 46 105
use M3_M2  M3_M2_1776
timestamp 1682952543
transform 1 0 412 0 1 3375
box -3 -3 3 3
use AOI22X1  AOI22X1_55
timestamp 1682952543
transform 1 0 360 0 1 3370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1682952543
transform 1 0 400 0 1 3370
box -8 -3 104 105
use M3_M2  M3_M2_1777
timestamp 1682952543
transform 1 0 516 0 1 3375
box -3 -3 3 3
use OAI22X1  OAI22X1_126
timestamp 1682952543
transform -1 0 536 0 1 3370
box -8 -3 46 105
use AOI22X1  AOI22X1_56
timestamp 1682952543
transform 1 0 536 0 1 3370
box -8 -3 46 105
use INVX2  INVX2_114
timestamp 1682952543
transform 1 0 576 0 1 3370
box -9 -3 26 105
use FILL  FILL_460
timestamp 1682952543
transform 1 0 592 0 1 3370
box -8 -3 16 105
use FILL  FILL_464
timestamp 1682952543
transform 1 0 600 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1682952543
transform 1 0 608 0 1 3370
box -8 -3 104 105
use OAI22X1  OAI22X1_128
timestamp 1682952543
transform 1 0 704 0 1 3370
box -8 -3 46 105
use INVX2  INVX2_121
timestamp 1682952543
transform -1 0 760 0 1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_59
timestamp 1682952543
transform -1 0 800 0 1 3370
box -8 -3 46 105
use FILL  FILL_466
timestamp 1682952543
transform 1 0 800 0 1 3370
box -8 -3 16 105
use FILL  FILL_469
timestamp 1682952543
transform 1 0 808 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_60
timestamp 1682952543
transform 1 0 816 0 1 3370
box -8 -3 46 105
use INVX2  INVX2_122
timestamp 1682952543
transform 1 0 856 0 1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_116
timestamp 1682952543
transform -1 0 968 0 1 3370
box -8 -3 104 105
use M3_M2  M3_M2_1778
timestamp 1682952543
transform 1 0 988 0 1 3375
box -3 -3 3 3
use NOR2X1  NOR2X1_13
timestamp 1682952543
transform 1 0 968 0 1 3370
box -8 -3 32 105
use FILL  FILL_471
timestamp 1682952543
transform 1 0 992 0 1 3370
box -8 -3 16 105
use FILL  FILL_472
timestamp 1682952543
transform 1 0 1000 0 1 3370
box -8 -3 16 105
use FILL  FILL_473
timestamp 1682952543
transform 1 0 1008 0 1 3370
box -8 -3 16 105
use FILL  FILL_474
timestamp 1682952543
transform 1 0 1016 0 1 3370
box -8 -3 16 105
use FILL  FILL_475
timestamp 1682952543
transform 1 0 1024 0 1 3370
box -8 -3 16 105
use FILL  FILL_476
timestamp 1682952543
transform 1 0 1032 0 1 3370
box -8 -3 16 105
use FILL  FILL_477
timestamp 1682952543
transform 1 0 1040 0 1 3370
box -8 -3 16 105
use FILL  FILL_478
timestamp 1682952543
transform 1 0 1048 0 1 3370
box -8 -3 16 105
use FILL  FILL_479
timestamp 1682952543
transform 1 0 1056 0 1 3370
box -8 -3 16 105
use FILL  FILL_480
timestamp 1682952543
transform 1 0 1064 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1682952543
transform 1 0 1072 0 1 3370
box -8 -3 32 105
use NOR2X1  NOR2X1_15
timestamp 1682952543
transform 1 0 1096 0 1 3370
box -8 -3 32 105
use FILL  FILL_481
timestamp 1682952543
transform 1 0 1120 0 1 3370
box -8 -3 16 105
use FILL  FILL_482
timestamp 1682952543
transform 1 0 1128 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_123
timestamp 1682952543
transform 1 0 1136 0 1 3370
box -9 -3 26 105
use FILL  FILL_483
timestamp 1682952543
transform 1 0 1152 0 1 3370
box -8 -3 16 105
use FILL  FILL_491
timestamp 1682952543
transform 1 0 1160 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1682952543
transform -1 0 1264 0 1 3370
box -8 -3 104 105
use OAI22X1  OAI22X1_130
timestamp 1682952543
transform -1 0 1304 0 1 3370
box -8 -3 46 105
use FILL  FILL_492
timestamp 1682952543
transform 1 0 1304 0 1 3370
box -8 -3 16 105
use FILL  FILL_493
timestamp 1682952543
transform 1 0 1312 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1779
timestamp 1682952543
transform 1 0 1332 0 1 3375
box -3 -3 3 3
use FILL  FILL_494
timestamp 1682952543
transform 1 0 1320 0 1 3370
box -8 -3 16 105
use FILL  FILL_495
timestamp 1682952543
transform 1 0 1328 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1780
timestamp 1682952543
transform 1 0 1348 0 1 3375
box -3 -3 3 3
use FILL  FILL_496
timestamp 1682952543
transform 1 0 1336 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_63
timestamp 1682952543
transform -1 0 1384 0 1 3370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1682952543
transform 1 0 1384 0 1 3370
box -8 -3 104 105
use INVX2  INVX2_125
timestamp 1682952543
transform -1 0 1496 0 1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_64
timestamp 1682952543
transform 1 0 1496 0 1 3370
box -8 -3 46 105
use FILL  FILL_497
timestamp 1682952543
transform 1 0 1536 0 1 3370
box -8 -3 16 105
use FILL  FILL_498
timestamp 1682952543
transform 1 0 1544 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_131
timestamp 1682952543
transform 1 0 1552 0 1 3370
box -8 -3 46 105
use INVX2  INVX2_126
timestamp 1682952543
transform 1 0 1592 0 1 3370
box -9 -3 26 105
use FILL  FILL_499
timestamp 1682952543
transform 1 0 1608 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_67
timestamp 1682952543
transform 1 0 1616 0 1 3370
box -8 -3 46 105
use FILL  FILL_509
timestamp 1682952543
transform 1 0 1656 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_130
timestamp 1682952543
transform 1 0 1664 0 1 3370
box -9 -3 26 105
use FILL  FILL_510
timestamp 1682952543
transform 1 0 1680 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1682952543
transform -1 0 1784 0 1 3370
box -8 -3 104 105
use FILL  FILL_511
timestamp 1682952543
transform 1 0 1784 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_124
timestamp 1682952543
transform -1 0 1888 0 1 3370
box -8 -3 104 105
use FILL  FILL_512
timestamp 1682952543
transform 1 0 1888 0 1 3370
box -8 -3 16 105
use FILL  FILL_513
timestamp 1682952543
transform 1 0 1896 0 1 3370
box -8 -3 16 105
use FILL  FILL_514
timestamp 1682952543
transform 1 0 1904 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_131
timestamp 1682952543
transform 1 0 1912 0 1 3370
box -9 -3 26 105
use M3_M2  M3_M2_1781
timestamp 1682952543
transform 1 0 1948 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_1782
timestamp 1682952543
transform 1 0 2020 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_125
timestamp 1682952543
transform 1 0 1928 0 1 3370
box -8 -3 104 105
use FILL  FILL_515
timestamp 1682952543
transform 1 0 2024 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1682952543
transform -1 0 2128 0 1 3370
box -8 -3 104 105
use FILL  FILL_516
timestamp 1682952543
transform 1 0 2128 0 1 3370
box -8 -3 16 105
use BUFX2  BUFX2_10
timestamp 1682952543
transform 1 0 2136 0 1 3370
box -5 -3 28 105
use FILL  FILL_532
timestamp 1682952543
transform 1 0 2160 0 1 3370
box -8 -3 16 105
use FILL  FILL_533
timestamp 1682952543
transform 1 0 2168 0 1 3370
box -8 -3 16 105
use FILL  FILL_534
timestamp 1682952543
transform 1 0 2176 0 1 3370
box -8 -3 16 105
use FILL  FILL_535
timestamp 1682952543
transform 1 0 2184 0 1 3370
box -8 -3 16 105
use FILL  FILL_536
timestamp 1682952543
transform 1 0 2192 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_135
timestamp 1682952543
transform 1 0 2200 0 1 3370
box -9 -3 26 105
use FILL  FILL_537
timestamp 1682952543
transform 1 0 2216 0 1 3370
box -8 -3 16 105
use FILL  FILL_538
timestamp 1682952543
transform 1 0 2224 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_136
timestamp 1682952543
transform 1 0 2232 0 1 3370
box -9 -3 26 105
use FILL  FILL_539
timestamp 1682952543
transform 1 0 2248 0 1 3370
box -8 -3 16 105
use FILL  FILL_543
timestamp 1682952543
transform 1 0 2256 0 1 3370
box -8 -3 16 105
use FILL  FILL_545
timestamp 1682952543
transform 1 0 2264 0 1 3370
box -8 -3 16 105
use FILL  FILL_546
timestamp 1682952543
transform 1 0 2272 0 1 3370
box -8 -3 16 105
use FILL  FILL_547
timestamp 1682952543
transform 1 0 2280 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_133
timestamp 1682952543
transform 1 0 2288 0 1 3370
box -8 -3 46 105
use FILL  FILL_548
timestamp 1682952543
transform 1 0 2328 0 1 3370
box -8 -3 16 105
use FILL  FILL_549
timestamp 1682952543
transform 1 0 2336 0 1 3370
box -8 -3 16 105
use FILL  FILL_550
timestamp 1682952543
transform 1 0 2344 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_134
timestamp 1682952543
transform 1 0 2352 0 1 3370
box -8 -3 46 105
use FILL  FILL_551
timestamp 1682952543
transform 1 0 2392 0 1 3370
box -8 -3 16 105
use FILL  FILL_552
timestamp 1682952543
transform 1 0 2400 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_24
timestamp 1682952543
transform 1 0 2408 0 1 3370
box -8 -3 34 105
use OAI21X1  OAI21X1_25
timestamp 1682952543
transform 1 0 2440 0 1 3370
box -8 -3 34 105
use INVX2  INVX2_137
timestamp 1682952543
transform 1 0 2472 0 1 3370
box -9 -3 26 105
use OAI21X1  OAI21X1_26
timestamp 1682952543
transform -1 0 2520 0 1 3370
box -8 -3 34 105
use FILL  FILL_553
timestamp 1682952543
transform 1 0 2520 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_27
timestamp 1682952543
transform -1 0 2560 0 1 3370
box -8 -3 34 105
use NAND2X1  NAND2X1_10
timestamp 1682952543
transform 1 0 2560 0 1 3370
box -8 -3 32 105
use FILL  FILL_554
timestamp 1682952543
transform 1 0 2584 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1783
timestamp 1682952543
transform 1 0 2612 0 1 3375
box -3 -3 3 3
use OAI21X1  OAI21X1_28
timestamp 1682952543
transform 1 0 2592 0 1 3370
box -8 -3 34 105
use NAND2X1  NAND2X1_11
timestamp 1682952543
transform 1 0 2624 0 1 3370
box -8 -3 32 105
use FILL  FILL_555
timestamp 1682952543
transform 1 0 2648 0 1 3370
box -8 -3 16 105
use FILL  FILL_556
timestamp 1682952543
transform 1 0 2656 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_12
timestamp 1682952543
transform -1 0 2688 0 1 3370
box -8 -3 32 105
use FILL  FILL_557
timestamp 1682952543
transform 1 0 2688 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_29
timestamp 1682952543
transform 1 0 2696 0 1 3370
box -8 -3 34 105
use FILL  FILL_558
timestamp 1682952543
transform 1 0 2728 0 1 3370
box -8 -3 16 105
use FILL  FILL_559
timestamp 1682952543
transform 1 0 2736 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_13
timestamp 1682952543
transform 1 0 2744 0 1 3370
box -8 -3 32 105
use FILL  FILL_560
timestamp 1682952543
transform 1 0 2768 0 1 3370
box -8 -3 16 105
use FILL  FILL_561
timestamp 1682952543
transform 1 0 2776 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_138
timestamp 1682952543
transform -1 0 2800 0 1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_131
timestamp 1682952543
transform -1 0 2896 0 1 3370
box -8 -3 104 105
use FILL  FILL_562
timestamp 1682952543
transform 1 0 2896 0 1 3370
box -8 -3 16 105
use FILL  FILL_563
timestamp 1682952543
transform 1 0 2904 0 1 3370
box -8 -3 16 105
use FILL  FILL_564
timestamp 1682952543
transform 1 0 2912 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_135
timestamp 1682952543
transform 1 0 2920 0 1 3370
box -8 -3 46 105
use M3_M2  M3_M2_1784
timestamp 1682952543
transform 1 0 2988 0 1 3375
box -3 -3 3 3
use OAI21X1  OAI21X1_30
timestamp 1682952543
transform 1 0 2960 0 1 3370
box -8 -3 34 105
use FILL  FILL_565
timestamp 1682952543
transform 1 0 2992 0 1 3370
box -8 -3 16 105
use FILL  FILL_566
timestamp 1682952543
transform 1 0 3000 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_139
timestamp 1682952543
transform -1 0 3024 0 1 3370
box -9 -3 26 105
use FILL  FILL_567
timestamp 1682952543
transform 1 0 3024 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_14
timestamp 1682952543
transform 1 0 3032 0 1 3370
box -8 -3 32 105
use FILL  FILL_568
timestamp 1682952543
transform 1 0 3056 0 1 3370
box -8 -3 16 105
use FILL  FILL_569
timestamp 1682952543
transform 1 0 3064 0 1 3370
box -8 -3 16 105
use FILL  FILL_570
timestamp 1682952543
transform 1 0 3072 0 1 3370
box -8 -3 16 105
use FILL  FILL_571
timestamp 1682952543
transform 1 0 3080 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1682952543
transform 1 0 3088 0 1 3370
box -8 -3 32 105
use FILL  FILL_572
timestamp 1682952543
transform 1 0 3112 0 1 3370
box -8 -3 16 105
use FILL  FILL_573
timestamp 1682952543
transform 1 0 3120 0 1 3370
box -8 -3 16 105
use FILL  FILL_574
timestamp 1682952543
transform 1 0 3128 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_31
timestamp 1682952543
transform -1 0 3168 0 1 3370
box -8 -3 34 105
use FILL  FILL_575
timestamp 1682952543
transform 1 0 3168 0 1 3370
box -8 -3 16 105
use FILL  FILL_576
timestamp 1682952543
transform 1 0 3176 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_140
timestamp 1682952543
transform 1 0 3184 0 1 3370
box -9 -3 26 105
use OAI22X1  OAI22X1_136
timestamp 1682952543
transform 1 0 3200 0 1 3370
box -8 -3 46 105
use FILL  FILL_577
timestamp 1682952543
transform 1 0 3240 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1785
timestamp 1682952543
transform 1 0 3260 0 1 3375
box -3 -3 3 3
use FILL  FILL_578
timestamp 1682952543
transform 1 0 3248 0 1 3370
box -8 -3 16 105
use FILL  FILL_588
timestamp 1682952543
transform 1 0 3256 0 1 3370
box -8 -3 16 105
use FILL  FILL_590
timestamp 1682952543
transform 1 0 3264 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_148
timestamp 1682952543
transform -1 0 3288 0 1 3370
box -9 -3 26 105
use FILL  FILL_591
timestamp 1682952543
transform 1 0 3288 0 1 3370
box -8 -3 16 105
use FILL  FILL_594
timestamp 1682952543
transform 1 0 3296 0 1 3370
box -8 -3 16 105
use FILL  FILL_595
timestamp 1682952543
transform 1 0 3304 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1786
timestamp 1682952543
transform 1 0 3332 0 1 3375
box -3 -3 3 3
use NAND2X1  NAND2X1_19
timestamp 1682952543
transform -1 0 3336 0 1 3370
box -8 -3 32 105
use FILL  FILL_596
timestamp 1682952543
transform 1 0 3336 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_36
timestamp 1682952543
transform -1 0 3376 0 1 3370
box -8 -3 34 105
use FILL  FILL_597
timestamp 1682952543
transform 1 0 3376 0 1 3370
box -8 -3 16 105
use FILL  FILL_598
timestamp 1682952543
transform 1 0 3384 0 1 3370
box -8 -3 16 105
use FILL  FILL_599
timestamp 1682952543
transform 1 0 3392 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_145
timestamp 1682952543
transform 1 0 3400 0 1 3370
box -8 -3 46 105
use FILL  FILL_600
timestamp 1682952543
transform 1 0 3440 0 1 3370
box -8 -3 16 105
use FILL  FILL_601
timestamp 1682952543
transform 1 0 3448 0 1 3370
box -8 -3 16 105
use FILL  FILL_602
timestamp 1682952543
transform 1 0 3456 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_150
timestamp 1682952543
transform 1 0 3464 0 1 3370
box -9 -3 26 105
use INVX2  INVX2_151
timestamp 1682952543
transform -1 0 3496 0 1 3370
box -9 -3 26 105
use FILL  FILL_603
timestamp 1682952543
transform 1 0 3496 0 1 3370
box -8 -3 16 105
use FILL  FILL_604
timestamp 1682952543
transform 1 0 3504 0 1 3370
box -8 -3 16 105
use FILL  FILL_605
timestamp 1682952543
transform 1 0 3512 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_152
timestamp 1682952543
transform 1 0 3520 0 1 3370
box -9 -3 26 105
use AND2X2  AND2X2_0
timestamp 1682952543
transform 1 0 3536 0 1 3370
box -8 -3 40 105
use OAI22X1  OAI22X1_146
timestamp 1682952543
transform 1 0 3568 0 1 3370
box -8 -3 46 105
use FILL  FILL_606
timestamp 1682952543
transform 1 0 3608 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1787
timestamp 1682952543
transform 1 0 3652 0 1 3375
box -3 -3 3 3
use OAI21X1  OAI21X1_37
timestamp 1682952543
transform 1 0 3616 0 1 3370
box -8 -3 34 105
use FILL  FILL_607
timestamp 1682952543
transform 1 0 3648 0 1 3370
box -8 -3 16 105
use FILL  FILL_608
timestamp 1682952543
transform 1 0 3656 0 1 3370
box -8 -3 16 105
use FILL  FILL_609
timestamp 1682952543
transform 1 0 3664 0 1 3370
box -8 -3 16 105
use FILL  FILL_610
timestamp 1682952543
transform 1 0 3672 0 1 3370
box -8 -3 16 105
use FILL  FILL_619
timestamp 1682952543
transform 1 0 3680 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_148
timestamp 1682952543
transform 1 0 3688 0 1 3370
box -8 -3 46 105
use FILL  FILL_621
timestamp 1682952543
transform 1 0 3728 0 1 3370
box -8 -3 16 105
use FILL  FILL_622
timestamp 1682952543
transform 1 0 3736 0 1 3370
box -8 -3 16 105
use FILL  FILL_623
timestamp 1682952543
transform 1 0 3744 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_149
timestamp 1682952543
transform 1 0 3752 0 1 3370
box -8 -3 46 105
use FILL  FILL_624
timestamp 1682952543
transform 1 0 3792 0 1 3370
box -8 -3 16 105
use FILL  FILL_625
timestamp 1682952543
transform 1 0 3800 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_150
timestamp 1682952543
transform 1 0 3808 0 1 3370
box -8 -3 46 105
use FILL  FILL_626
timestamp 1682952543
transform 1 0 3848 0 1 3370
box -8 -3 16 105
use FILL  FILL_627
timestamp 1682952543
transform 1 0 3856 0 1 3370
box -8 -3 16 105
use FILL  FILL_628
timestamp 1682952543
transform 1 0 3864 0 1 3370
box -8 -3 16 105
use FILL  FILL_629
timestamp 1682952543
transform 1 0 3872 0 1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_21
timestamp 1682952543
transform 1 0 3880 0 1 3370
box -8 -3 32 105
use FILL  FILL_630
timestamp 1682952543
transform 1 0 3904 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_1788
timestamp 1682952543
transform 1 0 3924 0 1 3375
box -3 -3 3 3
use OAI21X1  OAI21X1_39
timestamp 1682952543
transform -1 0 3944 0 1 3370
box -8 -3 34 105
use M3_M2  M3_M2_1789
timestamp 1682952543
transform 1 0 3956 0 1 3375
box -3 -3 3 3
use FILL  FILL_631
timestamp 1682952543
transform 1 0 3944 0 1 3370
box -8 -3 16 105
use FILL  FILL_632
timestamp 1682952543
transform 1 0 3952 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_151
timestamp 1682952543
transform 1 0 3960 0 1 3370
box -8 -3 46 105
use FILL  FILL_633
timestamp 1682952543
transform 1 0 4000 0 1 3370
box -8 -3 16 105
use FILL  FILL_636
timestamp 1682952543
transform 1 0 4008 0 1 3370
box -8 -3 16 105
use FILL  FILL_637
timestamp 1682952543
transform 1 0 4016 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_156
timestamp 1682952543
transform 1 0 4024 0 1 3370
box -8 -3 46 105
use FILL  FILL_638
timestamp 1682952543
transform 1 0 4064 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_158
timestamp 1682952543
transform -1 0 4088 0 1 3370
box -9 -3 26 105
use FILL  FILL_639
timestamp 1682952543
transform 1 0 4088 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_159
timestamp 1682952543
transform -1 0 4112 0 1 3370
box -9 -3 26 105
use FILL  FILL_640
timestamp 1682952543
transform 1 0 4112 0 1 3370
box -8 -3 16 105
use FILL  FILL_641
timestamp 1682952543
transform 1 0 4120 0 1 3370
box -8 -3 16 105
use FILL  FILL_642
timestamp 1682952543
transform 1 0 4128 0 1 3370
box -8 -3 16 105
use FILL  FILL_643
timestamp 1682952543
transform 1 0 4136 0 1 3370
box -8 -3 16 105
use FILL  FILL_644
timestamp 1682952543
transform 1 0 4144 0 1 3370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_15
timestamp 1682952543
transform 1 0 4177 0 1 3370
box -10 -3 10 3
use M3_M2  M3_M2_1790
timestamp 1682952543
transform 1 0 140 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1817
timestamp 1682952543
transform 1 0 148 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1851
timestamp 1682952543
transform 1 0 84 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1791
timestamp 1682952543
transform 1 0 180 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_1973
timestamp 1682952543
transform 1 0 132 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1682952543
transform 1 0 164 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1975
timestamp 1682952543
transform 1 0 172 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1931
timestamp 1682952543
transform 1 0 132 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1682952543
transform 1 0 172 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1682952543
transform 1 0 164 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1682952543
transform 1 0 220 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1682952543
transform 1 0 204 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1844
timestamp 1682952543
transform 1 0 276 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1852
timestamp 1682952543
transform 1 0 188 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1853
timestamp 1682952543
transform 1 0 196 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1854
timestamp 1682952543
transform 1 0 212 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1855
timestamp 1682952543
transform 1 0 220 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1856
timestamp 1682952543
transform 1 0 244 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1682952543
transform 1 0 252 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1858
timestamp 1682952543
transform 1 0 276 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1682952543
transform 1 0 284 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1682952543
transform 1 0 180 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1682952543
transform 1 0 204 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1978
timestamp 1682952543
transform 1 0 228 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1981
timestamp 1682952543
transform 1 0 196 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1682952543
transform 1 0 236 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_1979
timestamp 1682952543
transform 1 0 244 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1909
timestamp 1682952543
transform 1 0 252 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_1980
timestamp 1682952543
transform 1 0 260 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1981
timestamp 1682952543
transform 1 0 276 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1860
timestamp 1682952543
transform 1 0 300 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1682952543
transform 1 0 300 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1793
timestamp 1682952543
transform 1 0 332 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1794
timestamp 1682952543
transform 1 0 364 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1795
timestamp 1682952543
transform 1 0 404 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_1861
timestamp 1682952543
transform 1 0 324 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1862
timestamp 1682952543
transform 1 0 412 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1682952543
transform 1 0 308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1682952543
transform 1 0 348 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1985
timestamp 1682952543
transform 1 0 404 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1933
timestamp 1682952543
transform 1 0 308 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1682952543
transform 1 0 348 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1682952543
transform 1 0 444 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1863
timestamp 1682952543
transform 1 0 436 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1864
timestamp 1682952543
transform 1 0 452 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1682952543
transform 1 0 468 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1866
timestamp 1682952543
transform 1 0 476 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1682952543
transform 1 0 428 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1796
timestamp 1682952543
transform 1 0 532 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1846
timestamp 1682952543
transform 1 0 500 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1987
timestamp 1682952543
transform 1 0 444 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1682952543
transform 1 0 460 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1910
timestamp 1682952543
transform 1 0 476 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_1867
timestamp 1682952543
transform 1 0 500 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1682952543
transform 1 0 484 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1682952543
transform 1 0 524 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1982
timestamp 1682952543
transform 1 0 444 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1682952543
transform 1 0 460 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1911
timestamp 1682952543
transform 1 0 548 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_1991
timestamp 1682952543
transform 1 0 580 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1935
timestamp 1682952543
transform 1 0 484 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1936
timestamp 1682952543
transform 1 0 524 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1682952543
transform 1 0 580 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1847
timestamp 1682952543
transform 1 0 620 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1868
timestamp 1682952543
transform 1 0 636 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1682952543
transform 1 0 620 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1819
timestamp 1682952543
transform 1 0 700 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1869
timestamp 1682952543
transform 1 0 660 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1682952543
transform 1 0 676 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1682952543
transform 1 0 644 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1893
timestamp 1682952543
transform 1 0 724 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1682952543
transform 1 0 748 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1871
timestamp 1682952543
transform 1 0 764 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1872
timestamp 1682952543
transform 1 0 780 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1682952543
transform 1 0 724 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1995
timestamp 1682952543
transform 1 0 756 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1682952543
transform 1 0 772 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1682952543
transform 1 0 788 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1983
timestamp 1682952543
transform 1 0 660 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1682952543
transform 1 0 764 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1939
timestamp 1682952543
transform 1 0 788 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1682952543
transform 1 0 756 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1985
timestamp 1682952543
transform 1 0 772 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2008
timestamp 1682952543
transform 1 0 772 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2009
timestamp 1682952543
transform 1 0 788 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1682952543
transform 1 0 828 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1849
timestamp 1682952543
transform 1 0 852 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1873
timestamp 1682952543
transform 1 0 828 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1874
timestamp 1682952543
transform 1 0 836 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1682952543
transform 1 0 852 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1682952543
transform 1 0 820 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1940
timestamp 1682952543
transform 1 0 812 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1682952543
transform 1 0 804 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1682952543
transform 1 0 820 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_1999
timestamp 1682952543
transform 1 0 844 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1941
timestamp 1682952543
transform 1 0 844 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_1876
timestamp 1682952543
transform 1 0 868 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2000
timestamp 1682952543
transform 1 0 876 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1942
timestamp 1682952543
transform 1 0 868 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1682952543
transform 1 0 876 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1797
timestamp 1682952543
transform 1 0 948 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1798
timestamp 1682952543
transform 1 0 980 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1820
timestamp 1682952543
transform 1 0 908 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1682952543
transform 1 0 956 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1822
timestamp 1682952543
transform 1 0 988 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1682952543
transform 1 0 916 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1682952543
transform 1 0 924 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1896
timestamp 1682952543
transform 1 0 964 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1877
timestamp 1682952543
transform 1 0 988 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1682952543
transform 1 0 900 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1682952543
transform 1 0 908 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1912
timestamp 1682952543
transform 1 0 924 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2003
timestamp 1682952543
transform 1 0 940 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1943
timestamp 1682952543
transform 1 0 900 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1682952543
transform 1 0 940 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1823
timestamp 1682952543
transform 1 0 1012 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1878
timestamp 1682952543
transform 1 0 1012 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1682952543
transform 1 0 1036 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1851
timestamp 1682952543
transform 1 0 1132 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1897
timestamp 1682952543
transform 1 0 1116 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1879
timestamp 1682952543
transform 1 0 1124 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1682952543
transform 1 0 1108 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1682952543
transform 1 0 1116 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1682952543
transform 1 0 1132 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1682952543
transform 1 0 1148 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1945
timestamp 1682952543
transform 1 0 1116 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2023
timestamp 1682952543
transform 1 0 1116 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_1880
timestamp 1682952543
transform 1 0 1172 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1824
timestamp 1682952543
transform 1 0 1212 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1881
timestamp 1682952543
transform 1 0 1196 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1898
timestamp 1682952543
transform 1 0 1204 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1882
timestamp 1682952543
transform 1 0 1212 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1682952543
transform 1 0 1188 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1913
timestamp 1682952543
transform 1 0 1196 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1682952543
transform 1 0 1228 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1883
timestamp 1682952543
transform 1 0 1228 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1682952543
transform 1 0 1212 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1682952543
transform 1 0 1220 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1853
timestamp 1682952543
transform 1 0 1268 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1854
timestamp 1682952543
transform 1 0 1300 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1884
timestamp 1682952543
transform 1 0 1268 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1914
timestamp 1682952543
transform 1 0 1308 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2012
timestamp 1682952543
transform 1 0 1316 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1682952543
transform 1 0 1348 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1682952543
transform 1 0 1356 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1946
timestamp 1682952543
transform 1 0 1316 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1947
timestamp 1682952543
transform 1 0 1356 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1988
timestamp 1682952543
transform 1 0 1308 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1682952543
transform 1 0 1332 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1682952543
transform 1 0 1372 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1885
timestamp 1682952543
transform 1 0 1364 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1682952543
transform 1 0 1372 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1682952543
transform 1 0 1380 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1899
timestamp 1682952543
transform 1 0 1388 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1888
timestamp 1682952543
transform 1 0 1396 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1682952543
transform 1 0 1364 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1682952543
transform 1 0 1388 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1915
timestamp 1682952543
transform 1 0 1396 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_1889
timestamp 1682952543
transform 1 0 1420 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1682952543
transform 1 0 1404 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1682952543
transform 1 0 1468 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2019
timestamp 1682952543
transform 1 0 1500 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1682952543
transform 1 0 1508 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1990
timestamp 1682952543
transform 1 0 1364 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1682952543
transform 1 0 1468 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1991
timestamp 1682952543
transform 1 0 1500 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2024
timestamp 1682952543
transform 1 0 1492 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_1890
timestamp 1682952543
transform 1 0 1532 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1682952543
transform 1 0 1532 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1949
timestamp 1682952543
transform 1 0 1532 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2025
timestamp 1682952543
transform 1 0 1532 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1826
timestamp 1682952543
transform 1 0 1556 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1827
timestamp 1682952543
transform 1 0 1596 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1891
timestamp 1682952543
transform 1 0 1556 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1892
timestamp 1682952543
transform 1 0 1564 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1900
timestamp 1682952543
transform 1 0 1588 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1893
timestamp 1682952543
transform 1 0 1604 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2022
timestamp 1682952543
transform 1 0 1548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1682952543
transform 1 0 1572 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1682952543
transform 1 0 1588 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1682952543
transform 1 0 1596 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1992
timestamp 1682952543
transform 1 0 1564 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_1894
timestamp 1682952543
transform 1 0 1628 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1799
timestamp 1682952543
transform 1 0 1668 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_1895
timestamp 1682952543
transform 1 0 1716 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2026
timestamp 1682952543
transform 1 0 1684 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1950
timestamp 1682952543
transform 1 0 1684 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1682952543
transform 1 0 1716 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2027
timestamp 1682952543
transform 1 0 1732 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1951
timestamp 1682952543
transform 1 0 1732 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2010
timestamp 1682952543
transform 1 0 1748 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1828
timestamp 1682952543
transform 1 0 1772 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1855
timestamp 1682952543
transform 1 0 1788 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1896
timestamp 1682952543
transform 1 0 1764 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1897
timestamp 1682952543
transform 1 0 1772 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1898
timestamp 1682952543
transform 1 0 1796 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1682952543
transform 1 0 1804 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1900
timestamp 1682952543
transform 1 0 1812 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1916
timestamp 1682952543
transform 1 0 1764 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2028
timestamp 1682952543
transform 1 0 1772 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1917
timestamp 1682952543
transform 1 0 1780 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2029
timestamp 1682952543
transform 1 0 1788 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1952
timestamp 1682952543
transform 1 0 1772 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1682952543
transform 1 0 1788 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1682952543
transform 1 0 1780 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1682952543
transform 1 0 1828 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1953
timestamp 1682952543
transform 1 0 1820 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1682952543
transform 1 0 1924 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1901
timestamp 1682952543
transform 1 0 1924 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2030
timestamp 1682952543
transform 1 0 1836 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1682952543
transform 1 0 1844 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1682952543
transform 1 0 1900 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1994
timestamp 1682952543
transform 1 0 1924 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2033
timestamp 1682952543
transform 1 0 1956 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1901
timestamp 1682952543
transform 1 0 1972 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1858
timestamp 1682952543
transform 1 0 2020 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1859
timestamp 1682952543
transform 1 0 2036 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1902
timestamp 1682952543
transform 1 0 2020 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1829
timestamp 1682952543
transform 1 0 2116 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1860
timestamp 1682952543
transform 1 0 2116 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2034
timestamp 1682952543
transform 1 0 2004 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2035
timestamp 1682952543
transform 1 0 2044 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2036
timestamp 1682952543
transform 1 0 2100 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2037
timestamp 1682952543
transform 1 0 2108 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2027
timestamp 1682952543
transform 1 0 2100 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_1903
timestamp 1682952543
transform 1 0 2132 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1800
timestamp 1682952543
transform 1 0 2244 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1682952543
transform 1 0 2164 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1862
timestamp 1682952543
transform 1 0 2212 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1904
timestamp 1682952543
transform 1 0 2164 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2038
timestamp 1682952543
transform 1 0 2212 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1682952543
transform 1 0 2244 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1954
timestamp 1682952543
transform 1 0 2164 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1682952543
transform 1 0 2196 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2013
timestamp 1682952543
transform 1 0 2244 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2028
timestamp 1682952543
transform 1 0 2172 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1863
timestamp 1682952543
transform 1 0 2284 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1905
timestamp 1682952543
transform 1 0 2268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1906
timestamp 1682952543
transform 1 0 2284 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1682952543
transform 1 0 2300 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2040
timestamp 1682952543
transform 1 0 2260 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1918
timestamp 1682952543
transform 1 0 2268 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2041
timestamp 1682952543
transform 1 0 2292 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1830
timestamp 1682952543
transform 1 0 2324 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1682952543
transform 1 0 2316 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1908
timestamp 1682952543
transform 1 0 2324 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1909
timestamp 1682952543
transform 1 0 2340 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1682952543
transform 1 0 2356 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2042
timestamp 1682952543
transform 1 0 2332 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2043
timestamp 1682952543
transform 1 0 2348 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1919
timestamp 1682952543
transform 1 0 2356 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_1911
timestamp 1682952543
transform 1 0 2380 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1801
timestamp 1682952543
transform 1 0 2436 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1802
timestamp 1682952543
transform 1 0 2492 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1682952543
transform 1 0 2452 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1831
timestamp 1682952543
transform 1 0 2524 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1865
timestamp 1682952543
transform 1 0 2508 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1912
timestamp 1682952543
transform 1 0 2404 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1682952543
transform 1 0 2492 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1914
timestamp 1682952543
transform 1 0 2508 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1682952543
transform 1 0 2524 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1682952543
transform 1 0 2532 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1682952543
transform 1 0 2452 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1682952543
transform 1 0 2484 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2046
timestamp 1682952543
transform 1 0 2492 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1682952543
transform 1 0 2500 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1682952543
transform 1 0 2516 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1955
timestamp 1682952543
transform 1 0 2404 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1682952543
transform 1 0 2492 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1682952543
transform 1 0 2524 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2014
timestamp 1682952543
transform 1 0 2516 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_1917
timestamp 1682952543
transform 1 0 2548 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2049
timestamp 1682952543
transform 1 0 2548 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1832
timestamp 1682952543
transform 1 0 2572 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1918
timestamp 1682952543
transform 1 0 2580 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1833
timestamp 1682952543
transform 1 0 2596 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1919
timestamp 1682952543
transform 1 0 2596 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2050
timestamp 1682952543
transform 1 0 2564 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1682952543
transform 1 0 2580 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1682952543
transform 1 0 2588 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1682952543
transform 1 0 2556 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2029
timestamp 1682952543
transform 1 0 2548 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1682952543
transform 1 0 2580 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1682952543
transform 1 0 2596 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2108
timestamp 1682952543
transform 1 0 2596 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2030
timestamp 1682952543
transform 1 0 2604 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1682952543
transform 1 0 2628 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1920
timestamp 1682952543
transform 1 0 2620 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1958
timestamp 1682952543
transform 1 0 2620 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1803
timestamp 1682952543
transform 1 0 2660 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1866
timestamp 1682952543
transform 1 0 2652 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1835
timestamp 1682952543
transform 1 0 2676 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1921
timestamp 1682952543
transform 1 0 2652 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1922
timestamp 1682952543
transform 1 0 2668 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1923
timestamp 1682952543
transform 1 0 2676 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2053
timestamp 1682952543
transform 1 0 2636 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2054
timestamp 1682952543
transform 1 0 2660 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1804
timestamp 1682952543
transform 1 0 2708 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_1924
timestamp 1682952543
transform 1 0 2700 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1925
timestamp 1682952543
transform 1 0 2708 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1682952543
transform 1 0 2692 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1959
timestamp 1682952543
transform 1 0 2676 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1995
timestamp 1682952543
transform 1 0 2660 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1682952543
transform 1 0 2700 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1682952543
transform 1 0 2756 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_1926
timestamp 1682952543
transform 1 0 2748 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1927
timestamp 1682952543
transform 1 0 2756 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1682952543
transform 1 0 2780 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1682952543
transform 1 0 2732 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1923
timestamp 1682952543
transform 1 0 2772 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2109
timestamp 1682952543
transform 1 0 2756 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2110
timestamp 1682952543
transform 1 0 2772 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_1960
timestamp 1682952543
transform 1 0 2780 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1996
timestamp 1682952543
transform 1 0 2756 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1806
timestamp 1682952543
transform 1 0 2812 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1682952543
transform 1 0 2804 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1682952543
transform 1 0 2844 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1929
timestamp 1682952543
transform 1 0 2812 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1682952543
transform 1 0 2828 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1682952543
transform 1 0 2844 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2057
timestamp 1682952543
transform 1 0 2820 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2058
timestamp 1682952543
transform 1 0 2836 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2059
timestamp 1682952543
transform 1 0 2852 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2111
timestamp 1682952543
transform 1 0 2804 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_1997
timestamp 1682952543
transform 1 0 2804 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1682952543
transform 1 0 2868 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1682952543
transform 1 0 2940 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1682952543
transform 1 0 2900 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1870
timestamp 1682952543
transform 1 0 2924 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1809
timestamp 1682952543
transform 1 0 3044 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1682952543
transform 1 0 2980 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1682952543
transform 1 0 3052 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1932
timestamp 1682952543
transform 1 0 2868 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1682952543
transform 1 0 2884 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1682952543
transform 1 0 2900 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1682952543
transform 1 0 2924 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1682952543
transform 1 0 2940 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1682952543
transform 1 0 2956 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1682952543
transform 1 0 3044 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2060
timestamp 1682952543
transform 1 0 2868 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1682952543
transform 1 0 2876 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2062
timestamp 1682952543
transform 1 0 2892 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1961
timestamp 1682952543
transform 1 0 2852 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1682952543
transform 1 0 2900 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2063
timestamp 1682952543
transform 1 0 2916 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1682952543
transform 1 0 2932 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1962
timestamp 1682952543
transform 1 0 2876 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1682952543
transform 1 0 2916 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_2065
timestamp 1682952543
transform 1 0 2980 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1682952543
transform 1 0 3036 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1998
timestamp 1682952543
transform 1 0 3020 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1810
timestamp 1682952543
transform 1 0 3100 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1682952543
transform 1 0 3116 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1874
timestamp 1682952543
transform 1 0 3164 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1939
timestamp 1682952543
transform 1 0 3068 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1682952543
transform 1 0 3084 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1682952543
transform 1 0 3100 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1682952543
transform 1 0 3116 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1925
timestamp 1682952543
transform 1 0 3068 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1682952543
transform 1 0 3212 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1682952543
transform 1 0 3228 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1943
timestamp 1682952543
transform 1 0 3212 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1682952543
transform 1 0 3228 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1682952543
transform 1 0 3244 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2067
timestamp 1682952543
transform 1 0 3076 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1682952543
transform 1 0 3100 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2069
timestamp 1682952543
transform 1 0 3164 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1682952543
transform 1 0 3196 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1682952543
transform 1 0 3204 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2031
timestamp 1682952543
transform 1 0 3052 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1682952543
transform 1 0 3100 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1964
timestamp 1682952543
transform 1 0 3140 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1682952543
transform 1 0 3180 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1682952543
transform 1 0 3076 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1999
timestamp 1682952543
transform 1 0 3116 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1682952543
transform 1 0 3156 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1682952543
transform 1 0 3204 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2072
timestamp 1682952543
transform 1 0 3236 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1926
timestamp 1682952543
transform 1 0 3244 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2073
timestamp 1682952543
transform 1 0 3252 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1967
timestamp 1682952543
transform 1 0 3236 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_1946
timestamp 1682952543
transform 1 0 3260 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2018
timestamp 1682952543
transform 1 0 3252 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1876
timestamp 1682952543
transform 1 0 3276 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1682952543
transform 1 0 3324 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1682952543
transform 1 0 3372 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1947
timestamp 1682952543
transform 1 0 3324 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2074
timestamp 1682952543
transform 1 0 3300 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2075
timestamp 1682952543
transform 1 0 3308 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1682952543
transform 1 0 3372 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1968
timestamp 1682952543
transform 1 0 3356 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1836
timestamp 1682952543
transform 1 0 3428 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1682952543
transform 1 0 3444 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1682952543
transform 1 0 3460 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1948
timestamp 1682952543
transform 1 0 3428 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1682952543
transform 1 0 3444 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1903
timestamp 1682952543
transform 1 0 3452 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1950
timestamp 1682952543
transform 1 0 3460 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1881
timestamp 1682952543
transform 1 0 3508 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1682952543
transform 1 0 3532 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1951
timestamp 1682952543
transform 1 0 3492 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1952
timestamp 1682952543
transform 1 0 3524 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1682952543
transform 1 0 3532 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2077
timestamp 1682952543
transform 1 0 3436 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2078
timestamp 1682952543
transform 1 0 3452 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2079
timestamp 1682952543
transform 1 0 3468 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2080
timestamp 1682952543
transform 1 0 3484 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2081
timestamp 1682952543
transform 1 0 3500 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1682952543
transform 1 0 3516 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1969
timestamp 1682952543
transform 1 0 3452 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1682952543
transform 1 0 3428 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2032
timestamp 1682952543
transform 1 0 3324 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2033
timestamp 1682952543
transform 1 0 3348 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2034
timestamp 1682952543
transform 1 0 3404 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_1970
timestamp 1682952543
transform 1 0 3484 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1682952543
transform 1 0 3548 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1682952543
transform 1 0 3564 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2083
timestamp 1682952543
transform 1 0 3540 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1682952543
transform 1 0 3556 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1971
timestamp 1682952543
transform 1 0 3516 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1682952543
transform 1 0 3532 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2035
timestamp 1682952543
transform 1 0 3524 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1682952543
transform 1 0 3580 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1837
timestamp 1682952543
transform 1 0 3604 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_1954
timestamp 1682952543
transform 1 0 3604 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1682952543
transform 1 0 3604 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1973
timestamp 1682952543
transform 1 0 3620 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2112
timestamp 1682952543
transform 1 0 3628 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2019
timestamp 1682952543
transform 1 0 3628 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1838
timestamp 1682952543
transform 1 0 3644 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2086
timestamp 1682952543
transform 1 0 3668 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1884
timestamp 1682952543
transform 1 0 3692 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1955
timestamp 1682952543
transform 1 0 3692 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2087
timestamp 1682952543
transform 1 0 3692 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1812
timestamp 1682952543
transform 1 0 3732 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1682952543
transform 1 0 3716 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1839
timestamp 1682952543
transform 1 0 3748 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1682952543
transform 1 0 3756 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1956
timestamp 1682952543
transform 1 0 3716 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1905
timestamp 1682952543
transform 1 0 3724 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1957
timestamp 1682952543
transform 1 0 3732 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1906
timestamp 1682952543
transform 1 0 3740 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_1958
timestamp 1682952543
transform 1 0 3756 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1959
timestamp 1682952543
transform 1 0 3772 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1682952543
transform 1 0 3708 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1682952543
transform 1 0 3724 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1927
timestamp 1682952543
transform 1 0 3732 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2090
timestamp 1682952543
transform 1 0 3740 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2091
timestamp 1682952543
transform 1 0 3748 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2092
timestamp 1682952543
transform 1 0 3764 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2093
timestamp 1682952543
transform 1 0 3780 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2002
timestamp 1682952543
transform 1 0 3740 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1682952543
transform 1 0 3764 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2020
timestamp 1682952543
transform 1 0 3708 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1840
timestamp 1682952543
transform 1 0 3788 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1841
timestamp 1682952543
transform 1 0 3844 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1682952543
transform 1 0 3828 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1682952543
transform 1 0 3852 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1960
timestamp 1682952543
transform 1 0 3788 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1961
timestamp 1682952543
transform 1 0 3804 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1889
timestamp 1682952543
transform 1 0 3924 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1682952543
transform 1 0 3940 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1962
timestamp 1682952543
transform 1 0 3900 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1963
timestamp 1682952543
transform 1 0 3924 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1964
timestamp 1682952543
transform 1 0 3940 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1682952543
transform 1 0 3948 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1966
timestamp 1682952543
transform 1 0 3964 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1682952543
transform 1 0 3980 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1682952543
transform 1 0 3828 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2095
timestamp 1682952543
transform 1 0 3884 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2096
timestamp 1682952543
transform 1 0 3892 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2097
timestamp 1682952543
transform 1 0 3900 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2098
timestamp 1682952543
transform 1 0 3916 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2099
timestamp 1682952543
transform 1 0 3932 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1974
timestamp 1682952543
transform 1 0 3844 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1975
timestamp 1682952543
transform 1 0 3892 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1928
timestamp 1682952543
transform 1 0 3940 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2100
timestamp 1682952543
transform 1 0 3956 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2101
timestamp 1682952543
transform 1 0 3972 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1682952543
transform 1 0 3988 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1976
timestamp 1682952543
transform 1 0 3916 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1682952543
transform 1 0 3948 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1682952543
transform 1 0 3988 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1682952543
transform 1 0 3932 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_1813
timestamp 1682952543
transform 1 0 4020 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1842
timestamp 1682952543
transform 1 0 4044 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1682952543
transform 1 0 4028 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1968
timestamp 1682952543
transform 1 0 4004 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1682952543
transform 1 0 4012 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1682952543
transform 1 0 4028 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_1971
timestamp 1682952543
transform 1 0 4044 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2103
timestamp 1682952543
transform 1 0 4020 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1682952543
transform 1 0 4036 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2021
timestamp 1682952543
transform 1 0 4036 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1682952543
transform 1 0 4068 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1815
timestamp 1682952543
transform 1 0 4092 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1682952543
transform 1 0 4148 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_1843
timestamp 1682952543
transform 1 0 4060 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1682952543
transform 1 0 4092 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_1972
timestamp 1682952543
transform 1 0 4068 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_1907
timestamp 1682952543
transform 1 0 4156 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1682952543
transform 1 0 4068 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2105
timestamp 1682952543
transform 1 0 4092 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1930
timestamp 1682952543
transform 1 0 4108 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2106
timestamp 1682952543
transform 1 0 4148 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_1979
timestamp 1682952543
transform 1 0 4132 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1682952543
transform 1 0 4068 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1682952543
transform 1 0 4100 0 1 3305
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_16
timestamp 1682952543
transform 1 0 24 0 1 3270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_111
timestamp 1682952543
transform 1 0 72 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_115
timestamp 1682952543
transform -1 0 184 0 -1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_57
timestamp 1682952543
transform -1 0 224 0 -1 3370
box -8 -3 46 105
use INVX2  INVX2_116
timestamp 1682952543
transform -1 0 240 0 -1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_58
timestamp 1682952543
transform 1 0 240 0 -1 3370
box -8 -3 46 105
use INVX2  INVX2_117
timestamp 1682952543
transform 1 0 280 0 -1 3370
box -9 -3 26 105
use INVX2  INVX2_118
timestamp 1682952543
transform 1 0 296 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1682952543
transform 1 0 312 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_119
timestamp 1682952543
transform 1 0 408 0 -1 3370
box -9 -3 26 105
use FILL  FILL_461
timestamp 1682952543
transform 1 0 424 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_127
timestamp 1682952543
transform 1 0 432 0 -1 3370
box -8 -3 46 105
use INVX2  INVX2_120
timestamp 1682952543
transform 1 0 472 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1682952543
transform 1 0 488 0 -1 3370
box -8 -3 104 105
use FILL  FILL_462
timestamp 1682952543
transform 1 0 584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_463
timestamp 1682952543
transform 1 0 592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_465
timestamp 1682952543
transform 1 0 600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_467
timestamp 1682952543
transform 1 0 608 0 -1 3370
box -8 -3 16 105
use BUFX2  BUFX2_6
timestamp 1682952543
transform 1 0 616 0 -1 3370
box -5 -3 28 105
use BUFX2  BUFX2_7
timestamp 1682952543
transform 1 0 640 0 -1 3370
box -5 -3 28 105
use M3_M2  M3_M2_2036
timestamp 1682952543
transform 1 0 740 0 1 3275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_115
timestamp 1682952543
transform 1 0 664 0 -1 3370
box -8 -3 104 105
use OAI22X1  OAI22X1_129
timestamp 1682952543
transform 1 0 760 0 -1 3370
box -8 -3 46 105
use FILL  FILL_468
timestamp 1682952543
transform 1 0 800 0 -1 3370
box -8 -3 16 105
use FILL  FILL_470
timestamp 1682952543
transform 1 0 808 0 -1 3370
box -8 -3 16 105
use FILL  FILL_484
timestamp 1682952543
transform 1 0 816 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_61
timestamp 1682952543
transform 1 0 824 0 -1 3370
box -8 -3 46 105
use FILL  FILL_485
timestamp 1682952543
transform 1 0 864 0 -1 3370
box -8 -3 16 105
use FILL  FILL_486
timestamp 1682952543
transform 1 0 872 0 -1 3370
box -8 -3 16 105
use FILL  FILL_487
timestamp 1682952543
transform 1 0 880 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_124
timestamp 1682952543
transform 1 0 888 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1682952543
transform -1 0 1000 0 -1 3370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1682952543
transform 1 0 1000 0 -1 3370
box -8 -3 104 105
use FILL  FILL_488
timestamp 1682952543
transform 1 0 1096 0 -1 3370
box -8 -3 16 105
use FILL  FILL_489
timestamp 1682952543
transform 1 0 1104 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_62
timestamp 1682952543
transform 1 0 1112 0 -1 3370
box -8 -3 46 105
use FILL  FILL_490
timestamp 1682952543
transform 1 0 1152 0 -1 3370
box -8 -3 16 105
use FILL  FILL_500
timestamp 1682952543
transform 1 0 1160 0 -1 3370
box -8 -3 16 105
use FILL  FILL_501
timestamp 1682952543
transform 1 0 1168 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_132
timestamp 1682952543
transform -1 0 1216 0 -1 3370
box -8 -3 46 105
use FILL  FILL_502
timestamp 1682952543
transform 1 0 1216 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_127
timestamp 1682952543
transform 1 0 1224 0 -1 3370
box -9 -3 26 105
use FILL  FILL_503
timestamp 1682952543
transform 1 0 1240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_504
timestamp 1682952543
transform 1 0 1248 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1682952543
transform 1 0 1256 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_128
timestamp 1682952543
transform -1 0 1368 0 -1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_65
timestamp 1682952543
transform -1 0 1408 0 -1 3370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1682952543
transform 1 0 1408 0 -1 3370
box -8 -3 104 105
use BUFX2  BUFX2_8
timestamp 1682952543
transform 1 0 1504 0 -1 3370
box -5 -3 28 105
use FILL  FILL_505
timestamp 1682952543
transform 1 0 1528 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_129
timestamp 1682952543
transform -1 0 1552 0 -1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_66
timestamp 1682952543
transform -1 0 1592 0 -1 3370
box -8 -3 46 105
use FILL  FILL_506
timestamp 1682952543
transform 1 0 1592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_507
timestamp 1682952543
transform 1 0 1600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_508
timestamp 1682952543
transform 1 0 1608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_517
timestamp 1682952543
transform 1 0 1616 0 -1 3370
box -8 -3 16 105
use FILL  FILL_518
timestamp 1682952543
transform 1 0 1624 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1682952543
transform -1 0 1728 0 -1 3370
box -8 -3 104 105
use FILL  FILL_519
timestamp 1682952543
transform 1 0 1728 0 -1 3370
box -8 -3 16 105
use FILL  FILL_520
timestamp 1682952543
transform 1 0 1736 0 -1 3370
box -8 -3 16 105
use FILL  FILL_521
timestamp 1682952543
transform 1 0 1744 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_132
timestamp 1682952543
transform -1 0 1768 0 -1 3370
box -9 -3 26 105
use AOI22X1  AOI22X1_68
timestamp 1682952543
transform -1 0 1808 0 -1 3370
box -8 -3 46 105
use FILL  FILL_522
timestamp 1682952543
transform 1 0 1808 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_133
timestamp 1682952543
transform 1 0 1816 0 -1 3370
box -9 -3 26 105
use FILL  FILL_523
timestamp 1682952543
transform 1 0 1832 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2037
timestamp 1682952543
transform 1 0 1860 0 1 3275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_128
timestamp 1682952543
transform -1 0 1936 0 -1 3370
box -8 -3 104 105
use FILL  FILL_524
timestamp 1682952543
transform 1 0 1936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_525
timestamp 1682952543
transform 1 0 1944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_526
timestamp 1682952543
transform 1 0 1952 0 -1 3370
box -8 -3 16 105
use FILL  FILL_527
timestamp 1682952543
transform 1 0 1960 0 -1 3370
box -8 -3 16 105
use FILL  FILL_528
timestamp 1682952543
transform 1 0 1968 0 -1 3370
box -8 -3 16 105
use FILL  FILL_529
timestamp 1682952543
transform 1 0 1976 0 -1 3370
box -8 -3 16 105
use FILL  FILL_530
timestamp 1682952543
transform 1 0 1984 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_134
timestamp 1682952543
transform 1 0 1992 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_129
timestamp 1682952543
transform 1 0 2008 0 -1 3370
box -8 -3 104 105
use BUFX2  BUFX2_9
timestamp 1682952543
transform 1 0 2104 0 -1 3370
box -5 -3 28 105
use FILL  FILL_531
timestamp 1682952543
transform 1 0 2128 0 -1 3370
box -8 -3 16 105
use FILL  FILL_540
timestamp 1682952543
transform 1 0 2136 0 -1 3370
box -8 -3 16 105
use FILL  FILL_541
timestamp 1682952543
transform 1 0 2144 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_130
timestamp 1682952543
transform 1 0 2152 0 -1 3370
box -8 -3 104 105
use FILL  FILL_542
timestamp 1682952543
transform 1 0 2248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_544
timestamp 1682952543
transform 1 0 2256 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_137
timestamp 1682952543
transform 1 0 2264 0 -1 3370
box -8 -3 46 105
use FILL  FILL_579
timestamp 1682952543
transform 1 0 2304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_580
timestamp 1682952543
transform 1 0 2312 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_138
timestamp 1682952543
transform -1 0 2360 0 -1 3370
box -8 -3 46 105
use FILL  FILL_581
timestamp 1682952543
transform 1 0 2360 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_141
timestamp 1682952543
transform -1 0 2384 0 -1 3370
box -9 -3 26 105
use FILL  FILL_582
timestamp 1682952543
transform 1 0 2384 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1682952543
transform 1 0 2392 0 -1 3370
box -8 -3 104 105
use OAI22X1  OAI22X1_139
timestamp 1682952543
transform 1 0 2488 0 -1 3370
box -8 -3 46 105
use NAND2X1  NAND2X1_16
timestamp 1682952543
transform 1 0 2528 0 -1 3370
box -8 -3 32 105
use FILL  FILL_583
timestamp 1682952543
transform 1 0 2552 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_142
timestamp 1682952543
transform 1 0 2560 0 -1 3370
box -9 -3 26 105
use NAND2X1  NAND2X1_17
timestamp 1682952543
transform 1 0 2576 0 -1 3370
box -8 -3 32 105
use INVX2  INVX2_143
timestamp 1682952543
transform 1 0 2600 0 -1 3370
box -9 -3 26 105
use FILL  FILL_584
timestamp 1682952543
transform 1 0 2616 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_32
timestamp 1682952543
transform 1 0 2624 0 -1 3370
box -8 -3 34 105
use INVX2  INVX2_144
timestamp 1682952543
transform -1 0 2672 0 -1 3370
box -9 -3 26 105
use OAI21X1  OAI21X1_33
timestamp 1682952543
transform -1 0 2704 0 -1 3370
box -8 -3 34 105
use INVX2  INVX2_145
timestamp 1682952543
transform 1 0 2704 0 -1 3370
box -9 -3 26 105
use OAI21X1  OAI21X1_34
timestamp 1682952543
transform 1 0 2720 0 -1 3370
box -8 -3 34 105
use NAND2X1  NAND2X1_18
timestamp 1682952543
transform 1 0 2752 0 -1 3370
box -8 -3 32 105
use OAI21X1  OAI21X1_35
timestamp 1682952543
transform 1 0 2776 0 -1 3370
box -8 -3 34 105
use OAI22X1  OAI22X1_140
timestamp 1682952543
transform 1 0 2808 0 -1 3370
box -8 -3 46 105
use INVX2  INVX2_146
timestamp 1682952543
transform -1 0 2864 0 -1 3370
box -9 -3 26 105
use OAI22X1  OAI22X1_141
timestamp 1682952543
transform 1 0 2864 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_142
timestamp 1682952543
transform -1 0 2944 0 -1 3370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1682952543
transform 1 0 2944 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_147
timestamp 1682952543
transform 1 0 3040 0 -1 3370
box -9 -3 26 105
use FILL  FILL_585
timestamp 1682952543
transform 1 0 3056 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_143
timestamp 1682952543
transform -1 0 3104 0 -1 3370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1682952543
transform 1 0 3104 0 -1 3370
box -8 -3 104 105
use FILL  FILL_586
timestamp 1682952543
transform 1 0 3200 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_144
timestamp 1682952543
transform 1 0 3208 0 -1 3370
box -8 -3 46 105
use FILL  FILL_587
timestamp 1682952543
transform 1 0 3248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_589
timestamp 1682952543
transform 1 0 3256 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_149
timestamp 1682952543
transform 1 0 3264 0 -1 3370
box -9 -3 26 105
use FILL  FILL_592
timestamp 1682952543
transform 1 0 3280 0 -1 3370
box -8 -3 16 105
use FILL  FILL_593
timestamp 1682952543
transform 1 0 3288 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_153
timestamp 1682952543
transform 1 0 3296 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1682952543
transform 1 0 3312 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_154
timestamp 1682952543
transform 1 0 3408 0 -1 3370
box -9 -3 26 105
use OAI22X1  OAI22X1_147
timestamp 1682952543
transform 1 0 3424 0 -1 3370
box -8 -3 46 105
use AND2X2  AND2X2_1
timestamp 1682952543
transform -1 0 3496 0 -1 3370
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1682952543
transform -1 0 3528 0 -1 3370
box -8 -3 40 105
use M3_M2  M3_M2_2038
timestamp 1682952543
transform 1 0 3540 0 1 3275
box -3 -3 3 3
use M3_M2  M3_M2_2039
timestamp 1682952543
transform 1 0 3564 0 1 3275
box -3 -3 3 3
use AND2X2  AND2X2_3
timestamp 1682952543
transform 1 0 3528 0 -1 3370
box -8 -3 40 105
use FILL  FILL_611
timestamp 1682952543
transform 1 0 3560 0 -1 3370
box -8 -3 16 105
use FILL  FILL_612
timestamp 1682952543
transform 1 0 3568 0 -1 3370
box -8 -3 16 105
use FILL  FILL_613
timestamp 1682952543
transform 1 0 3576 0 -1 3370
box -8 -3 16 105
use FILL  FILL_614
timestamp 1682952543
transform 1 0 3584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_615
timestamp 1682952543
transform 1 0 3592 0 -1 3370
box -8 -3 16 105
use NAND2X1  NAND2X1_20
timestamp 1682952543
transform 1 0 3600 0 -1 3370
box -8 -3 32 105
use FILL  FILL_616
timestamp 1682952543
transform 1 0 3624 0 -1 3370
box -8 -3 16 105
use FILL  FILL_617
timestamp 1682952543
transform 1 0 3632 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_38
timestamp 1682952543
transform -1 0 3672 0 -1 3370
box -8 -3 34 105
use FILL  FILL_618
timestamp 1682952543
transform 1 0 3672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_620
timestamp 1682952543
transform 1 0 3680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_634
timestamp 1682952543
transform 1 0 3688 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2040
timestamp 1682952543
transform 1 0 3724 0 1 3275
box -3 -3 3 3
use OAI22X1  OAI22X1_152
timestamp 1682952543
transform 1 0 3696 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_153
timestamp 1682952543
transform 1 0 3736 0 -1 3370
box -8 -3 46 105
use INVX2  INVX2_155
timestamp 1682952543
transform -1 0 3792 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_136
timestamp 1682952543
transform 1 0 3792 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_156
timestamp 1682952543
transform -1 0 3904 0 -1 3370
box -9 -3 26 105
use OAI22X1  OAI22X1_154
timestamp 1682952543
transform 1 0 3904 0 -1 3370
box -8 -3 46 105
use OAI22X1  OAI22X1_155
timestamp 1682952543
transform 1 0 3944 0 -1 3370
box -8 -3 46 105
use M3_M2  M3_M2_2041
timestamp 1682952543
transform 1 0 4004 0 1 3275
box -3 -3 3 3
use INVX2  INVX2_157
timestamp 1682952543
transform -1 0 4000 0 -1 3370
box -9 -3 26 105
use FILL  FILL_635
timestamp 1682952543
transform 1 0 4000 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_157
timestamp 1682952543
transform 1 0 4008 0 -1 3370
box -8 -3 46 105
use M3_M2  M3_M2_2042
timestamp 1682952543
transform 1 0 4060 0 1 3275
box -3 -3 3 3
use FILL  FILL_645
timestamp 1682952543
transform 1 0 4048 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1682952543
transform 1 0 4056 0 -1 3370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_17
timestamp 1682952543
transform 1 0 4201 0 1 3270
box -10 -3 10 3
use M3_M2  M3_M2_2082
timestamp 1682952543
transform 1 0 164 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2110
timestamp 1682952543
transform 1 0 132 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2111
timestamp 1682952543
transform 1 0 172 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2120
timestamp 1682952543
transform 1 0 132 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2121
timestamp 1682952543
transform 1 0 164 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2122
timestamp 1682952543
transform 1 0 172 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1682952543
transform 1 0 84 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2193
timestamp 1682952543
transform 1 0 164 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2064
timestamp 1682952543
transform 1 0 220 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1682952543
transform 1 0 188 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2083
timestamp 1682952543
transform 1 0 236 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2113
timestamp 1682952543
transform 1 0 228 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2043
timestamp 1682952543
transform 1 0 284 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2044
timestamp 1682952543
transform 1 0 380 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2065
timestamp 1682952543
transform 1 0 364 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1682952543
transform 1 0 356 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2115
timestamp 1682952543
transform 1 0 388 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2123
timestamp 1682952543
transform 1 0 180 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2124
timestamp 1682952543
transform 1 0 204 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2125
timestamp 1682952543
transform 1 0 220 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1682952543
transform 1 0 228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2127
timestamp 1682952543
transform 1 0 244 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1682952543
transform 1 0 260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1682952543
transform 1 0 188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2250
timestamp 1682952543
transform 1 0 196 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1682952543
transform 1 0 212 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2194
timestamp 1682952543
transform 1 0 196 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1682952543
transform 1 0 188 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1682952543
transform 1 0 276 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2129
timestamp 1682952543
transform 1 0 300 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2147
timestamp 1682952543
transform 1 0 324 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2130
timestamp 1682952543
transform 1 0 356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1682952543
transform 1 0 364 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1682952543
transform 1 0 380 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1682952543
transform 1 0 396 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2252
timestamp 1682952543
transform 1 0 236 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1682952543
transform 1 0 252 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2169
timestamp 1682952543
transform 1 0 260 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2254
timestamp 1682952543
transform 1 0 276 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2170
timestamp 1682952543
transform 1 0 300 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2255
timestamp 1682952543
transform 1 0 364 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2256
timestamp 1682952543
transform 1 0 372 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2257
timestamp 1682952543
transform 1 0 388 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2227
timestamp 1682952543
transform 1 0 244 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2134
timestamp 1682952543
transform 1 0 420 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2066
timestamp 1682952543
transform 1 0 452 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2084
timestamp 1682952543
transform 1 0 468 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2135
timestamp 1682952543
transform 1 0 444 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1682952543
transform 1 0 460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2258
timestamp 1682952543
transform 1 0 452 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2259
timestamp 1682952543
transform 1 0 468 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2195
timestamp 1682952543
transform 1 0 468 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2228
timestamp 1682952543
transform 1 0 452 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2137
timestamp 1682952543
transform 1 0 484 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2055
timestamp 1682952543
transform 1 0 492 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_2138
timestamp 1682952543
transform 1 0 508 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2171
timestamp 1682952543
transform 1 0 508 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2045
timestamp 1682952543
transform 1 0 532 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_2139
timestamp 1682952543
transform 1 0 532 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2140
timestamp 1682952543
transform 1 0 548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2141
timestamp 1682952543
transform 1 0 564 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1682952543
transform 1 0 532 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1682952543
transform 1 0 540 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2196
timestamp 1682952543
transform 1 0 524 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2197
timestamp 1682952543
transform 1 0 540 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2262
timestamp 1682952543
transform 1 0 572 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2085
timestamp 1682952543
transform 1 0 588 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1682952543
transform 1 0 636 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1682952543
transform 1 0 612 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1682952543
transform 1 0 676 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1682952543
transform 1 0 676 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2142
timestamp 1682952543
transform 1 0 636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1682952543
transform 1 0 668 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1682952543
transform 1 0 676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2263
timestamp 1682952543
transform 1 0 588 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2198
timestamp 1682952543
transform 1 0 668 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1682952543
transform 1 0 708 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2145
timestamp 1682952543
transform 1 0 708 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2149
timestamp 1682952543
transform 1 0 716 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2146
timestamp 1682952543
transform 1 0 724 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1682952543
transform 1 0 708 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1682952543
transform 1 0 716 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1682952543
transform 1 0 732 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2199
timestamp 1682952543
transform 1 0 732 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1682952543
transform 1 0 780 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2267
timestamp 1682952543
transform 1 0 788 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2046
timestamp 1682952543
transform 1 0 820 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_2147
timestamp 1682952543
transform 1 0 804 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2150
timestamp 1682952543
transform 1 0 812 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2148
timestamp 1682952543
transform 1 0 820 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2151
timestamp 1682952543
transform 1 0 828 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2056
timestamp 1682952543
transform 1 0 844 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_2149
timestamp 1682952543
transform 1 0 844 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2268
timestamp 1682952543
transform 1 0 828 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1682952543
transform 1 0 836 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1682952543
transform 1 0 852 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2173
timestamp 1682952543
transform 1 0 876 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2347
timestamp 1682952543
transform 1 0 876 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_2270
timestamp 1682952543
transform 1 0 900 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2067
timestamp 1682952543
transform 1 0 916 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_2151
timestamp 1682952543
transform 1 0 924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1682952543
transform 1 0 924 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1682952543
transform 1 0 916 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1682952543
transform 1 0 940 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2229
timestamp 1682952543
transform 1 0 940 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1682952543
transform 1 0 964 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2152
timestamp 1682952543
transform 1 0 964 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2152
timestamp 1682952543
transform 1 0 972 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1682952543
transform 1 0 996 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2272
timestamp 1682952543
transform 1 0 988 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1682952543
transform 1 0 980 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1682952543
transform 1 0 1004 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1682952543
transform 1 0 1012 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2200
timestamp 1682952543
transform 1 0 1004 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2154
timestamp 1682952543
transform 1 0 1028 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1682952543
transform 1 0 1036 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2174
timestamp 1682952543
transform 1 0 1028 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2121
timestamp 1682952543
transform 1 0 1068 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2274
timestamp 1682952543
transform 1 0 1068 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2230
timestamp 1682952543
transform 1 0 1060 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2047
timestamp 1682952543
transform 1 0 1100 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1682952543
transform 1 0 1084 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1682952543
transform 1 0 1092 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2156
timestamp 1682952543
transform 1 0 1084 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1682952543
transform 1 0 1100 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2275
timestamp 1682952543
transform 1 0 1092 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2276
timestamp 1682952543
transform 1 0 1108 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2158
timestamp 1682952543
transform 1 0 1124 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1682952543
transform 1 0 1140 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2231
timestamp 1682952543
transform 1 0 1140 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1682952543
transform 1 0 1172 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2048
timestamp 1682952543
transform 1 0 1196 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2059
timestamp 1682952543
transform 1 0 1212 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2068
timestamp 1682952543
transform 1 0 1156 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1682952543
transform 1 0 1188 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2087
timestamp 1682952543
transform 1 0 1188 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1682952543
transform 1 0 1244 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1682952543
transform 1 0 1284 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2160
timestamp 1682952543
transform 1 0 1156 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2161
timestamp 1682952543
transform 1 0 1172 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1682952543
transform 1 0 1188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1682952543
transform 1 0 1244 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1682952543
transform 1 0 1284 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2175
timestamp 1682952543
transform 1 0 1156 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2277
timestamp 1682952543
transform 1 0 1164 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2278
timestamp 1682952543
transform 1 0 1268 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1682952543
transform 1 0 1308 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2070
timestamp 1682952543
transform 1 0 1348 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2088
timestamp 1682952543
transform 1 0 1324 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2166
timestamp 1682952543
transform 1 0 1332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2279
timestamp 1682952543
transform 1 0 1316 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1682952543
transform 1 0 1324 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1682952543
transform 1 0 1340 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2282
timestamp 1682952543
transform 1 0 1348 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2232
timestamp 1682952543
transform 1 0 1340 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1682952543
transform 1 0 1364 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2049
timestamp 1682952543
transform 1 0 1420 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2050
timestamp 1682952543
transform 1 0 1492 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1682952543
transform 1 0 1484 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2071
timestamp 1682952543
transform 1 0 1404 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1682952543
transform 1 0 1388 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1682952543
transform 1 0 1484 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2125
timestamp 1682952543
transform 1 0 1380 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1682952543
transform 1 0 1420 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2167
timestamp 1682952543
transform 1 0 1380 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1682952543
transform 1 0 1388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2169
timestamp 1682952543
transform 1 0 1420 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1682952543
transform 1 0 1372 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1682952543
transform 1 0 1468 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2285
timestamp 1682952543
transform 1 0 1484 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1682952543
transform 1 0 1508 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2051
timestamp 1682952543
transform 1 0 1548 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2092
timestamp 1682952543
transform 1 0 1548 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2127
timestamp 1682952543
transform 1 0 1532 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2171
timestamp 1682952543
transform 1 0 1532 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2153
timestamp 1682952543
transform 1 0 1540 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2172
timestamp 1682952543
transform 1 0 1548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1682952543
transform 1 0 1556 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1682952543
transform 1 0 1516 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1682952543
transform 1 0 1540 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2154
timestamp 1682952543
transform 1 0 1564 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1682952543
transform 1 0 1596 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1682952543
transform 1 0 1580 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2128
timestamp 1682952543
transform 1 0 1596 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2174
timestamp 1682952543
transform 1 0 1596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2288
timestamp 1682952543
transform 1 0 1564 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1682952543
transform 1 0 1572 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2176
timestamp 1682952543
transform 1 0 1580 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2290
timestamp 1682952543
transform 1 0 1588 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2201
timestamp 1682952543
transform 1 0 1588 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2175
timestamp 1682952543
transform 1 0 1612 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2052
timestamp 1682952543
transform 1 0 1660 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_2176
timestamp 1682952543
transform 1 0 1636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1682952543
transform 1 0 1660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1682952543
transform 1 0 1628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2292
timestamp 1682952543
transform 1 0 1644 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2293
timestamp 1682952543
transform 1 0 1652 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2202
timestamp 1682952543
transform 1 0 1612 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2233
timestamp 1682952543
transform 1 0 1604 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2352
timestamp 1682952543
transform 1 0 1612 0 1 3185
box -2 -2 2 2
use M3_M2  M3_M2_2234
timestamp 1682952543
transform 1 0 1620 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2235
timestamp 1682952543
transform 1 0 1644 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2129
timestamp 1682952543
transform 1 0 1676 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2094
timestamp 1682952543
transform 1 0 1740 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2130
timestamp 1682952543
transform 1 0 1716 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2178
timestamp 1682952543
transform 1 0 1676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1682952543
transform 1 0 1684 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2180
timestamp 1682952543
transform 1 0 1716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1682952543
transform 1 0 1764 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2236
timestamp 1682952543
transform 1 0 1684 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2181
timestamp 1682952543
transform 1 0 1780 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2203
timestamp 1682952543
transform 1 0 1780 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1682952543
transform 1 0 1820 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2182
timestamp 1682952543
transform 1 0 1804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2183
timestamp 1682952543
transform 1 0 1820 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2295
timestamp 1682952543
transform 1 0 1796 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2177
timestamp 1682952543
transform 1 0 1804 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2296
timestamp 1682952543
transform 1 0 1812 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2204
timestamp 1682952543
transform 1 0 1796 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1682952543
transform 1 0 1836 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1682952543
transform 1 0 1940 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1682952543
transform 1 0 1964 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1682952543
transform 1 0 1876 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1682952543
transform 1 0 1900 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1682952543
transform 1 0 1948 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1682952543
transform 1 0 1972 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2184
timestamp 1682952543
transform 1 0 1876 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1682952543
transform 1 0 1940 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2297
timestamp 1682952543
transform 1 0 1924 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2155
timestamp 1682952543
transform 1 0 1948 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2186
timestamp 1682952543
transform 1 0 1956 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2187
timestamp 1682952543
transform 1 0 1972 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2298
timestamp 1682952543
transform 1 0 1948 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2178
timestamp 1682952543
transform 1 0 1956 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2299
timestamp 1682952543
transform 1 0 1964 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2205
timestamp 1682952543
transform 1 0 1964 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2073
timestamp 1682952543
transform 1 0 2084 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1682952543
transform 1 0 2036 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2188
timestamp 1682952543
transform 1 0 1988 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2179
timestamp 1682952543
transform 1 0 1980 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1682952543
transform 1 0 1996 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2189
timestamp 1682952543
transform 1 0 2020 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2157
timestamp 1682952543
transform 1 0 2068 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2190
timestamp 1682952543
transform 1 0 2084 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2158
timestamp 1682952543
transform 1 0 2092 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2191
timestamp 1682952543
transform 1 0 2100 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2180
timestamp 1682952543
transform 1 0 2020 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2300
timestamp 1682952543
transform 1 0 2068 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2301
timestamp 1682952543
transform 1 0 2092 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2237
timestamp 1682952543
transform 1 0 2004 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1682952543
transform 1 0 2068 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2061
timestamp 1682952543
transform 1 0 2188 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2136
timestamp 1682952543
transform 1 0 2196 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2192
timestamp 1682952543
transform 1 0 2180 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2159
timestamp 1682952543
transform 1 0 2220 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2302
timestamp 1682952543
transform 1 0 2116 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2303
timestamp 1682952543
transform 1 0 2132 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2206
timestamp 1682952543
transform 1 0 2116 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2207
timestamp 1682952543
transform 1 0 2132 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2208
timestamp 1682952543
transform 1 0 2180 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2239
timestamp 1682952543
transform 1 0 2116 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2240
timestamp 1682952543
transform 1 0 2132 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2074
timestamp 1682952543
transform 1 0 2244 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1682952543
transform 1 0 2260 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2193
timestamp 1682952543
transform 1 0 2228 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2194
timestamp 1682952543
transform 1 0 2244 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2160
timestamp 1682952543
transform 1 0 2252 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1682952543
transform 1 0 2396 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1682952543
transform 1 0 2388 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2195
timestamp 1682952543
transform 1 0 2260 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1682952543
transform 1 0 2268 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1682952543
transform 1 0 2284 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1682952543
transform 1 0 2340 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1682952543
transform 1 0 2380 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1682952543
transform 1 0 2388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1682952543
transform 1 0 2444 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1682952543
transform 1 0 2236 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2181
timestamp 1682952543
transform 1 0 2244 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2305
timestamp 1682952543
transform 1 0 2252 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2306
timestamp 1682952543
transform 1 0 2276 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2209
timestamp 1682952543
transform 1 0 2252 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2182
timestamp 1682952543
transform 1 0 2284 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2307
timestamp 1682952543
transform 1 0 2300 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2241
timestamp 1682952543
transform 1 0 2300 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2308
timestamp 1682952543
transform 1 0 2468 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2210
timestamp 1682952543
transform 1 0 2468 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2113
timestamp 1682952543
transform 1 0 2676 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1682952543
transform 1 0 2516 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2203
timestamp 1682952543
transform 1 0 2572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1682952543
transform 1 0 2636 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1682952543
transform 1 0 2668 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1682952543
transform 1 0 2492 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2211
timestamp 1682952543
transform 1 0 2492 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2212
timestamp 1682952543
transform 1 0 2524 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2310
timestamp 1682952543
transform 1 0 2588 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2183
timestamp 1682952543
transform 1 0 2636 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2184
timestamp 1682952543
transform 1 0 2676 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2206
timestamp 1682952543
transform 1 0 2692 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1682952543
transform 1 0 2700 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2351
timestamp 1682952543
transform 1 0 2708 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2242
timestamp 1682952543
transform 1 0 2708 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2207
timestamp 1682952543
transform 1 0 2732 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2312
timestamp 1682952543
transform 1 0 2732 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2075
timestamp 1682952543
transform 1 0 2780 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1682952543
transform 1 0 2772 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1682952543
transform 1 0 2788 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1682952543
transform 1 0 2780 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2114
timestamp 1682952543
transform 1 0 2788 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2138
timestamp 1682952543
transform 1 0 2836 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1682952543
transform 1 0 2852 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1682952543
transform 1 0 2884 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2208
timestamp 1682952543
transform 1 0 2772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2209
timestamp 1682952543
transform 1 0 2780 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1682952543
transform 1 0 2748 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1682952543
transform 1 0 2772 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2243
timestamp 1682952543
transform 1 0 2748 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1682952543
transform 1 0 2788 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2210
timestamp 1682952543
transform 1 0 2852 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1682952543
transform 1 0 2884 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2212
timestamp 1682952543
transform 1 0 2892 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2315
timestamp 1682952543
transform 1 0 2804 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1682952543
transform 1 0 2892 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2213
timestamp 1682952543
transform 1 0 2804 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2115
timestamp 1682952543
transform 1 0 2916 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2162
timestamp 1682952543
transform 1 0 2916 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2213
timestamp 1682952543
transform 1 0 2924 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1682952543
transform 1 0 2980 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2317
timestamp 1682952543
transform 1 0 3020 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2214
timestamp 1682952543
transform 1 0 2956 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2215
timestamp 1682952543
transform 1 0 3084 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1682952543
transform 1 0 3044 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2185
timestamp 1682952543
transform 1 0 3092 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2215
timestamp 1682952543
transform 1 0 3044 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2076
timestamp 1682952543
transform 1 0 3148 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_2116
timestamp 1682952543
transform 1 0 3148 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1682952543
transform 1 0 3140 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2163
timestamp 1682952543
transform 1 0 3148 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2217
timestamp 1682952543
transform 1 0 3156 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1682952543
transform 1 0 3164 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1682952543
transform 1 0 3188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1682952543
transform 1 0 3204 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2186
timestamp 1682952543
transform 1 0 3140 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2319
timestamp 1682952543
transform 1 0 3164 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2164
timestamp 1682952543
transform 1 0 3212 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2221
timestamp 1682952543
transform 1 0 3220 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2320
timestamp 1682952543
transform 1 0 3196 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2216
timestamp 1682952543
transform 1 0 3188 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2321
timestamp 1682952543
transform 1 0 3228 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2322
timestamp 1682952543
transform 1 0 3236 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2244
timestamp 1682952543
transform 1 0 3220 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1682952543
transform 1 0 3236 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2323
timestamp 1682952543
transform 1 0 3260 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2217
timestamp 1682952543
transform 1 0 3260 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1682952543
transform 1 0 3276 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1682952543
transform 1 0 3316 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1682952543
transform 1 0 3332 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2222
timestamp 1682952543
transform 1 0 3276 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1682952543
transform 1 0 3292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1682952543
transform 1 0 3300 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2225
timestamp 1682952543
transform 1 0 3316 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1682952543
transform 1 0 3332 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2324
timestamp 1682952543
transform 1 0 3324 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2325
timestamp 1682952543
transform 1 0 3332 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2246
timestamp 1682952543
transform 1 0 3324 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2187
timestamp 1682952543
transform 1 0 3348 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2227
timestamp 1682952543
transform 1 0 3388 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1682952543
transform 1 0 3364 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2077
timestamp 1682952543
transform 1 0 3468 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_2117
timestamp 1682952543
transform 1 0 3468 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_2228
timestamp 1682952543
transform 1 0 3460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1682952543
transform 1 0 3468 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2078
timestamp 1682952543
transform 1 0 3492 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1682952543
transform 1 0 3500 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2118
timestamp 1682952543
transform 1 0 3492 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2218
timestamp 1682952543
transform 1 0 3468 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1682952543
transform 1 0 3484 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2229
timestamp 1682952543
transform 1 0 3500 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2188
timestamp 1682952543
transform 1 0 3500 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2230
timestamp 1682952543
transform 1 0 3516 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2104
timestamp 1682952543
transform 1 0 3556 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2231
timestamp 1682952543
transform 1 0 3556 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1682952543
transform 1 0 3540 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2329
timestamp 1682952543
transform 1 0 3548 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2189
timestamp 1682952543
transform 1 0 3556 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2330
timestamp 1682952543
transform 1 0 3564 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1682952543
transform 1 0 3580 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2247
timestamp 1682952543
transform 1 0 3540 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2220
timestamp 1682952543
transform 1 0 3580 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2232
timestamp 1682952543
transform 1 0 3596 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2248
timestamp 1682952543
transform 1 0 3604 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2332
timestamp 1682952543
transform 1 0 3620 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2221
timestamp 1682952543
transform 1 0 3620 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2333
timestamp 1682952543
transform 1 0 3660 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2105
timestamp 1682952543
transform 1 0 3708 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2165
timestamp 1682952543
transform 1 0 3684 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2233
timestamp 1682952543
transform 1 0 3692 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2234
timestamp 1682952543
transform 1 0 3708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2334
timestamp 1682952543
transform 1 0 3684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2335
timestamp 1682952543
transform 1 0 3700 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2079
timestamp 1682952543
transform 1 0 3764 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1682952543
transform 1 0 3748 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2235
timestamp 1682952543
transform 1 0 3740 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1682952543
transform 1 0 3748 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2237
timestamp 1682952543
transform 1 0 3764 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1682952543
transform 1 0 3732 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2249
timestamp 1682952543
transform 1 0 3732 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2337
timestamp 1682952543
transform 1 0 3756 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2190
timestamp 1682952543
transform 1 0 3764 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2053
timestamp 1682952543
transform 1 0 3868 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1682952543
transform 1 0 3780 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2338
timestamp 1682952543
transform 1 0 3772 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2222
timestamp 1682952543
transform 1 0 3756 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2238
timestamp 1682952543
transform 1 0 3788 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2239
timestamp 1682952543
transform 1 0 3820 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2339
timestamp 1682952543
transform 1 0 3868 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2223
timestamp 1682952543
transform 1 0 3820 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2224
timestamp 1682952543
transform 1 0 3868 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1682952543
transform 1 0 3844 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2080
timestamp 1682952543
transform 1 0 3916 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2108
timestamp 1682952543
transform 1 0 3924 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2144
timestamp 1682952543
transform 1 0 3908 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1682952543
transform 1 0 3892 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2240
timestamp 1682952543
transform 1 0 3900 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2167
timestamp 1682952543
transform 1 0 3908 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2241
timestamp 1682952543
transform 1 0 3916 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2168
timestamp 1682952543
transform 1 0 3924 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_2242
timestamp 1682952543
transform 1 0 3932 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2191
timestamp 1682952543
transform 1 0 3884 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2340
timestamp 1682952543
transform 1 0 3892 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2192
timestamp 1682952543
transform 1 0 3900 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_2341
timestamp 1682952543
transform 1 0 3908 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_2342
timestamp 1682952543
transform 1 0 3924 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2251
timestamp 1682952543
transform 1 0 3924 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_2243
timestamp 1682952543
transform 1 0 3940 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2145
timestamp 1682952543
transform 1 0 3948 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_2343
timestamp 1682952543
transform 1 0 3956 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2109
timestamp 1682952543
transform 1 0 4004 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_2244
timestamp 1682952543
transform 1 0 4004 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1682952543
transform 1 0 4060 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2246
timestamp 1682952543
transform 1 0 4068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_2344
timestamp 1682952543
transform 1 0 3980 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2225
timestamp 1682952543
transform 1 0 3980 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_2345
timestamp 1682952543
transform 1 0 4068 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2063
timestamp 1682952543
transform 1 0 4092 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2081
timestamp 1682952543
transform 1 0 4108 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_2119
timestamp 1682952543
transform 1 0 4092 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_2247
timestamp 1682952543
transform 1 0 4108 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2054
timestamp 1682952543
transform 1 0 4156 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_2346
timestamp 1682952543
transform 1 0 4148 0 1 3205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_18
timestamp 1682952543
transform 1 0 48 0 1 3170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_138
timestamp 1682952543
transform 1 0 72 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_160
timestamp 1682952543
transform -1 0 184 0 1 3170
box -9 -3 26 105
use M3_M2  M3_M2_2252
timestamp 1682952543
transform 1 0 212 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_69
timestamp 1682952543
transform -1 0 224 0 1 3170
box -8 -3 46 105
use M3_M2  M3_M2_2253
timestamp 1682952543
transform 1 0 252 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_70
timestamp 1682952543
transform -1 0 264 0 1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1682952543
transform 1 0 264 0 1 3170
box -8 -3 104 105
use AOI22X1  AOI22X1_71
timestamp 1682952543
transform 1 0 360 0 1 3170
box -8 -3 46 105
use FILL  FILL_646
timestamp 1682952543
transform 1 0 400 0 1 3170
box -8 -3 16 105
use FILL  FILL_647
timestamp 1682952543
transform 1 0 408 0 1 3170
box -8 -3 16 105
use FILL  FILL_648
timestamp 1682952543
transform 1 0 416 0 1 3170
box -8 -3 16 105
use FILL  FILL_649
timestamp 1682952543
transform 1 0 424 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_158
timestamp 1682952543
transform 1 0 432 0 1 3170
box -8 -3 46 105
use FILL  FILL_650
timestamp 1682952543
transform 1 0 472 0 1 3170
box -8 -3 16 105
use FILL  FILL_651
timestamp 1682952543
transform 1 0 480 0 1 3170
box -8 -3 16 105
use FILL  FILL_652
timestamp 1682952543
transform 1 0 488 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_162
timestamp 1682952543
transform -1 0 512 0 1 3170
box -9 -3 26 105
use FILL  FILL_653
timestamp 1682952543
transform 1 0 512 0 1 3170
box -8 -3 16 105
use FILL  FILL_654
timestamp 1682952543
transform 1 0 520 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_72
timestamp 1682952543
transform 1 0 528 0 1 3170
box -8 -3 46 105
use FILL  FILL_657
timestamp 1682952543
transform 1 0 568 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_143
timestamp 1682952543
transform 1 0 576 0 1 3170
box -8 -3 104 105
use FILL  FILL_658
timestamp 1682952543
transform 1 0 672 0 1 3170
box -8 -3 16 105
use FILL  FILL_659
timestamp 1682952543
transform 1 0 680 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_164
timestamp 1682952543
transform -1 0 704 0 1 3170
box -9 -3 26 105
use M3_M2  M3_M2_2254
timestamp 1682952543
transform 1 0 748 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_76
timestamp 1682952543
transform 1 0 704 0 1 3170
box -8 -3 46 105
use FILL  FILL_660
timestamp 1682952543
transform 1 0 744 0 1 3170
box -8 -3 16 105
use FILL  FILL_665
timestamp 1682952543
transform 1 0 752 0 1 3170
box -8 -3 16 105
use FILL  FILL_666
timestamp 1682952543
transform 1 0 760 0 1 3170
box -8 -3 16 105
use FILL  FILL_667
timestamp 1682952543
transform 1 0 768 0 1 3170
box -8 -3 16 105
use FILL  FILL_668
timestamp 1682952543
transform 1 0 776 0 1 3170
box -8 -3 16 105
use FILL  FILL_669
timestamp 1682952543
transform 1 0 784 0 1 3170
box -8 -3 16 105
use FILL  FILL_670
timestamp 1682952543
transform 1 0 792 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_77
timestamp 1682952543
transform -1 0 840 0 1 3170
box -8 -3 46 105
use FILL  FILL_671
timestamp 1682952543
transform 1 0 840 0 1 3170
box -8 -3 16 105
use FILL  FILL_672
timestamp 1682952543
transform 1 0 848 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_166
timestamp 1682952543
transform 1 0 856 0 1 3170
box -9 -3 26 105
use FILL  FILL_673
timestamp 1682952543
transform 1 0 872 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2255
timestamp 1682952543
transform 1 0 892 0 1 3175
box -3 -3 3 3
use FILL  FILL_674
timestamp 1682952543
transform 1 0 880 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_16
timestamp 1682952543
transform 1 0 888 0 1 3170
box -8 -3 32 105
use FILL  FILL_675
timestamp 1682952543
transform 1 0 912 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_17
timestamp 1682952543
transform 1 0 920 0 1 3170
box -8 -3 32 105
use FILL  FILL_678
timestamp 1682952543
transform 1 0 944 0 1 3170
box -8 -3 16 105
use FILL  FILL_680
timestamp 1682952543
transform 1 0 952 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_19
timestamp 1682952543
transform 1 0 960 0 1 3170
box -8 -3 32 105
use FILL  FILL_681
timestamp 1682952543
transform 1 0 984 0 1 3170
box -8 -3 16 105
use FILL  FILL_682
timestamp 1682952543
transform 1 0 992 0 1 3170
box -8 -3 16 105
use FILL  FILL_683
timestamp 1682952543
transform 1 0 1000 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_20
timestamp 1682952543
transform 1 0 1008 0 1 3170
box -8 -3 32 105
use FILL  FILL_684
timestamp 1682952543
transform 1 0 1032 0 1 3170
box -8 -3 16 105
use FILL  FILL_685
timestamp 1682952543
transform 1 0 1040 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_168
timestamp 1682952543
transform -1 0 1064 0 1 3170
box -9 -3 26 105
use FILL  FILL_686
timestamp 1682952543
transform 1 0 1064 0 1 3170
box -8 -3 16 105
use FILL  FILL_687
timestamp 1682952543
transform 1 0 1072 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_78
timestamp 1682952543
transform 1 0 1080 0 1 3170
box -8 -3 46 105
use FILL  FILL_690
timestamp 1682952543
transform 1 0 1120 0 1 3170
box -8 -3 16 105
use FILL  FILL_691
timestamp 1682952543
transform 1 0 1128 0 1 3170
box -8 -3 16 105
use FILL  FILL_694
timestamp 1682952543
transform 1 0 1136 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2256
timestamp 1682952543
transform 1 0 1156 0 1 3175
box -3 -3 3 3
use OAI22X1  OAI22X1_162
timestamp 1682952543
transform -1 0 1184 0 1 3170
box -8 -3 46 105
use M3_M2  M3_M2_2257
timestamp 1682952543
transform 1 0 1236 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_147
timestamp 1682952543
transform -1 0 1280 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_170
timestamp 1682952543
transform -1 0 1296 0 1 3170
box -9 -3 26 105
use FILL  FILL_695
timestamp 1682952543
transform 1 0 1296 0 1 3170
box -8 -3 16 105
use FILL  FILL_696
timestamp 1682952543
transform 1 0 1304 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_80
timestamp 1682952543
transform -1 0 1352 0 1 3170
box -8 -3 46 105
use FILL  FILL_697
timestamp 1682952543
transform 1 0 1352 0 1 3170
box -8 -3 16 105
use FILL  FILL_704
timestamp 1682952543
transform 1 0 1360 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_171
timestamp 1682952543
transform 1 0 1368 0 1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_149
timestamp 1682952543
transform -1 0 1480 0 1 3170
box -8 -3 104 105
use FILL  FILL_706
timestamp 1682952543
transform 1 0 1480 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_11
timestamp 1682952543
transform -1 0 1512 0 1 3170
box -5 -3 28 105
use FILL  FILL_707
timestamp 1682952543
transform 1 0 1512 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_164
timestamp 1682952543
transform -1 0 1560 0 1 3170
box -8 -3 46 105
use FILL  FILL_708
timestamp 1682952543
transform 1 0 1560 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_165
timestamp 1682952543
transform 1 0 1568 0 1 3170
box -8 -3 46 105
use FILL  FILL_709
timestamp 1682952543
transform 1 0 1608 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_82
timestamp 1682952543
transform 1 0 1616 0 1 3170
box -8 -3 46 105
use INVX2  INVX2_173
timestamp 1682952543
transform 1 0 1656 0 1 3170
box -9 -3 26 105
use FILL  FILL_710
timestamp 1682952543
transform 1 0 1672 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_152
timestamp 1682952543
transform -1 0 1776 0 1 3170
box -8 -3 104 105
use FILL  FILL_711
timestamp 1682952543
transform 1 0 1776 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_84
timestamp 1682952543
transform 1 0 1784 0 1 3170
box -8 -3 46 105
use FILL  FILL_712
timestamp 1682952543
transform 1 0 1824 0 1 3170
box -8 -3 16 105
use FILL  FILL_713
timestamp 1682952543
transform 1 0 1832 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_153
timestamp 1682952543
transform -1 0 1936 0 1 3170
box -8 -3 104 105
use AOI22X1  AOI22X1_85
timestamp 1682952543
transform -1 0 1976 0 1 3170
box -8 -3 46 105
use FILL  FILL_714
timestamp 1682952543
transform 1 0 1976 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2258
timestamp 1682952543
transform 1 0 2036 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2259
timestamp 1682952543
transform 1 0 2060 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2260
timestamp 1682952543
transform 1 0 2076 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_154
timestamp 1682952543
transform -1 0 2080 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_175
timestamp 1682952543
transform -1 0 2096 0 1 3170
box -9 -3 26 105
use M3_M2  M3_M2_2261
timestamp 1682952543
transform 1 0 2108 0 1 3175
box -3 -3 3 3
use BUFX2  BUFX2_12
timestamp 1682952543
transform 1 0 2096 0 1 3170
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_155
timestamp 1682952543
transform 1 0 2120 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_176
timestamp 1682952543
transform 1 0 2216 0 1 3170
box -9 -3 26 105
use OAI22X1  OAI22X1_167
timestamp 1682952543
transform -1 0 2272 0 1 3170
box -8 -3 46 105
use INVX2  INVX2_177
timestamp 1682952543
transform 1 0 2272 0 1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_156
timestamp 1682952543
transform 1 0 2288 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_157
timestamp 1682952543
transform -1 0 2480 0 1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2262
timestamp 1682952543
transform 1 0 2524 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_158
timestamp 1682952543
transform 1 0 2480 0 1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2263
timestamp 1682952543
transform 1 0 2588 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2264
timestamp 1682952543
transform 1 0 2628 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_159
timestamp 1682952543
transform 1 0 2576 0 1 3170
box -8 -3 104 105
use FILL  FILL_715
timestamp 1682952543
transform 1 0 2672 0 1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_22
timestamp 1682952543
transform -1 0 2704 0 1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_21
timestamp 1682952543
transform 1 0 2704 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_23
timestamp 1682952543
transform 1 0 2728 0 1 3170
box -8 -3 32 105
use INVX2  INVX2_178
timestamp 1682952543
transform 1 0 2752 0 1 3170
box -9 -3 26 105
use NAND2X1  NAND2X1_24
timestamp 1682952543
transform 1 0 2768 0 1 3170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_160
timestamp 1682952543
transform 1 0 2792 0 1 3170
box -8 -3 104 105
use NAND2X1  NAND2X1_25
timestamp 1682952543
transform 1 0 2888 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_26
timestamp 1682952543
transform -1 0 2936 0 1 3170
box -8 -3 32 105
use M3_M2  M3_M2_2265
timestamp 1682952543
transform 1 0 3020 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_161
timestamp 1682952543
transform -1 0 3032 0 1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_162
timestamp 1682952543
transform 1 0 3032 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_179
timestamp 1682952543
transform 1 0 3128 0 1 3170
box -9 -3 26 105
use NAND2X1  NAND2X1_27
timestamp 1682952543
transform -1 0 3168 0 1 3170
box -8 -3 32 105
use AND2X2  AND2X2_4
timestamp 1682952543
transform -1 0 3200 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_5
timestamp 1682952543
transform -1 0 3232 0 1 3170
box -8 -3 40 105
use INVX2  INVX2_180
timestamp 1682952543
transform 1 0 3232 0 1 3170
box -9 -3 26 105
use FILL  FILL_716
timestamp 1682952543
transform 1 0 3248 0 1 3170
box -8 -3 16 105
use FILL  FILL_746
timestamp 1682952543
transform 1 0 3256 0 1 3170
box -8 -3 16 105
use AND2X2  AND2X2_7
timestamp 1682952543
transform 1 0 3264 0 1 3170
box -8 -3 40 105
use AND2X2  AND2X2_8
timestamp 1682952543
transform -1 0 3328 0 1 3170
box -8 -3 40 105
use INVX2  INVX2_183
timestamp 1682952543
transform 1 0 3328 0 1 3170
box -9 -3 26 105
use FILL  FILL_748
timestamp 1682952543
transform 1 0 3344 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2266
timestamp 1682952543
transform 1 0 3364 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1682952543
transform 1 0 3404 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_172
timestamp 1682952543
transform 1 0 3352 0 1 3170
box -8 -3 104 105
use NAND2X1  NAND2X1_29
timestamp 1682952543
transform 1 0 3448 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_30
timestamp 1682952543
transform 1 0 3472 0 1 3170
box -8 -3 32 105
use FILL  FILL_749
timestamp 1682952543
transform 1 0 3496 0 1 3170
box -8 -3 16 105
use FILL  FILL_750
timestamp 1682952543
transform 1 0 3504 0 1 3170
box -8 -3 16 105
use FILL  FILL_751
timestamp 1682952543
transform 1 0 3512 0 1 3170
box -8 -3 16 105
use FILL  FILL_752
timestamp 1682952543
transform 1 0 3520 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_184
timestamp 1682952543
transform -1 0 3544 0 1 3170
box -9 -3 26 105
use OAI22X1  OAI22X1_168
timestamp 1682952543
transform -1 0 3584 0 1 3170
box -8 -3 46 105
use FILL  FILL_753
timestamp 1682952543
transform 1 0 3584 0 1 3170
box -8 -3 16 105
use FILL  FILL_754
timestamp 1682952543
transform 1 0 3592 0 1 3170
box -8 -3 16 105
use FILL  FILL_755
timestamp 1682952543
transform 1 0 3600 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_185
timestamp 1682952543
transform -1 0 3624 0 1 3170
box -9 -3 26 105
use FILL  FILL_756
timestamp 1682952543
transform 1 0 3624 0 1 3170
box -8 -3 16 105
use FILL  FILL_757
timestamp 1682952543
transform 1 0 3632 0 1 3170
box -8 -3 16 105
use FILL  FILL_758
timestamp 1682952543
transform 1 0 3640 0 1 3170
box -8 -3 16 105
use FILL  FILL_759
timestamp 1682952543
transform 1 0 3648 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_186
timestamp 1682952543
transform 1 0 3656 0 1 3170
box -9 -3 26 105
use FILL  FILL_760
timestamp 1682952543
transform 1 0 3672 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_169
timestamp 1682952543
transform 1 0 3680 0 1 3170
box -8 -3 46 105
use FILL  FILL_761
timestamp 1682952543
transform 1 0 3720 0 1 3170
box -8 -3 16 105
use FILL  FILL_762
timestamp 1682952543
transform 1 0 3728 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_170
timestamp 1682952543
transform 1 0 3736 0 1 3170
box -8 -3 46 105
use FILL  FILL_763
timestamp 1682952543
transform 1 0 3776 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_173
timestamp 1682952543
transform -1 0 3880 0 1 3170
box -8 -3 104 105
use FILL  FILL_764
timestamp 1682952543
transform 1 0 3880 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_171
timestamp 1682952543
transform 1 0 3888 0 1 3170
box -8 -3 46 105
use FILL  FILL_765
timestamp 1682952543
transform 1 0 3928 0 1 3170
box -8 -3 16 105
use FILL  FILL_766
timestamp 1682952543
transform 1 0 3936 0 1 3170
box -8 -3 16 105
use FILL  FILL_767
timestamp 1682952543
transform 1 0 3944 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_187
timestamp 1682952543
transform 1 0 3952 0 1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_174
timestamp 1682952543
transform 1 0 3968 0 1 3170
box -8 -3 104 105
use FILL  FILL_768
timestamp 1682952543
transform 1 0 4064 0 1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_31
timestamp 1682952543
transform 1 0 4072 0 1 3170
box -8 -3 32 105
use NAND2X1  NAND2X1_32
timestamp 1682952543
transform -1 0 4120 0 1 3170
box -8 -3 32 105
use FILL  FILL_769
timestamp 1682952543
transform 1 0 4120 0 1 3170
box -8 -3 16 105
use FILL  FILL_770
timestamp 1682952543
transform 1 0 4128 0 1 3170
box -8 -3 16 105
use FILL  FILL_771
timestamp 1682952543
transform 1 0 4136 0 1 3170
box -8 -3 16 105
use FILL  FILL_772
timestamp 1682952543
transform 1 0 4144 0 1 3170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_19
timestamp 1682952543
transform 1 0 4177 0 1 3170
box -10 -3 10 3
use M3_M2  M3_M2_2305
timestamp 1682952543
transform 1 0 84 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2360
timestamp 1682952543
transform 1 0 84 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2362
timestamp 1682952543
transform 1 0 84 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1682952543
transform 1 0 116 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_2439
timestamp 1682952543
transform 1 0 132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1682952543
transform 1 0 164 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1682952543
transform 1 0 172 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2374
timestamp 1682952543
transform 1 0 84 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1682952543
transform 1 0 132 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2376
timestamp 1682952543
transform 1 0 172 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1682952543
transform 1 0 196 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2361
timestamp 1682952543
transform 1 0 188 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1682952543
transform 1 0 196 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1682952543
transform 1 0 212 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2307
timestamp 1682952543
transform 1 0 316 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2364
timestamp 1682952543
transform 1 0 236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1682952543
transform 1 0 324 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1682952543
transform 1 0 188 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1682952543
transform 1 0 204 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2444
timestamp 1682952543
transform 1 0 220 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2377
timestamp 1682952543
transform 1 0 196 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2378
timestamp 1682952543
transform 1 0 212 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2364
timestamp 1682952543
transform 1 0 236 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_2366
timestamp 1682952543
transform 1 0 348 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2280
timestamp 1682952543
transform 1 0 388 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2308
timestamp 1682952543
transform 1 0 380 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2367
timestamp 1682952543
transform 1 0 380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1682952543
transform 1 0 260 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1682952543
transform 1 0 316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1682952543
transform 1 0 332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1682952543
transform 1 0 340 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1682952543
transform 1 0 356 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2450
timestamp 1682952543
transform 1 0 372 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2379
timestamp 1682952543
transform 1 0 324 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1682952543
transform 1 0 228 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2422
timestamp 1682952543
transform 1 0 260 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2442
timestamp 1682952543
transform 1 0 220 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1682952543
transform 1 0 356 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2443
timestamp 1682952543
transform 1 0 340 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_2368
timestamp 1682952543
transform 1 0 388 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1682952543
transform 1 0 388 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2281
timestamp 1682952543
transform 1 0 444 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2282
timestamp 1682952543
transform 1 0 516 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1682952543
transform 1 0 428 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2310
timestamp 1682952543
transform 1 0 556 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2369
timestamp 1682952543
transform 1 0 412 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2370
timestamp 1682952543
transform 1 0 428 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1682952543
transform 1 0 444 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1682952543
transform 1 0 532 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1682952543
transform 1 0 556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1682952543
transform 1 0 404 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1682952543
transform 1 0 420 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2381
timestamp 1682952543
transform 1 0 404 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_2454
timestamp 1682952543
transform 1 0 484 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2455
timestamp 1682952543
transform 1 0 524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2456
timestamp 1682952543
transform 1 0 532 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2365
timestamp 1682952543
transform 1 0 540 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2283
timestamp 1682952543
transform 1 0 580 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2374
timestamp 1682952543
transform 1 0 580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1682952543
transform 1 0 668 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1682952543
transform 1 0 548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1682952543
transform 1 0 564 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2459
timestamp 1682952543
transform 1 0 628 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2460
timestamp 1682952543
transform 1 0 660 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1682952543
transform 1 0 668 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2382
timestamp 1682952543
transform 1 0 476 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2383
timestamp 1682952543
transform 1 0 524 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2384
timestamp 1682952543
transform 1 0 556 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2423
timestamp 1682952543
transform 1 0 492 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1682952543
transform 1 0 532 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1682952543
transform 1 0 516 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2385
timestamp 1682952543
transform 1 0 628 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1682952543
transform 1 0 668 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2425
timestamp 1682952543
transform 1 0 628 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2445
timestamp 1682952543
transform 1 0 612 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_2376
timestamp 1682952543
transform 1 0 684 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2366
timestamp 1682952543
transform 1 0 684 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2426
timestamp 1682952543
transform 1 0 676 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1682952543
transform 1 0 692 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2284
timestamp 1682952543
transform 1 0 716 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1682952543
transform 1 0 740 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2377
timestamp 1682952543
transform 1 0 716 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2378
timestamp 1682952543
transform 1 0 732 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1682952543
transform 1 0 740 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1682952543
transform 1 0 708 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2463
timestamp 1682952543
transform 1 0 724 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2387
timestamp 1682952543
transform 1 0 708 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2427
timestamp 1682952543
transform 1 0 724 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_2464
timestamp 1682952543
transform 1 0 740 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2388
timestamp 1682952543
transform 1 0 740 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1682952543
transform 1 0 772 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_2380
timestamp 1682952543
transform 1 0 772 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1682952543
transform 1 0 788 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2465
timestamp 1682952543
transform 1 0 756 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2466
timestamp 1682952543
transform 1 0 780 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2389
timestamp 1682952543
transform 1 0 780 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2428
timestamp 1682952543
transform 1 0 772 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1682952543
transform 1 0 844 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2313
timestamp 1682952543
transform 1 0 884 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2382
timestamp 1682952543
transform 1 0 884 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1682952543
transform 1 0 852 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2468
timestamp 1682952543
transform 1 0 900 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2390
timestamp 1682952543
transform 1 0 900 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2447
timestamp 1682952543
transform 1 0 884 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2285
timestamp 1682952543
transform 1 0 916 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2353
timestamp 1682952543
transform 1 0 916 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1682952543
transform 1 0 916 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2367
timestamp 1682952543
transform 1 0 916 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_2384
timestamp 1682952543
transform 1 0 932 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2314
timestamp 1682952543
transform 1 0 948 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2469
timestamp 1682952543
transform 1 0 948 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2269
timestamp 1682952543
transform 1 0 980 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_2385
timestamp 1682952543
transform 1 0 964 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2339
timestamp 1682952543
transform 1 0 1036 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2470
timestamp 1682952543
transform 1 0 1004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1682952543
transform 1 0 1044 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2391
timestamp 1682952543
transform 1 0 1004 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2429
timestamp 1682952543
transform 1 0 996 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2286
timestamp 1682952543
transform 1 0 1068 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2472
timestamp 1682952543
transform 1 0 1060 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2392
timestamp 1682952543
transform 1 0 1060 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1682952543
transform 1 0 1084 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2287
timestamp 1682952543
transform 1 0 1092 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2386
timestamp 1682952543
transform 1 0 1084 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1682952543
transform 1 0 1092 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2340
timestamp 1682952543
transform 1 0 1108 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2388
timestamp 1682952543
transform 1 0 1116 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2473
timestamp 1682952543
transform 1 0 1092 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1682952543
transform 1 0 1108 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2475
timestamp 1682952543
transform 1 0 1124 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2393
timestamp 1682952543
transform 1 0 1084 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2394
timestamp 1682952543
transform 1 0 1108 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2456
timestamp 1682952543
transform 1 0 1092 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1682952543
transform 1 0 1180 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2389
timestamp 1682952543
transform 1 0 1180 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2476
timestamp 1682952543
transform 1 0 1172 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2477
timestamp 1682952543
transform 1 0 1188 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2316
timestamp 1682952543
transform 1 0 1212 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2390
timestamp 1682952543
transform 1 0 1212 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2288
timestamp 1682952543
transform 1 0 1228 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2289
timestamp 1682952543
transform 1 0 1268 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1682952543
transform 1 0 1340 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1682952543
transform 1 0 1316 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2391
timestamp 1682952543
transform 1 0 1228 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1682952543
transform 1 0 1316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1682952543
transform 1 0 1340 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1682952543
transform 1 0 1348 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1682952543
transform 1 0 1356 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2478
timestamp 1682952543
transform 1 0 1252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1682952543
transform 1 0 1308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1682952543
transform 1 0 1316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2481
timestamp 1682952543
transform 1 0 1332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2482
timestamp 1682952543
transform 1 0 1348 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2430
timestamp 1682952543
transform 1 0 1220 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2395
timestamp 1682952543
transform 1 0 1332 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2448
timestamp 1682952543
transform 1 0 1340 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2457
timestamp 1682952543
transform 1 0 1340 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2396
timestamp 1682952543
transform 1 0 1356 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1682952543
transform 1 0 1436 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1682952543
transform 1 0 1468 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2290
timestamp 1682952543
transform 1 0 1468 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1682952543
transform 1 0 1388 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2396
timestamp 1682952543
transform 1 0 1468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2483
timestamp 1682952543
transform 1 0 1380 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1682952543
transform 1 0 1388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2485
timestamp 1682952543
transform 1 0 1420 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2397
timestamp 1682952543
transform 1 0 1380 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2398
timestamp 1682952543
transform 1 0 1420 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2291
timestamp 1682952543
transform 1 0 1620 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2292
timestamp 1682952543
transform 1 0 1644 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2397
timestamp 1682952543
transform 1 0 1492 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2398
timestamp 1682952543
transform 1 0 1580 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2341
timestamp 1682952543
transform 1 0 1588 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1682952543
transform 1 0 1636 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1682952543
transform 1 0 1652 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2399
timestamp 1682952543
transform 1 0 1596 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2400
timestamp 1682952543
transform 1 0 1620 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1682952543
transform 1 0 1628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1682952543
transform 1 0 1644 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1682952543
transform 1 0 1652 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1682952543
transform 1 0 1516 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2487
timestamp 1682952543
transform 1 0 1572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2488
timestamp 1682952543
transform 1 0 1580 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2489
timestamp 1682952543
transform 1 0 1604 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2490
timestamp 1682952543
transform 1 0 1620 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2491
timestamp 1682952543
transform 1 0 1636 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2492
timestamp 1682952543
transform 1 0 1652 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2399
timestamp 1682952543
transform 1 0 1556 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1682952543
transform 1 0 1580 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2431
timestamp 1682952543
transform 1 0 1436 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2432
timestamp 1682952543
transform 1 0 1484 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2458
timestamp 1682952543
transform 1 0 1460 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2459
timestamp 1682952543
transform 1 0 1524 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2449
timestamp 1682952543
transform 1 0 1620 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2293
timestamp 1682952543
transform 1 0 1692 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2404
timestamp 1682952543
transform 1 0 1772 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1682952543
transform 1 0 1684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2494
timestamp 1682952543
transform 1 0 1692 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2495
timestamp 1682952543
transform 1 0 1724 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2401
timestamp 1682952543
transform 1 0 1684 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2402
timestamp 1682952543
transform 1 0 1724 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2450
timestamp 1682952543
transform 1 0 1692 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1682952543
transform 1 0 1796 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2496
timestamp 1682952543
transform 1 0 1796 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2321
timestamp 1682952543
transform 1 0 1892 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1682952543
transform 1 0 1844 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1682952543
transform 1 0 1868 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2405
timestamp 1682952543
transform 1 0 1892 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1682952543
transform 1 0 1844 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2451
timestamp 1682952543
transform 1 0 1828 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2322
timestamp 1682952543
transform 1 0 1924 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2323
timestamp 1682952543
transform 1 0 1996 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2406
timestamp 1682952543
transform 1 0 1996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1682952543
transform 1 0 1916 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2499
timestamp 1682952543
transform 1 0 1956 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2274
timestamp 1682952543
transform 1 0 2020 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1682952543
transform 1 0 2068 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1682952543
transform 1 0 2100 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2324
timestamp 1682952543
transform 1 0 2028 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2407
timestamp 1682952543
transform 1 0 2028 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2500
timestamp 1682952543
transform 1 0 2052 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1682952543
transform 1 0 2108 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2502
timestamp 1682952543
transform 1 0 2116 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2295
timestamp 1682952543
transform 1 0 2140 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1682952543
transform 1 0 2172 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2408
timestamp 1682952543
transform 1 0 2140 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1682952543
transform 1 0 2156 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2503
timestamp 1682952543
transform 1 0 2172 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2325
timestamp 1682952543
transform 1 0 2204 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1682952543
transform 1 0 2236 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2410
timestamp 1682952543
transform 1 0 2204 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2411
timestamp 1682952543
transform 1 0 2212 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1682952543
transform 1 0 2236 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2345
timestamp 1682952543
transform 1 0 2276 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1682952543
transform 1 0 2324 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2504
timestamp 1682952543
transform 1 0 2220 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2505
timestamp 1682952543
transform 1 0 2284 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1682952543
transform 1 0 2316 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1682952543
transform 1 0 2324 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1682952543
transform 1 0 2332 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2403
timestamp 1682952543
transform 1 0 2212 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2297
timestamp 1682952543
transform 1 0 2372 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1682952543
transform 1 0 2412 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1682952543
transform 1 0 2356 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2328
timestamp 1682952543
transform 1 0 2380 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2413
timestamp 1682952543
transform 1 0 2356 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1682952543
transform 1 0 2372 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1682952543
transform 1 0 2380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1682952543
transform 1 0 2412 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2509
timestamp 1682952543
transform 1 0 2364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1682952543
transform 1 0 2380 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1682952543
transform 1 0 2388 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2512
timestamp 1682952543
transform 1 0 2404 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1682952543
transform 1 0 2420 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2404
timestamp 1682952543
transform 1 0 2380 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2433
timestamp 1682952543
transform 1 0 2388 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1682952543
transform 1 0 2428 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1682952543
transform 1 0 2444 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2417
timestamp 1682952543
transform 1 0 2524 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2368
timestamp 1682952543
transform 1 0 2444 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_2514
timestamp 1682952543
transform 1 0 2476 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1682952543
transform 1 0 2500 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2516
timestamp 1682952543
transform 1 0 2540 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2329
timestamp 1682952543
transform 1 0 2628 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1682952543
transform 1 0 2580 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2418
timestamp 1682952543
transform 1 0 2628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2517
timestamp 1682952543
transform 1 0 2580 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1682952543
transform 1 0 2588 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2519
timestamp 1682952543
transform 1 0 2652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2354
timestamp 1682952543
transform 1 0 2668 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_2520
timestamp 1682952543
transform 1 0 2708 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2330
timestamp 1682952543
transform 1 0 2812 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1682952543
transform 1 0 2732 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1682952543
transform 1 0 2772 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1682952543
transform 1 0 2788 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2419
timestamp 1682952543
transform 1 0 2812 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1682952543
transform 1 0 2732 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1682952543
transform 1 0 2788 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2554
timestamp 1682952543
transform 1 0 2724 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1682952543
transform 1 0 2828 0 1 3145
box -2 -2 2 2
use M3_M2  M3_M2_2352
timestamp 1682952543
transform 1 0 2828 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2420
timestamp 1682952543
transform 1 0 2844 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2523
timestamp 1682952543
transform 1 0 2852 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2405
timestamp 1682952543
transform 1 0 2852 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1682952543
transform 1 0 2868 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1682952543
transform 1 0 2892 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1682952543
transform 1 0 2948 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2421
timestamp 1682952543
transform 1 0 2948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2524
timestamp 1682952543
transform 1 0 2868 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1682952543
transform 1 0 2924 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2460
timestamp 1682952543
transform 1 0 2940 0 1 3085
box -3 -3 3 3
use M2_M1  M2_M1_2356
timestamp 1682952543
transform 1 0 2972 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1682952543
transform 1 0 2964 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2406
timestamp 1682952543
transform 1 0 2964 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1682952543
transform 1 0 2988 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1682952543
transform 1 0 3012 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2423
timestamp 1682952543
transform 1 0 2996 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2526
timestamp 1682952543
transform 1 0 2988 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2461
timestamp 1682952543
transform 1 0 2980 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1682952543
transform 1 0 3004 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2527
timestamp 1682952543
transform 1 0 3012 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1682952543
transform 1 0 3036 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2407
timestamp 1682952543
transform 1 0 3012 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_2424
timestamp 1682952543
transform 1 0 3068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2529
timestamp 1682952543
transform 1 0 3092 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2408
timestamp 1682952543
transform 1 0 3092 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1682952543
transform 1 0 3124 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2425
timestamp 1682952543
transform 1 0 3116 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2278
timestamp 1682952543
transform 1 0 3164 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1682952543
transform 1 0 3228 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2357
timestamp 1682952543
transform 1 0 3236 0 1 3145
box -2 -2 2 2
use M3_M2  M3_M2_2355
timestamp 1682952543
transform 1 0 3140 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2530
timestamp 1682952543
transform 1 0 3132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2531
timestamp 1682952543
transform 1 0 3140 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1682952543
transform 1 0 3148 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2435
timestamp 1682952543
transform 1 0 3188 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2334
timestamp 1682952543
transform 1 0 3252 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2426
timestamp 1682952543
transform 1 0 3252 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2409
timestamp 1682952543
transform 1 0 3252 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1682952543
transform 1 0 3332 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2358
timestamp 1682952543
transform 1 0 3372 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1682952543
transform 1 0 3268 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2356
timestamp 1682952543
transform 1 0 3324 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1682952543
transform 1 0 3380 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2428
timestamp 1682952543
transform 1 0 3388 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2369
timestamp 1682952543
transform 1 0 3268 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_2533
timestamp 1682952543
transform 1 0 3276 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2534
timestamp 1682952543
transform 1 0 3284 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2370
timestamp 1682952543
transform 1 0 3316 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2436
timestamp 1682952543
transform 1 0 3260 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_2558
timestamp 1682952543
transform 1 0 3260 0 1 3095
box -2 -2 2 2
use M3_M2  M3_M2_2410
timestamp 1682952543
transform 1 0 3284 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2437
timestamp 1682952543
transform 1 0 3300 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2438
timestamp 1682952543
transform 1 0 3316 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2439
timestamp 1682952543
transform 1 0 3348 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2452
timestamp 1682952543
transform 1 0 3276 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1682952543
transform 1 0 3324 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1682952543
transform 1 0 3404 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2429
timestamp 1682952543
transform 1 0 3404 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2371
timestamp 1682952543
transform 1 0 3404 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1682952543
transform 1 0 3500 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2430
timestamp 1682952543
transform 1 0 3500 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2279
timestamp 1682952543
transform 1 0 3684 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2336
timestamp 1682952543
transform 1 0 3596 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2431
timestamp 1682952543
transform 1 0 3596 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2358
timestamp 1682952543
transform 1 0 3644 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2535
timestamp 1682952543
transform 1 0 3428 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2536
timestamp 1682952543
transform 1 0 3484 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1682952543
transform 1 0 3548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2538
timestamp 1682952543
transform 1 0 3580 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2411
timestamp 1682952543
transform 1 0 3388 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2412
timestamp 1682952543
transform 1 0 3548 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2462
timestamp 1682952543
transform 1 0 3572 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2372
timestamp 1682952543
transform 1 0 3636 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2302
timestamp 1682952543
transform 1 0 3764 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2359
timestamp 1682952543
transform 1 0 3780 0 1 3145
box -2 -2 2 2
use M3_M2  M3_M2_2359
timestamp 1682952543
transform 1 0 3700 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2432
timestamp 1682952543
transform 1 0 3764 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2539
timestamp 1682952543
transform 1 0 3644 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2540
timestamp 1682952543
transform 1 0 3676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2541
timestamp 1682952543
transform 1 0 3684 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1682952543
transform 1 0 3740 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2373
timestamp 1682952543
transform 1 0 3780 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2413
timestamp 1682952543
transform 1 0 3740 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2414
timestamp 1682952543
transform 1 0 3780 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2454
timestamp 1682952543
transform 1 0 3692 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1682952543
transform 1 0 3804 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2433
timestamp 1682952543
transform 1 0 3796 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2543
timestamp 1682952543
transform 1 0 3796 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2544
timestamp 1682952543
transform 1 0 3820 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2545
timestamp 1682952543
transform 1 0 3836 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2415
timestamp 1682952543
transform 1 0 3796 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_2555
timestamp 1682952543
transform 1 0 3804 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_2416
timestamp 1682952543
transform 1 0 3820 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_2556
timestamp 1682952543
transform 1 0 3828 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1682952543
transform 1 0 3812 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1682952543
transform 1 0 3844 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2360
timestamp 1682952543
transform 1 0 3852 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_2546
timestamp 1682952543
transform 1 0 3844 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2417
timestamp 1682952543
transform 1 0 3844 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2338
timestamp 1682952543
transform 1 0 3876 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_2435
timestamp 1682952543
transform 1 0 3860 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1682952543
transform 1 0 3876 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2303
timestamp 1682952543
transform 1 0 3972 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2437
timestamp 1682952543
transform 1 0 3972 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2361
timestamp 1682952543
transform 1 0 3996 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2304
timestamp 1682952543
transform 1 0 4068 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_2438
timestamp 1682952543
transform 1 0 4068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1682952543
transform 1 0 3908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2548
timestamp 1682952543
transform 1 0 3956 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2549
timestamp 1682952543
transform 1 0 3996 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2550
timestamp 1682952543
transform 1 0 4020 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1682952543
transform 1 0 4052 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1682952543
transform 1 0 4092 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1682952543
transform 1 0 4148 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2418
timestamp 1682952543
transform 1 0 3860 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1682952543
transform 1 0 3908 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2441
timestamp 1682952543
transform 1 0 3948 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2455
timestamp 1682952543
transform 1 0 3892 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2463
timestamp 1682952543
transform 1 0 3884 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2419
timestamp 1682952543
transform 1 0 4036 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2464
timestamp 1682952543
transform 1 0 4028 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1682952543
transform 1 0 4092 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2465
timestamp 1682952543
transform 1 0 4140 0 1 3085
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_20
timestamp 1682952543
transform 1 0 24 0 1 3070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_139
timestamp 1682952543
transform 1 0 72 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_161
timestamp 1682952543
transform -1 0 184 0 -1 3170
box -9 -3 26 105
use AOI22X1  AOI22X1_73
timestamp 1682952543
transform -1 0 224 0 -1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_141
timestamp 1682952543
transform 1 0 224 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_163
timestamp 1682952543
transform 1 0 320 0 -1 3170
box -9 -3 26 105
use AOI22X1  AOI22X1_74
timestamp 1682952543
transform 1 0 336 0 -1 3170
box -8 -3 46 105
use FILL  FILL_655
timestamp 1682952543
transform 1 0 376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_656
timestamp 1682952543
transform 1 0 384 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_159
timestamp 1682952543
transform -1 0 432 0 -1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_142
timestamp 1682952543
transform 1 0 432 0 -1 3170
box -8 -3 104 105
use AOI22X1  AOI22X1_75
timestamp 1682952543
transform 1 0 528 0 -1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_144
timestamp 1682952543
transform 1 0 568 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_165
timestamp 1682952543
transform 1 0 664 0 -1 3170
box -9 -3 26 105
use FILL  FILL_661
timestamp 1682952543
transform 1 0 680 0 -1 3170
box -8 -3 16 105
use FILL  FILL_662
timestamp 1682952543
transform 1 0 688 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2466
timestamp 1682952543
transform 1 0 740 0 1 3075
box -3 -3 3 3
use OAI22X1  OAI22X1_160
timestamp 1682952543
transform 1 0 696 0 -1 3170
box -8 -3 46 105
use FILL  FILL_663
timestamp 1682952543
transform 1 0 736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_664
timestamp 1682952543
transform 1 0 744 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_161
timestamp 1682952543
transform 1 0 752 0 -1 3170
box -8 -3 46 105
use FILL  FILL_676
timestamp 1682952543
transform 1 0 792 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2467
timestamp 1682952543
transform 1 0 860 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2468
timestamp 1682952543
transform 1 0 876 0 1 3075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_145
timestamp 1682952543
transform -1 0 896 0 -1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2469
timestamp 1682952543
transform 1 0 908 0 1 3075
box -3 -3 3 3
use INVX2  INVX2_167
timestamp 1682952543
transform -1 0 912 0 -1 3170
box -9 -3 26 105
use FILL  FILL_677
timestamp 1682952543
transform 1 0 912 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2470
timestamp 1682952543
transform 1 0 932 0 1 3075
box -3 -3 3 3
use NOR2X1  NOR2X1_18
timestamp 1682952543
transform 1 0 920 0 -1 3170
box -8 -3 32 105
use FILL  FILL_679
timestamp 1682952543
transform 1 0 944 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_146
timestamp 1682952543
transform 1 0 952 0 -1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2471
timestamp 1682952543
transform 1 0 1060 0 1 3075
box -3 -3 3 3
use FILL  FILL_688
timestamp 1682952543
transform 1 0 1048 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_169
timestamp 1682952543
transform -1 0 1072 0 -1 3170
box -9 -3 26 105
use FILL  FILL_689
timestamp 1682952543
transform 1 0 1072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_692
timestamp 1682952543
transform 1 0 1080 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_79
timestamp 1682952543
transform 1 0 1088 0 -1 3170
box -8 -3 46 105
use FILL  FILL_693
timestamp 1682952543
transform 1 0 1128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_698
timestamp 1682952543
transform 1 0 1136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_699
timestamp 1682952543
transform 1 0 1144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_700
timestamp 1682952543
transform 1 0 1152 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_163
timestamp 1682952543
transform -1 0 1200 0 -1 3170
box -8 -3 46 105
use FILL  FILL_701
timestamp 1682952543
transform 1 0 1200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_702
timestamp 1682952543
transform 1 0 1208 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_148
timestamp 1682952543
transform 1 0 1216 0 -1 3170
box -8 -3 104 105
use AOI22X1  AOI22X1_81
timestamp 1682952543
transform -1 0 1352 0 -1 3170
box -8 -3 46 105
use FILL  FILL_703
timestamp 1682952543
transform 1 0 1352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_705
timestamp 1682952543
transform 1 0 1360 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_172
timestamp 1682952543
transform 1 0 1368 0 -1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_150
timestamp 1682952543
transform -1 0 1480 0 -1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2472
timestamp 1682952543
transform 1 0 1524 0 1 3075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_151
timestamp 1682952543
transform 1 0 1480 0 -1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2473
timestamp 1682952543
transform 1 0 1604 0 1 3075
box -3 -3 3 3
use OAI22X1  OAI22X1_166
timestamp 1682952543
transform 1 0 1576 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_83
timestamp 1682952543
transform 1 0 1616 0 -1 3170
box -8 -3 46 105
use INVX2  INVX2_174
timestamp 1682952543
transform 1 0 1656 0 -1 3170
box -9 -3 26 105
use FILL  FILL_717
timestamp 1682952543
transform 1 0 1672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_718
timestamp 1682952543
transform 1 0 1680 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_163
timestamp 1682952543
transform -1 0 1784 0 -1 3170
box -8 -3 104 105
use FILL  FILL_719
timestamp 1682952543
transform 1 0 1784 0 -1 3170
box -8 -3 16 105
use FILL  FILL_720
timestamp 1682952543
transform 1 0 1792 0 -1 3170
box -8 -3 16 105
use FILL  FILL_721
timestamp 1682952543
transform 1 0 1800 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_164
timestamp 1682952543
transform -1 0 1904 0 -1 3170
box -8 -3 104 105
use FILL  FILL_722
timestamp 1682952543
transform 1 0 1904 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_165
timestamp 1682952543
transform -1 0 2008 0 -1 3170
box -8 -3 104 105
use FILL  FILL_723
timestamp 1682952543
transform 1 0 2008 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2474
timestamp 1682952543
transform 1 0 2060 0 1 3075
box -3 -3 3 3
use M3_M2  M3_M2_2475
timestamp 1682952543
transform 1 0 2084 0 1 3075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_166
timestamp 1682952543
transform 1 0 2016 0 -1 3170
box -8 -3 104 105
use FILL  FILL_724
timestamp 1682952543
transform 1 0 2112 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_13
timestamp 1682952543
transform 1 0 2120 0 -1 3170
box -5 -3 28 105
use FILL  FILL_725
timestamp 1682952543
transform 1 0 2144 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_14
timestamp 1682952543
transform -1 0 2176 0 -1 3170
box -5 -3 28 105
use BUFX2  BUFX2_15
timestamp 1682952543
transform 1 0 2176 0 -1 3170
box -5 -3 28 105
use FILL  FILL_726
timestamp 1682952543
transform 1 0 2200 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_181
timestamp 1682952543
transform 1 0 2208 0 -1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_167
timestamp 1682952543
transform 1 0 2224 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_182
timestamp 1682952543
transform -1 0 2336 0 -1 3170
box -9 -3 26 105
use FILL  FILL_727
timestamp 1682952543
transform 1 0 2336 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_86
timestamp 1682952543
transform 1 0 2344 0 -1 3170
box -8 -3 46 105
use AOI22X1  AOI22X1_87
timestamp 1682952543
transform 1 0 2384 0 -1 3170
box -8 -3 46 105
use FILL  FILL_728
timestamp 1682952543
transform 1 0 2424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_729
timestamp 1682952543
transform 1 0 2432 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_168
timestamp 1682952543
transform -1 0 2536 0 -1 3170
box -8 -3 104 105
use FILL  FILL_730
timestamp 1682952543
transform 1 0 2536 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_169
timestamp 1682952543
transform -1 0 2640 0 -1 3170
box -8 -3 104 105
use FILL  FILL_731
timestamp 1682952543
transform 1 0 2640 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_22
timestamp 1682952543
transform -1 0 2672 0 -1 3170
box -8 -3 32 105
use FILL  FILL_732
timestamp 1682952543
transform 1 0 2672 0 -1 3170
box -8 -3 16 105
use FILL  FILL_733
timestamp 1682952543
transform 1 0 2680 0 -1 3170
box -8 -3 16 105
use FILL  FILL_734
timestamp 1682952543
transform 1 0 2688 0 -1 3170
box -8 -3 16 105
use FILL  FILL_735
timestamp 1682952543
transform 1 0 2696 0 -1 3170
box -8 -3 16 105
use NAND2X1  NAND2X1_28
timestamp 1682952543
transform 1 0 2704 0 -1 3170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_170
timestamp 1682952543
transform -1 0 2824 0 -1 3170
box -8 -3 104 105
use FILL  FILL_736
timestamp 1682952543
transform 1 0 2824 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_23
timestamp 1682952543
transform 1 0 2832 0 -1 3170
box -8 -3 32 105
use FILL  FILL_737
timestamp 1682952543
transform 1 0 2856 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_171
timestamp 1682952543
transform -1 0 2960 0 -1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2476
timestamp 1682952543
transform 1 0 2972 0 1 3075
box -3 -3 3 3
use FILL  FILL_738
timestamp 1682952543
transform 1 0 2960 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_24
timestamp 1682952543
transform 1 0 2968 0 -1 3170
box -8 -3 32 105
use FILL  FILL_739
timestamp 1682952543
transform 1 0 2992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_740
timestamp 1682952543
transform 1 0 3000 0 -1 3170
box -8 -3 16 105
use XOR2X1  XOR2X1_0
timestamp 1682952543
transform -1 0 3064 0 -1 3170
box -8 -3 64 105
use FILL  FILL_741
timestamp 1682952543
transform 1 0 3064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_742
timestamp 1682952543
transform 1 0 3072 0 -1 3170
box -8 -3 16 105
use AND2X2  AND2X2_6
timestamp 1682952543
transform 1 0 3080 0 -1 3170
box -8 -3 40 105
use FILL  FILL_743
timestamp 1682952543
transform 1 0 3112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_744
timestamp 1682952543
transform 1 0 3120 0 -1 3170
box -8 -3 16 105
use FAX1  FAX1_0
timestamp 1682952543
transform 1 0 3128 0 -1 3170
box -5 -3 126 105
use FILL  FILL_745
timestamp 1682952543
transform 1 0 3248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_747
timestamp 1682952543
transform 1 0 3256 0 -1 3170
box -8 -3 16 105
use FAX1  FAX1_1
timestamp 1682952543
transform 1 0 3264 0 -1 3170
box -5 -3 126 105
use FILL  FILL_773
timestamp 1682952543
transform 1 0 3384 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_175
timestamp 1682952543
transform 1 0 3392 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_176
timestamp 1682952543
transform 1 0 3488 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_177
timestamp 1682952543
transform 1 0 3584 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_178
timestamp 1682952543
transform -1 0 3776 0 -1 3170
box -8 -3 104 105
use M3_M2  M3_M2_2477
timestamp 1682952543
transform 1 0 3804 0 1 3075
box -3 -3 3 3
use NOR2X1  NOR2X1_25
timestamp 1682952543
transform 1 0 3776 0 -1 3170
box -8 -3 32 105
use NAND3X1  NAND3X1_0
timestamp 1682952543
transform -1 0 3832 0 -1 3170
box -8 -3 40 105
use INVX2  INVX2_188
timestamp 1682952543
transform -1 0 3848 0 -1 3170
box -9 -3 26 105
use INVX2  INVX2_189
timestamp 1682952543
transform -1 0 3864 0 -1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_179
timestamp 1682952543
transform 1 0 3864 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_180
timestamp 1682952543
transform 1 0 3960 0 -1 3170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_181
timestamp 1682952543
transform 1 0 4056 0 -1 3170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_21
timestamp 1682952543
transform 1 0 4201 0 1 3070
box -10 -3 10 3
use M2_M1  M2_M1_2570
timestamp 1682952543
transform 1 0 132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2571
timestamp 1682952543
transform 1 0 164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1682952543
transform 1 0 172 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2710
timestamp 1682952543
transform 1 0 84 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1682952543
transform 1 0 188 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1682952543
transform 1 0 188 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2712
timestamp 1682952543
transform 1 0 196 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2713
timestamp 1682952543
transform 1 0 220 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2541
timestamp 1682952543
transform 1 0 236 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2574
timestamp 1682952543
transform 1 0 228 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1682952543
transform 1 0 236 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2513
timestamp 1682952543
transform 1 0 252 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1682952543
transform 1 0 268 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2575
timestamp 1682952543
transform 1 0 244 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1682952543
transform 1 0 268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2715
timestamp 1682952543
transform 1 0 252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1682952543
transform 1 0 260 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2667
timestamp 1682952543
transform 1 0 276 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2708
timestamp 1682952543
transform 1 0 260 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_2577
timestamp 1682952543
transform 1 0 292 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2633
timestamp 1682952543
transform 1 0 292 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2717
timestamp 1682952543
transform 1 0 300 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2478
timestamp 1682952543
transform 1 0 412 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2543
timestamp 1682952543
transform 1 0 460 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2544
timestamp 1682952543
transform 1 0 500 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2578
timestamp 1682952543
transform 1 0 340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1682952543
transform 1 0 396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2718
timestamp 1682952543
transform 1 0 316 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2634
timestamp 1682952543
transform 1 0 356 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1682952543
transform 1 0 316 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1682952543
transform 1 0 380 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2709
timestamp 1682952543
transform 1 0 308 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1682952543
transform 1 0 348 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2589
timestamp 1682952543
transform 1 0 412 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2590
timestamp 1682952543
transform 1 0 444 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1682952543
transform 1 0 548 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2580
timestamp 1682952543
transform 1 0 460 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1682952543
transform 1 0 492 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1682952543
transform 1 0 500 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1682952543
transform 1 0 516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1682952543
transform 1 0 412 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2591
timestamp 1682952543
transform 1 0 524 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2584
timestamp 1682952543
transform 1 0 532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1682952543
transform 1 0 548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1682952543
transform 1 0 556 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1682952543
transform 1 0 516 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2721
timestamp 1682952543
transform 1 0 524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1682952543
transform 1 0 540 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2670
timestamp 1682952543
transform 1 0 492 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1682952543
transform 1 0 540 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1682952543
transform 1 0 572 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2514
timestamp 1682952543
transform 1 0 572 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2546
timestamp 1682952543
transform 1 0 564 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1682952543
transform 1 0 612 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1682952543
transform 1 0 620 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2516
timestamp 1682952543
transform 1 0 636 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1682952543
transform 1 0 604 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2592
timestamp 1682952543
transform 1 0 564 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2587
timestamp 1682952543
transform 1 0 572 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2593
timestamp 1682952543
transform 1 0 580 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1682952543
transform 1 0 644 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2588
timestamp 1682952543
transform 1 0 588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2589
timestamp 1682952543
transform 1 0 604 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2594
timestamp 1682952543
transform 1 0 620 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1682952543
transform 1 0 748 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2590
timestamp 1682952543
transform 1 0 628 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1682952543
transform 1 0 644 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2595
timestamp 1682952543
transform 1 0 660 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2550
timestamp 1682952543
transform 1 0 780 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2592
timestamp 1682952543
transform 1 0 708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1682952543
transform 1 0 748 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1682952543
transform 1 0 756 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1682952543
transform 1 0 772 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1682952543
transform 1 0 788 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2723
timestamp 1682952543
transform 1 0 572 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1682952543
transform 1 0 580 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1682952543
transform 1 0 596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2726
timestamp 1682952543
transform 1 0 612 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2727
timestamp 1682952543
transform 1 0 620 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2728
timestamp 1682952543
transform 1 0 644 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1682952543
transform 1 0 660 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2635
timestamp 1682952543
transform 1 0 708 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1682952543
transform 1 0 804 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1682952543
transform 1 0 836 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1682952543
transform 1 0 812 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1682952543
transform 1 0 868 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2552
timestamp 1682952543
transform 1 0 860 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2597
timestamp 1682952543
transform 1 0 804 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1682952543
transform 1 0 820 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2599
timestamp 1682952543
transform 1 0 836 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1682952543
transform 1 0 748 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2731
timestamp 1682952543
transform 1 0 764 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1682952543
transform 1 0 780 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2672
timestamp 1682952543
transform 1 0 644 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2636
timestamp 1682952543
transform 1 0 788 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2733
timestamp 1682952543
transform 1 0 804 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1682952543
transform 1 0 812 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2735
timestamp 1682952543
transform 1 0 828 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2673
timestamp 1682952543
transform 1 0 748 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1682952543
transform 1 0 764 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2711
timestamp 1682952543
transform 1 0 660 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1682952543
transform 1 0 692 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1682952543
transform 1 0 724 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2637
timestamp 1682952543
transform 1 0 844 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1682952543
transform 1 0 900 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1682952543
transform 1 0 900 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2479
timestamp 1682952543
transform 1 0 1004 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_2600
timestamp 1682952543
transform 1 0 860 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1682952543
transform 1 0 868 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1682952543
transform 1 0 884 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1682952543
transform 1 0 900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1682952543
transform 1 0 908 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1682952543
transform 1 0 956 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2736
timestamp 1682952543
transform 1 0 852 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1682952543
transform 1 0 860 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2738
timestamp 1682952543
transform 1 0 892 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2675
timestamp 1682952543
transform 1 0 836 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2825
timestamp 1682952543
transform 1 0 844 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2676
timestamp 1682952543
transform 1 0 860 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1682952543
transform 1 0 828 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2596
timestamp 1682952543
transform 1 0 988 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2739
timestamp 1682952543
transform 1 0 988 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2677
timestamp 1682952543
transform 1 0 908 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1682952543
transform 1 0 972 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1682952543
transform 1 0 988 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2826
timestamp 1682952543
transform 1 0 1004 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2715
timestamp 1682952543
transform 1 0 892 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1682952543
transform 1 0 972 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1682952543
transform 1 0 988 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2490
timestamp 1682952543
transform 1 0 1020 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_2606
timestamp 1682952543
transform 1 0 1020 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2597
timestamp 1682952543
transform 1 0 1028 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2607
timestamp 1682952543
transform 1 0 1036 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2740
timestamp 1682952543
transform 1 0 1020 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1682952543
transform 1 0 1028 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2742
timestamp 1682952543
transform 1 0 1068 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2500
timestamp 1682952543
transform 1 0 1084 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1682952543
transform 1 0 1116 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2608
timestamp 1682952543
transform 1 0 1084 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2598
timestamp 1682952543
transform 1 0 1092 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2609
timestamp 1682952543
transform 1 0 1100 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2599
timestamp 1682952543
transform 1 0 1116 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2610
timestamp 1682952543
transform 1 0 1124 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1682952543
transform 1 0 1092 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2638
timestamp 1682952543
transform 1 0 1100 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2744
timestamp 1682952543
transform 1 0 1108 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2718
timestamp 1682952543
transform 1 0 1084 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_2827
timestamp 1682952543
transform 1 0 1124 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2501
timestamp 1682952543
transform 1 0 1132 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2639
timestamp 1682952543
transform 1 0 1140 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2828
timestamp 1682952543
transform 1 0 1148 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2502
timestamp 1682952543
transform 1 0 1188 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1682952543
transform 1 0 1164 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1682952543
transform 1 0 1172 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2611
timestamp 1682952543
transform 1 0 1164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1682952543
transform 1 0 1180 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1682952543
transform 1 0 1172 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2503
timestamp 1682952543
transform 1 0 1244 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1682952543
transform 1 0 1236 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2746
timestamp 1682952543
transform 1 0 1228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1682952543
transform 1 0 1236 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2680
timestamp 1682952543
transform 1 0 1228 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1682952543
transform 1 0 1260 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2613
timestamp 1682952543
transform 1 0 1252 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2748
timestamp 1682952543
transform 1 0 1252 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2719
timestamp 1682952543
transform 1 0 1252 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2504
timestamp 1682952543
transform 1 0 1292 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1682952543
transform 1 0 1308 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2555
timestamp 1682952543
transform 1 0 1292 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1682952543
transform 1 0 1316 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2614
timestamp 1682952543
transform 1 0 1276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1682952543
transform 1 0 1292 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2640
timestamp 1682952543
transform 1 0 1276 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2600
timestamp 1682952543
transform 1 0 1308 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2616
timestamp 1682952543
transform 1 0 1316 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2749
timestamp 1682952543
transform 1 0 1300 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2750
timestamp 1682952543
transform 1 0 1308 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2681
timestamp 1682952543
transform 1 0 1300 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2617
timestamp 1682952543
transform 1 0 1324 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2601
timestamp 1682952543
transform 1 0 1332 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2557
timestamp 1682952543
transform 1 0 1372 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2618
timestamp 1682952543
transform 1 0 1340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1682952543
transform 1 0 1356 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2641
timestamp 1682952543
transform 1 0 1324 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2602
timestamp 1682952543
transform 1 0 1364 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2620
timestamp 1682952543
transform 1 0 1372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1682952543
transform 1 0 1364 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1682952543
transform 1 0 1372 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2558
timestamp 1682952543
transform 1 0 1388 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1682952543
transform 1 0 1420 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2481
timestamp 1682952543
transform 1 0 1492 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2505
timestamp 1682952543
transform 1 0 1452 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2506
timestamp 1682952543
transform 1 0 1468 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1682952543
transform 1 0 1436 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2621
timestamp 1682952543
transform 1 0 1388 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2622
timestamp 1682952543
transform 1 0 1404 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2603
timestamp 1682952543
transform 1 0 1412 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2623
timestamp 1682952543
transform 1 0 1436 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1682952543
transform 1 0 1516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2753
timestamp 1682952543
transform 1 0 1484 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2754
timestamp 1682952543
transform 1 0 1500 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2642
timestamp 1682952543
transform 1 0 1508 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2682
timestamp 1682952543
transform 1 0 1508 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1682952543
transform 1 0 1460 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1682952543
transform 1 0 1500 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1682952543
transform 1 0 1532 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2560
timestamp 1682952543
transform 1 0 1564 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2625
timestamp 1682952543
transform 1 0 1532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1682952543
transform 1 0 1548 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2627
timestamp 1682952543
transform 1 0 1564 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2755
timestamp 1682952543
transform 1 0 1540 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2643
timestamp 1682952543
transform 1 0 1548 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2756
timestamp 1682952543
transform 1 0 1556 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2722
timestamp 1682952543
transform 1 0 1540 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_2757
timestamp 1682952543
transform 1 0 1572 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1682952543
transform 1 0 1572 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2482
timestamp 1682952543
transform 1 0 1588 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1682952543
transform 1 0 1580 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2491
timestamp 1682952543
transform 1 0 1596 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2492
timestamp 1682952543
transform 1 0 1612 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1682952543
transform 1 0 1596 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1682952543
transform 1 0 1628 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1682952543
transform 1 0 1604 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1682952543
transform 1 0 1620 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2628
timestamp 1682952543
transform 1 0 1588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2629
timestamp 1682952543
transform 1 0 1604 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2605
timestamp 1682952543
transform 1 0 1612 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2630
timestamp 1682952543
transform 1 0 1620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2758
timestamp 1682952543
transform 1 0 1588 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1682952543
transform 1 0 1596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2760
timestamp 1682952543
transform 1 0 1612 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1682952543
transform 1 0 1620 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2723
timestamp 1682952543
transform 1 0 1588 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2526
timestamp 1682952543
transform 1 0 1652 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1682952543
transform 1 0 1724 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1682952543
transform 1 0 1764 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2562
timestamp 1682952543
transform 1 0 1636 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2563
timestamp 1682952543
transform 1 0 1676 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2564
timestamp 1682952543
transform 1 0 1740 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2631
timestamp 1682952543
transform 1 0 1636 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2632
timestamp 1682952543
transform 1 0 1644 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2606
timestamp 1682952543
transform 1 0 1652 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1682952543
transform 1 0 1772 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2633
timestamp 1682952543
transform 1 0 1676 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1682952543
transform 1 0 1740 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2635
timestamp 1682952543
transform 1 0 1756 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2607
timestamp 1682952543
transform 1 0 1764 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2636
timestamp 1682952543
transform 1 0 1772 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1682952543
transform 1 0 1780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2762
timestamp 1682952543
transform 1 0 1724 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2763
timestamp 1682952543
transform 1 0 1740 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2764
timestamp 1682952543
transform 1 0 1764 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1682952543
transform 1 0 1772 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2565
timestamp 1682952543
transform 1 0 1796 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2566
timestamp 1682952543
transform 1 0 1820 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2638
timestamp 1682952543
transform 1 0 1796 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1682952543
transform 1 0 1812 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2608
timestamp 1682952543
transform 1 0 1820 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2640
timestamp 1682952543
transform 1 0 1828 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2609
timestamp 1682952543
transform 1 0 1836 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2641
timestamp 1682952543
transform 1 0 1844 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1682952543
transform 1 0 1804 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2767
timestamp 1682952543
transform 1 0 1820 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1682952543
transform 1 0 1828 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2724
timestamp 1682952543
transform 1 0 1796 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1682952543
transform 1 0 1860 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1682952543
transform 1 0 1860 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2642
timestamp 1682952543
transform 1 0 1860 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1682952543
transform 1 0 1860 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2683
timestamp 1682952543
transform 1 0 1860 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1682952543
transform 1 0 1908 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2529
timestamp 1682952543
transform 1 0 1908 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1682952543
transform 1 0 1940 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2643
timestamp 1682952543
transform 1 0 1876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1682952543
transform 1 0 1892 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2725
timestamp 1682952543
transform 1 0 1868 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2610
timestamp 1682952543
transform 1 0 1900 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2568
timestamp 1682952543
transform 1 0 1924 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1682952543
transform 1 0 1980 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2645
timestamp 1682952543
transform 1 0 1908 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2646
timestamp 1682952543
transform 1 0 1924 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1682952543
transform 1 0 1932 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2770
timestamp 1682952543
transform 1 0 1900 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1682952543
transform 1 0 1908 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2611
timestamp 1682952543
transform 1 0 1964 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2648
timestamp 1682952543
transform 1 0 1980 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1682952543
transform 1 0 2012 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2684
timestamp 1682952543
transform 1 0 1932 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1682952543
transform 1 0 2108 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1682952543
transform 1 0 2092 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1682952543
transform 1 0 2060 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1682952543
transform 1 0 2268 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2531
timestamp 1682952543
transform 1 0 2244 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2570
timestamp 1682952543
transform 1 0 2260 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2649
timestamp 1682952543
transform 1 0 2076 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1682952543
transform 1 0 2116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1682952543
transform 1 0 2180 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1682952543
transform 1 0 2212 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1682952543
transform 1 0 2228 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2654
timestamp 1682952543
transform 1 0 2244 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1682952543
transform 1 0 2260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2773
timestamp 1682952543
transform 1 0 2036 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2774
timestamp 1682952543
transform 1 0 2132 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2644
timestamp 1682952543
transform 1 0 2212 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2775
timestamp 1682952543
transform 1 0 2220 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2645
timestamp 1682952543
transform 1 0 2228 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2776
timestamp 1682952543
transform 1 0 2236 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2777
timestamp 1682952543
transform 1 0 2252 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2685
timestamp 1682952543
transform 1 0 2132 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2686
timestamp 1682952543
transform 1 0 2164 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2687
timestamp 1682952543
transform 1 0 2180 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1682952543
transform 1 0 2084 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1682952543
transform 1 0 2124 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2728
timestamp 1682952543
transform 1 0 2212 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2688
timestamp 1682952543
transform 1 0 2252 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2656
timestamp 1682952543
transform 1 0 2276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1682952543
transform 1 0 2276 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2532
timestamp 1682952543
transform 1 0 2292 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2571
timestamp 1682952543
transform 1 0 2308 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2657
timestamp 1682952543
transform 1 0 2292 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1682952543
transform 1 0 2308 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2646
timestamp 1682952543
transform 1 0 2292 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2779
timestamp 1682952543
transform 1 0 2300 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2689
timestamp 1682952543
transform 1 0 2276 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2659
timestamp 1682952543
transform 1 0 2332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1682952543
transform 1 0 2340 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2612
timestamp 1682952543
transform 1 0 2348 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2661
timestamp 1682952543
transform 1 0 2356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1682952543
transform 1 0 2324 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2647
timestamp 1682952543
transform 1 0 2332 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2781
timestamp 1682952543
transform 1 0 2340 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2648
timestamp 1682952543
transform 1 0 2348 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2782
timestamp 1682952543
transform 1 0 2356 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2729
timestamp 1682952543
transform 1 0 2340 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1682952543
transform 1 0 2356 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1682952543
transform 1 0 2388 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2562
timestamp 1682952543
transform 1 0 2404 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_2573
timestamp 1682952543
transform 1 0 2412 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2662
timestamp 1682952543
transform 1 0 2388 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1682952543
transform 1 0 2372 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2690
timestamp 1682952543
transform 1 0 2372 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1682952543
transform 1 0 2460 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_2663
timestamp 1682952543
transform 1 0 2412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1682952543
transform 1 0 2404 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2613
timestamp 1682952543
transform 1 0 2420 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2664
timestamp 1682952543
transform 1 0 2428 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1682952543
transform 1 0 2484 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2785
timestamp 1682952543
transform 1 0 2420 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2649
timestamp 1682952543
transform 1 0 2484 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2786
timestamp 1682952543
transform 1 0 2508 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2731
timestamp 1682952543
transform 1 0 2428 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1682952543
transform 1 0 2580 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2666
timestamp 1682952543
transform 1 0 2532 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2614
timestamp 1682952543
transform 1 0 2540 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2667
timestamp 1682952543
transform 1 0 2580 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2615
timestamp 1682952543
transform 1 0 2612 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2787
timestamp 1682952543
transform 1 0 2612 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2574
timestamp 1682952543
transform 1 0 2660 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2616
timestamp 1682952543
transform 1 0 2636 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2668
timestamp 1682952543
transform 1 0 2660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2669
timestamp 1682952543
transform 1 0 2724 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1682952543
transform 1 0 2636 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2650
timestamp 1682952543
transform 1 0 2716 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2789
timestamp 1682952543
transform 1 0 2724 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2691
timestamp 1682952543
transform 1 0 2636 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2830
timestamp 1682952543
transform 1 0 2724 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2732
timestamp 1682952543
transform 1 0 2628 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2733
timestamp 1682952543
transform 1 0 2668 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2575
timestamp 1682952543
transform 1 0 2740 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2563
timestamp 1682952543
transform 1 0 2748 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_2617
timestamp 1682952543
transform 1 0 2748 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1682952543
transform 1 0 2764 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1682952543
transform 1 0 2796 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2576
timestamp 1682952543
transform 1 0 2788 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2790
timestamp 1682952543
transform 1 0 2780 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2692
timestamp 1682952543
transform 1 0 2780 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2791
timestamp 1682952543
transform 1 0 2796 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1682952543
transform 1 0 2788 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1682952543
transform 1 0 2812 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_2618
timestamp 1682952543
transform 1 0 2812 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1682952543
transform 1 0 2836 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1682952543
transform 1 0 2828 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2792
timestamp 1682952543
transform 1 0 2836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1682952543
transform 1 0 2844 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2693
timestamp 1682952543
transform 1 0 2844 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2620
timestamp 1682952543
transform 1 0 2852 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2670
timestamp 1682952543
transform 1 0 2860 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2652
timestamp 1682952543
transform 1 0 2852 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2794
timestamp 1682952543
transform 1 0 2860 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1682952543
transform 1 0 2876 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_2577
timestamp 1682952543
transform 1 0 2884 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2671
timestamp 1682952543
transform 1 0 2876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2672
timestamp 1682952543
transform 1 0 2884 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2621
timestamp 1682952543
transform 1 0 2900 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2795
timestamp 1682952543
transform 1 0 2892 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1682952543
transform 1 0 2900 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2535
timestamp 1682952543
transform 1 0 2924 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2673
timestamp 1682952543
transform 1 0 2916 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1682952543
transform 1 0 2924 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2559
timestamp 1682952543
transform 1 0 2980 0 1 3035
box -2 -2 2 2
use M3_M2  M3_M2_2578
timestamp 1682952543
transform 1 0 2948 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2566
timestamp 1682952543
transform 1 0 2964 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_2579
timestamp 1682952543
transform 1 0 2972 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2567
timestamp 1682952543
transform 1 0 2988 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1682952543
transform 1 0 2948 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2675
timestamp 1682952543
transform 1 0 2956 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2676
timestamp 1682952543
transform 1 0 2972 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1682952543
transform 1 0 2940 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2622
timestamp 1682952543
transform 1 0 2980 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1682952543
transform 1 0 2956 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2694
timestamp 1682952543
transform 1 0 2948 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2799
timestamp 1682952543
transform 1 0 2996 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2695
timestamp 1682952543
transform 1 0 2996 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2654
timestamp 1682952543
transform 1 0 3004 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2677
timestamp 1682952543
transform 1 0 3020 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2678
timestamp 1682952543
transform 1 0 3036 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1682952543
transform 1 0 3052 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2511
timestamp 1682952543
transform 1 0 3092 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1682952543
transform 1 0 3068 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2581
timestamp 1682952543
transform 1 0 3100 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2679
timestamp 1682952543
transform 1 0 3076 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1682952543
transform 1 0 3092 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2681
timestamp 1682952543
transform 1 0 3100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1682952543
transform 1 0 3124 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2512
timestamp 1682952543
transform 1 0 3172 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_2682
timestamp 1682952543
transform 1 0 3148 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2683
timestamp 1682952543
transform 1 0 3164 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1682952543
transform 1 0 3172 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1682952543
transform 1 0 3140 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2655
timestamp 1682952543
transform 1 0 3164 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2803
timestamp 1682952543
transform 1 0 3172 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2734
timestamp 1682952543
transform 1 0 3140 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_2560
timestamp 1682952543
transform 1 0 3236 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1682952543
transform 1 0 3220 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1682952543
transform 1 0 3196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2686
timestamp 1682952543
transform 1 0 3212 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2623
timestamp 1682952543
transform 1 0 3220 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2687
timestamp 1682952543
transform 1 0 3228 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1682952543
transform 1 0 3188 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2656
timestamp 1682952543
transform 1 0 3196 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2805
timestamp 1682952543
transform 1 0 3204 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2657
timestamp 1682952543
transform 1 0 3220 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1682952543
transform 1 0 3180 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2496
timestamp 1682952543
transform 1 0 3260 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1682952543
transform 1 0 3260 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2569
timestamp 1682952543
transform 1 0 3260 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_2624
timestamp 1682952543
transform 1 0 3252 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2806
timestamp 1682952543
transform 1 0 3252 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2735
timestamp 1682952543
transform 1 0 3252 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2497
timestamp 1682952543
transform 1 0 3276 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1682952543
transform 1 0 3308 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2688
timestamp 1682952543
transform 1 0 3268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2689
timestamp 1682952543
transform 1 0 3284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2690
timestamp 1682952543
transform 1 0 3300 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1682952543
transform 1 0 3308 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1682952543
transform 1 0 3292 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2808
timestamp 1682952543
transform 1 0 3300 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2697
timestamp 1682952543
transform 1 0 3292 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2809
timestamp 1682952543
transform 1 0 3316 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2582
timestamp 1682952543
transform 1 0 3372 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2692
timestamp 1682952543
transform 1 0 3340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2693
timestamp 1682952543
transform 1 0 3356 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2625
timestamp 1682952543
transform 1 0 3364 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2658
timestamp 1682952543
transform 1 0 3356 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2694
timestamp 1682952543
transform 1 0 3380 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2810
timestamp 1682952543
transform 1 0 3364 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1682952543
transform 1 0 3372 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2698
timestamp 1682952543
transform 1 0 3364 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1682952543
transform 1 0 3348 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_2695
timestamp 1682952543
transform 1 0 3404 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2538
timestamp 1682952543
transform 1 0 3436 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_2696
timestamp 1682952543
transform 1 0 3428 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2697
timestamp 1682952543
transform 1 0 3436 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1682952543
transform 1 0 3436 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2659
timestamp 1682952543
transform 1 0 3452 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1682952543
transform 1 0 3468 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2698
timestamp 1682952543
transform 1 0 3484 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2626
timestamp 1682952543
transform 1 0 3492 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2812
timestamp 1682952543
transform 1 0 3468 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1682952543
transform 1 0 3492 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2584
timestamp 1682952543
transform 1 0 3508 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2699
timestamp 1682952543
transform 1 0 3508 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2487
timestamp 1682952543
transform 1 0 3660 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1682952543
transform 1 0 3724 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1682952543
transform 1 0 3772 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_2585
timestamp 1682952543
transform 1 0 3652 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1682952543
transform 1 0 3524 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2700
timestamp 1682952543
transform 1 0 3540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2701
timestamp 1682952543
transform 1 0 3548 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2628
timestamp 1682952543
transform 1 0 3580 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2814
timestamp 1682952543
transform 1 0 3508 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2660
timestamp 1682952543
transform 1 0 3516 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2815
timestamp 1682952543
transform 1 0 3524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2816
timestamp 1682952543
transform 1 0 3532 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2661
timestamp 1682952543
transform 1 0 3636 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2702
timestamp 1682952543
transform 1 0 3660 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2703
timestamp 1682952543
transform 1 0 3676 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2629
timestamp 1682952543
transform 1 0 3772 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1682952543
transform 1 0 3860 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2561
timestamp 1682952543
transform 1 0 4028 0 1 3035
box -2 -2 2 2
use M3_M2  M3_M2_2586
timestamp 1682952543
transform 1 0 3924 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2587
timestamp 1682952543
transform 1 0 4028 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_2588
timestamp 1682952543
transform 1 0 4052 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_2704
timestamp 1682952543
transform 1 0 3876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1682952543
transform 1 0 3884 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2706
timestamp 1682952543
transform 1 0 3900 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1682952543
transform 1 0 3924 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1682952543
transform 1 0 3652 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1682952543
transform 1 0 3660 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2699
timestamp 1682952543
transform 1 0 3524 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2700
timestamp 1682952543
transform 1 0 3572 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1682952543
transform 1 0 3588 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2833
timestamp 1682952543
transform 1 0 3636 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2737
timestamp 1682952543
transform 1 0 3540 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2738
timestamp 1682952543
transform 1 0 3596 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1682952543
transform 1 0 3676 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1682952543
transform 1 0 3772 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2819
timestamp 1682952543
transform 1 0 3780 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2664
timestamp 1682952543
transform 1 0 3788 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1682952543
transform 1 0 3876 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2820
timestamp 1682952543
transform 1 0 3892 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2702
timestamp 1682952543
transform 1 0 3660 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2703
timestamp 1682952543
transform 1 0 3676 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1682952543
transform 1 0 3716 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2834
timestamp 1682952543
transform 1 0 3764 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1682952543
transform 1 0 3788 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2705
timestamp 1682952543
transform 1 0 3804 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2821
timestamp 1682952543
transform 1 0 3908 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2631
timestamp 1682952543
transform 1 0 4036 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2708
timestamp 1682952543
transform 1 0 4044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_2709
timestamp 1682952543
transform 1 0 4052 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_2632
timestamp 1682952543
transform 1 0 4068 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_2822
timestamp 1682952543
transform 1 0 4028 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2823
timestamp 1682952543
transform 1 0 4036 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_2706
timestamp 1682952543
transform 1 0 3908 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_2707
timestamp 1682952543
transform 1 0 3940 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_2836
timestamp 1682952543
transform 1 0 4012 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2739
timestamp 1682952543
transform 1 0 3980 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1682952543
transform 1 0 4020 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1682952543
transform 1 0 4140 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_2824
timestamp 1682952543
transform 1 0 4148 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_2837
timestamp 1682952543
transform 1 0 4140 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_2741
timestamp 1682952543
transform 1 0 4068 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1682952543
transform 1 0 4108 0 1 2985
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_22
timestamp 1682952543
transform 1 0 48 0 1 2970
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_182
timestamp 1682952543
transform 1 0 72 0 1 2970
box -8 -3 104 105
use FILL  FILL_774
timestamp 1682952543
transform 1 0 168 0 1 2970
box -8 -3 16 105
use FILL  FILL_775
timestamp 1682952543
transform 1 0 176 0 1 2970
box -8 -3 16 105
use FILL  FILL_776
timestamp 1682952543
transform 1 0 184 0 1 2970
box -8 -3 16 105
use FILL  FILL_777
timestamp 1682952543
transform 1 0 192 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_191
timestamp 1682952543
transform 1 0 200 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_192
timestamp 1682952543
transform 1 0 216 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_193
timestamp 1682952543
transform 1 0 232 0 1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_89
timestamp 1682952543
transform 1 0 248 0 1 2970
box -8 -3 46 105
use FILL  FILL_787
timestamp 1682952543
transform 1 0 288 0 1 2970
box -8 -3 16 105
use FILL  FILL_788
timestamp 1682952543
transform 1 0 296 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_183
timestamp 1682952543
transform 1 0 304 0 1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_184
timestamp 1682952543
transform 1 0 400 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_194
timestamp 1682952543
transform -1 0 512 0 1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_90
timestamp 1682952543
transform 1 0 512 0 1 2970
box -8 -3 46 105
use INVX2  INVX2_195
timestamp 1682952543
transform -1 0 568 0 1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_91
timestamp 1682952543
transform 1 0 568 0 1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_92
timestamp 1682952543
transform 1 0 608 0 1 2970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_185
timestamp 1682952543
transform 1 0 648 0 1 2970
box -8 -3 104 105
use M3_M2  M3_M2_2743
timestamp 1682952543
transform 1 0 756 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1682952543
transform 1 0 796 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_172
timestamp 1682952543
transform 1 0 744 0 1 2970
box -8 -3 46 105
use INVX2  INVX2_196
timestamp 1682952543
transform -1 0 800 0 1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_93
timestamp 1682952543
transform -1 0 840 0 1 2970
box -8 -3 46 105
use M3_M2  M3_M2_2745
timestamp 1682952543
transform 1 0 868 0 1 2975
box -3 -3 3 3
use NOR2X1  NOR2X1_26
timestamp 1682952543
transform 1 0 840 0 1 2970
box -8 -3 32 105
use AOI22X1  AOI22X1_94
timestamp 1682952543
transform -1 0 904 0 1 2970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_186
timestamp 1682952543
transform -1 0 1000 0 1 2970
box -8 -3 104 105
use M3_M2  M3_M2_2746
timestamp 1682952543
transform 1 0 1012 0 1 2975
box -3 -3 3 3
use NOR2X1  NOR2X1_27
timestamp 1682952543
transform 1 0 1000 0 1 2970
box -8 -3 32 105
use INVX2  INVX2_197
timestamp 1682952543
transform 1 0 1024 0 1 2970
box -9 -3 26 105
use FILL  FILL_789
timestamp 1682952543
transform 1 0 1040 0 1 2970
box -8 -3 16 105
use FILL  FILL_790
timestamp 1682952543
transform 1 0 1048 0 1 2970
box -8 -3 16 105
use FILL  FILL_791
timestamp 1682952543
transform 1 0 1056 0 1 2970
box -8 -3 16 105
use FILL  FILL_792
timestamp 1682952543
transform 1 0 1064 0 1 2970
box -8 -3 16 105
use FILL  FILL_793
timestamp 1682952543
transform 1 0 1072 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_95
timestamp 1682952543
transform 1 0 1080 0 1 2970
box -8 -3 46 105
use FILL  FILL_794
timestamp 1682952543
transform 1 0 1120 0 1 2970
box -8 -3 16 105
use FILL  FILL_795
timestamp 1682952543
transform 1 0 1128 0 1 2970
box -8 -3 16 105
use FILL  FILL_796
timestamp 1682952543
transform 1 0 1136 0 1 2970
box -8 -3 16 105
use FILL  FILL_797
timestamp 1682952543
transform 1 0 1144 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_173
timestamp 1682952543
transform -1 0 1192 0 1 2970
box -8 -3 46 105
use FILL  FILL_798
timestamp 1682952543
transform 1 0 1192 0 1 2970
box -8 -3 16 105
use FILL  FILL_799
timestamp 1682952543
transform 1 0 1200 0 1 2970
box -8 -3 16 105
use FILL  FILL_800
timestamp 1682952543
transform 1 0 1208 0 1 2970
box -8 -3 16 105
use FILL  FILL_801
timestamp 1682952543
transform 1 0 1216 0 1 2970
box -8 -3 16 105
use FILL  FILL_802
timestamp 1682952543
transform 1 0 1224 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_198
timestamp 1682952543
transform 1 0 1232 0 1 2970
box -9 -3 26 105
use FILL  FILL_803
timestamp 1682952543
transform 1 0 1248 0 1 2970
box -8 -3 16 105
use FILL  FILL_804
timestamp 1682952543
transform 1 0 1256 0 1 2970
box -8 -3 16 105
use FILL  FILL_805
timestamp 1682952543
transform 1 0 1264 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_96
timestamp 1682952543
transform 1 0 1272 0 1 2970
box -8 -3 46 105
use FILL  FILL_806
timestamp 1682952543
transform 1 0 1312 0 1 2970
box -8 -3 16 105
use FILL  FILL_807
timestamp 1682952543
transform 1 0 1320 0 1 2970
box -8 -3 16 105
use FILL  FILL_808
timestamp 1682952543
transform 1 0 1328 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_97
timestamp 1682952543
transform 1 0 1336 0 1 2970
box -8 -3 46 105
use FILL  FILL_809
timestamp 1682952543
transform 1 0 1376 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_199
timestamp 1682952543
transform 1 0 1384 0 1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_187
timestamp 1682952543
transform -1 0 1496 0 1 2970
box -8 -3 104 105
use M3_M2  M3_M2_2747
timestamp 1682952543
transform 1 0 1516 0 1 2975
box -3 -3 3 3
use INVX2  INVX2_200
timestamp 1682952543
transform 1 0 1496 0 1 2970
box -9 -3 26 105
use FILL  FILL_810
timestamp 1682952543
transform 1 0 1512 0 1 2970
box -8 -3 16 105
use FILL  FILL_811
timestamp 1682952543
transform 1 0 1520 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_98
timestamp 1682952543
transform 1 0 1528 0 1 2970
box -8 -3 46 105
use FILL  FILL_812
timestamp 1682952543
transform 1 0 1568 0 1 2970
box -8 -3 16 105
use FILL  FILL_813
timestamp 1682952543
transform 1 0 1576 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_99
timestamp 1682952543
transform 1 0 1584 0 1 2970
box -8 -3 46 105
use INVX2  INVX2_204
timestamp 1682952543
transform 1 0 1624 0 1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_196
timestamp 1682952543
transform -1 0 1736 0 1 2970
box -8 -3 104 105
use AOI22X1  AOI22X1_104
timestamp 1682952543
transform -1 0 1776 0 1 2970
box -8 -3 46 105
use INVX2  INVX2_206
timestamp 1682952543
transform 1 0 1776 0 1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_105
timestamp 1682952543
transform -1 0 1832 0 1 2970
box -8 -3 46 105
use INVX2  INVX2_207
timestamp 1682952543
transform 1 0 1832 0 1 2970
box -9 -3 26 105
use FILL  FILL_825
timestamp 1682952543
transform 1 0 1848 0 1 2970
box -8 -3 16 105
use FILL  FILL_826
timestamp 1682952543
transform 1 0 1856 0 1 2970
box -8 -3 16 105
use FILL  FILL_827
timestamp 1682952543
transform 1 0 1864 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_106
timestamp 1682952543
transform -1 0 1912 0 1 2970
box -8 -3 46 105
use INVX2  INVX2_208
timestamp 1682952543
transform 1 0 1912 0 1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_197
timestamp 1682952543
transform -1 0 2024 0 1 2970
box -8 -3 104 105
use M3_M2  M3_M2_2748
timestamp 1682952543
transform 1 0 2084 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_198
timestamp 1682952543
transform 1 0 2024 0 1 2970
box -8 -3 104 105
use M3_M2  M3_M2_2749
timestamp 1682952543
transform 1 0 2220 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_199
timestamp 1682952543
transform 1 0 2120 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_209
timestamp 1682952543
transform 1 0 2216 0 1 2970
box -9 -3 26 105
use OAI22X1  OAI22X1_180
timestamp 1682952543
transform 1 0 2232 0 1 2970
box -8 -3 46 105
use FILL  FILL_828
timestamp 1682952543
transform 1 0 2272 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_181
timestamp 1682952543
transform 1 0 2280 0 1 2970
box -8 -3 46 105
use FILL  FILL_829
timestamp 1682952543
transform 1 0 2320 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_210
timestamp 1682952543
transform -1 0 2344 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_211
timestamp 1682952543
transform -1 0 2360 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_212
timestamp 1682952543
transform -1 0 2376 0 1 2970
box -9 -3 26 105
use M3_M2  M3_M2_2750
timestamp 1682952543
transform 1 0 2396 0 1 2975
box -3 -3 3 3
use OAI21X1  OAI21X1_40
timestamp 1682952543
transform 1 0 2376 0 1 2970
box -8 -3 34 105
use INVX2  INVX2_213
timestamp 1682952543
transform -1 0 2424 0 1 2970
box -9 -3 26 105
use M3_M2  M3_M2_2751
timestamp 1682952543
transform 1 0 2492 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_200
timestamp 1682952543
transform -1 0 2520 0 1 2970
box -8 -3 104 105
use FILL  FILL_830
timestamp 1682952543
transform 1 0 2520 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_201
timestamp 1682952543
transform -1 0 2624 0 1 2970
box -8 -3 104 105
use M3_M2  M3_M2_2752
timestamp 1682952543
transform 1 0 2724 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_202
timestamp 1682952543
transform 1 0 2624 0 1 2970
box -8 -3 104 105
use NOR2X1  NOR2X1_31
timestamp 1682952543
transform 1 0 2720 0 1 2970
box -8 -3 32 105
use FILL  FILL_831
timestamp 1682952543
transform 1 0 2744 0 1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_33
timestamp 1682952543
transform -1 0 2776 0 1 2970
box -8 -3 32 105
use FILL  FILL_832
timestamp 1682952543
transform 1 0 2776 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_32
timestamp 1682952543
transform 1 0 2784 0 1 2970
box -8 -3 32 105
use FILL  FILL_833
timestamp 1682952543
transform 1 0 2808 0 1 2970
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1682952543
transform -1 0 2840 0 1 2970
box -8 -3 32 105
use INVX2  INVX2_214
timestamp 1682952543
transform 1 0 2840 0 1 2970
box -9 -3 26 105
use INVX2  INVX2_215
timestamp 1682952543
transform 1 0 2856 0 1 2970
box -9 -3 26 105
use M3_M2  M3_M2_2753
timestamp 1682952543
transform 1 0 2900 0 1 2975
box -3 -3 3 3
use NAND2X1  NAND2X1_35
timestamp 1682952543
transform -1 0 2896 0 1 2970
box -8 -3 32 105
use INVX2  INVX2_216
timestamp 1682952543
transform 1 0 2896 0 1 2970
box -9 -3 26 105
use FILL  FILL_834
timestamp 1682952543
transform 1 0 2912 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_217
timestamp 1682952543
transform 1 0 2920 0 1 2970
box -9 -3 26 105
use FILL  FILL_835
timestamp 1682952543
transform 1 0 2936 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_218
timestamp 1682952543
transform 1 0 2944 0 1 2970
box -9 -3 26 105
use NAND3X1  NAND3X1_1
timestamp 1682952543
transform 1 0 2960 0 1 2970
box -8 -3 40 105
use FILL  FILL_836
timestamp 1682952543
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_837
timestamp 1682952543
transform 1 0 3000 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_219
timestamp 1682952543
transform 1 0 3008 0 1 2970
box -9 -3 26 105
use FILL  FILL_838
timestamp 1682952543
transform 1 0 3024 0 1 2970
box -8 -3 16 105
use FILL  FILL_839
timestamp 1682952543
transform 1 0 3032 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_2754
timestamp 1682952543
transform 1 0 3052 0 1 2975
box -3 -3 3 3
use FILL  FILL_840
timestamp 1682952543
transform 1 0 3040 0 1 2970
box -8 -3 16 105
use FILL  FILL_841
timestamp 1682952543
transform 1 0 3048 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_107
timestamp 1682952543
transform -1 0 3096 0 1 2970
box -8 -3 46 105
use FILL  FILL_842
timestamp 1682952543
transform 1 0 3096 0 1 2970
box -8 -3 16 105
use FILL  FILL_843
timestamp 1682952543
transform 1 0 3104 0 1 2970
box -8 -3 16 105
use FILL  FILL_844
timestamp 1682952543
transform 1 0 3112 0 1 2970
box -8 -3 16 105
use FILL  FILL_845
timestamp 1682952543
transform 1 0 3120 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_108
timestamp 1682952543
transform 1 0 3128 0 1 2970
box -8 -3 46 105
use FILL  FILL_846
timestamp 1682952543
transform 1 0 3168 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_2755
timestamp 1682952543
transform 1 0 3204 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_109
timestamp 1682952543
transform 1 0 3176 0 1 2970
box -8 -3 46 105
use NAND3X1  NAND3X1_2
timestamp 1682952543
transform 1 0 3216 0 1 2970
box -8 -3 40 105
use FILL  FILL_850
timestamp 1682952543
transform 1 0 3248 0 1 2970
box -8 -3 16 105
use FILL  FILL_852
timestamp 1682952543
transform 1 0 3256 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_2756
timestamp 1682952543
transform 1 0 3276 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_112
timestamp 1682952543
transform 1 0 3264 0 1 2970
box -8 -3 46 105
use M3_M2  M3_M2_2757
timestamp 1682952543
transform 1 0 3316 0 1 2975
box -3 -3 3 3
use FILL  FILL_854
timestamp 1682952543
transform 1 0 3304 0 1 2970
box -8 -3 16 105
use FILL  FILL_855
timestamp 1682952543
transform 1 0 3312 0 1 2970
box -8 -3 16 105
use FILL  FILL_856
timestamp 1682952543
transform 1 0 3320 0 1 2970
box -8 -3 16 105
use FILL  FILL_858
timestamp 1682952543
transform 1 0 3328 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_2758
timestamp 1682952543
transform 1 0 3356 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1682952543
transform 1 0 3372 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_113
timestamp 1682952543
transform 1 0 3336 0 1 2970
box -8 -3 46 105
use FILL  FILL_860
timestamp 1682952543
transform 1 0 3376 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_2760
timestamp 1682952543
transform 1 0 3396 0 1 2975
box -3 -3 3 3
use FILL  FILL_862
timestamp 1682952543
transform 1 0 3384 0 1 2970
box -8 -3 16 105
use FILL  FILL_864
timestamp 1682952543
transform 1 0 3392 0 1 2970
box -8 -3 16 105
use FILL  FILL_865
timestamp 1682952543
transform 1 0 3400 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_34
timestamp 1682952543
transform -1 0 3432 0 1 2970
box -8 -3 32 105
use FILL  FILL_866
timestamp 1682952543
transform 1 0 3432 0 1 2970
box -8 -3 16 105
use FILL  FILL_867
timestamp 1682952543
transform 1 0 3440 0 1 2970
box -8 -3 16 105
use FILL  FILL_868
timestamp 1682952543
transform 1 0 3448 0 1 2970
box -8 -3 16 105
use FILL  FILL_869
timestamp 1682952543
transform 1 0 3456 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_2761
timestamp 1682952543
transform 1 0 3476 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1682952543
transform 1 0 3492 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_115
timestamp 1682952543
transform 1 0 3464 0 1 2970
box -8 -3 46 105
use FILL  FILL_870
timestamp 1682952543
transform 1 0 3504 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_225
timestamp 1682952543
transform -1 0 3528 0 1 2970
box -9 -3 26 105
use FAX1  FAX1_2
timestamp 1682952543
transform 1 0 3528 0 1 2970
box -5 -3 126 105
use FILL  FILL_871
timestamp 1682952543
transform 1 0 3648 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_2763
timestamp 1682952543
transform 1 0 3756 0 1 2975
box -3 -3 3 3
use FAX1  FAX1_3
timestamp 1682952543
transform 1 0 3656 0 1 2970
box -5 -3 126 105
use M3_M2  M3_M2_2764
timestamp 1682952543
transform 1 0 3812 0 1 2975
box -3 -3 3 3
use FAX1  FAX1_4
timestamp 1682952543
transform -1 0 3896 0 1 2970
box -5 -3 126 105
use FILL  FILL_872
timestamp 1682952543
transform 1 0 3896 0 1 2970
box -8 -3 16 105
use FAX1  FAX1_5
timestamp 1682952543
transform 1 0 3904 0 1 2970
box -5 -3 126 105
use FILL  FILL_877
timestamp 1682952543
transform 1 0 4024 0 1 2970
box -8 -3 16 105
use FAX1  FAX1_6
timestamp 1682952543
transform 1 0 4032 0 1 2970
box -5 -3 126 105
use top_level_VIA0  top_level_VIA0_23
timestamp 1682952543
transform 1 0 4177 0 1 2970
box -10 -3 10 3
use M3_M2  M3_M2_2826
timestamp 1682952543
transform 1 0 148 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1682952543
transform 1 0 140 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2851
timestamp 1682952543
transform 1 0 148 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1682952543
transform 1 0 132 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1682952543
transform 1 0 140 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2926
timestamp 1682952543
transform 1 0 148 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1682952543
transform 1 0 164 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2852
timestamp 1682952543
transform 1 0 164 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2873
timestamp 1682952543
transform 1 0 172 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2853
timestamp 1682952543
transform 1 0 188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1682952543
transform 1 0 172 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2927
timestamp 1682952543
transform 1 0 172 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1682952543
transform 1 0 204 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_2974
timestamp 1682952543
transform 1 0 204 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2766
timestamp 1682952543
transform 1 0 252 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2827
timestamp 1682952543
transform 1 0 220 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2828
timestamp 1682952543
transform 1 0 260 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2829
timestamp 1682952543
transform 1 0 300 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2854
timestamp 1682952543
transform 1 0 220 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2899
timestamp 1682952543
transform 1 0 220 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_2855
timestamp 1682952543
transform 1 0 308 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2975
timestamp 1682952543
transform 1 0 244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1682952543
transform 1 0 300 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1682952543
transform 1 0 340 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1682952543
transform 1 0 348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2977
timestamp 1682952543
transform 1 0 316 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1682952543
transform 1 0 332 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2900
timestamp 1682952543
transform 1 0 340 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_2979
timestamp 1682952543
transform 1 0 356 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2767
timestamp 1682952543
transform 1 0 420 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1682952543
transform 1 0 468 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2795
timestamp 1682952543
transform 1 0 484 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2768
timestamp 1682952543
transform 1 0 612 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1682952543
transform 1 0 500 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2831
timestamp 1682952543
transform 1 0 596 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2858
timestamp 1682952543
transform 1 0 380 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1682952543
transform 1 0 468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2860
timestamp 1682952543
transform 1 0 484 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1682952543
transform 1 0 500 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1682952543
transform 1 0 516 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2863
timestamp 1682952543
transform 1 0 604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1682952543
transform 1 0 364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2981
timestamp 1682952543
transform 1 0 404 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2901
timestamp 1682952543
transform 1 0 452 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_2982
timestamp 1682952543
transform 1 0 460 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2983
timestamp 1682952543
transform 1 0 476 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2984
timestamp 1682952543
transform 1 0 500 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1682952543
transform 1 0 556 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2986
timestamp 1682952543
transform 1 0 596 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2928
timestamp 1682952543
transform 1 0 364 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2929
timestamp 1682952543
transform 1 0 404 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1682952543
transform 1 0 460 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1682952543
transform 1 0 444 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2930
timestamp 1682952543
transform 1 0 500 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1682952543
transform 1 0 508 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2902
timestamp 1682952543
transform 1 0 604 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1682952543
transform 1 0 604 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3018
timestamp 1682952543
transform 1 0 524 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3019
timestamp 1682952543
transform 1 0 556 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2796
timestamp 1682952543
transform 1 0 628 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2838
timestamp 1682952543
transform 1 0 628 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_2832
timestamp 1682952543
transform 1 0 644 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2839
timestamp 1682952543
transform 1 0 692 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1682952543
transform 1 0 628 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2865
timestamp 1682952543
transform 1 0 644 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1682952543
transform 1 0 668 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2987
timestamp 1682952543
transform 1 0 620 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2903
timestamp 1682952543
transform 1 0 636 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2874
timestamp 1682952543
transform 1 0 676 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2867
timestamp 1682952543
transform 1 0 684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1682952543
transform 1 0 700 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1682952543
transform 1 0 644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1682952543
transform 1 0 652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1682952543
transform 1 0 676 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2932
timestamp 1682952543
transform 1 0 652 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2933
timestamp 1682952543
transform 1 0 692 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_2869
timestamp 1682952543
transform 1 0 716 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2769
timestamp 1682952543
transform 1 0 732 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2875
timestamp 1682952543
transform 1 0 732 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2870
timestamp 1682952543
transform 1 0 740 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2991
timestamp 1682952543
transform 1 0 732 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1682952543
transform 1 0 740 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2979
timestamp 1682952543
transform 1 0 724 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2770
timestamp 1682952543
transform 1 0 780 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2833
timestamp 1682952543
transform 1 0 788 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2834
timestamp 1682952543
transform 1 0 828 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2871
timestamp 1682952543
transform 1 0 828 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1682952543
transform 1 0 796 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2934
timestamp 1682952543
transform 1 0 764 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1682952543
transform 1 0 828 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3020
timestamp 1682952543
transform 1 0 804 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1682952543
transform 1 0 852 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2797
timestamp 1682952543
transform 1 0 860 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2840
timestamp 1682952543
transform 1 0 852 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1682952543
transform 1 0 844 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2772
timestamp 1682952543
transform 1 0 892 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1682952543
transform 1 0 964 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1682952543
transform 1 0 980 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2835
timestamp 1682952543
transform 1 0 908 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2873
timestamp 1682952543
transform 1 0 884 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1682952543
transform 1 0 876 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2995
timestamp 1682952543
transform 1 0 884 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2935
timestamp 1682952543
transform 1 0 884 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3006
timestamp 1682952543
transform 1 0 876 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_2874
timestamp 1682952543
transform 1 0 908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1682952543
transform 1 0 948 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2936
timestamp 1682952543
transform 1 0 956 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1682952543
transform 1 0 940 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3021
timestamp 1682952543
transform 1 0 908 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1682952543
transform 1 0 972 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_2997
timestamp 1682952543
transform 1 0 996 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2937
timestamp 1682952543
transform 1 0 996 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1682952543
transform 1 0 996 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1682952543
transform 1 0 1020 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2776
timestamp 1682952543
transform 1 0 1092 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2836
timestamp 1682952543
transform 1 0 1012 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2875
timestamp 1682952543
transform 1 0 1012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2998
timestamp 1682952543
transform 1 0 1036 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2938
timestamp 1682952543
transform 1 0 1084 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1682952543
transform 1 0 1084 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1682952543
transform 1 0 1092 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2777
timestamp 1682952543
transform 1 0 1124 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1682952543
transform 1 0 1196 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2838
timestamp 1682952543
transform 1 0 1212 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2798
timestamp 1682952543
transform 1 0 1284 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2839
timestamp 1682952543
transform 1 0 1276 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2876
timestamp 1682952543
transform 1 0 1116 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1682952543
transform 1 0 1124 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2878
timestamp 1682952543
transform 1 0 1140 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1682952543
transform 1 0 1148 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2880
timestamp 1682952543
transform 1 0 1164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2881
timestamp 1682952543
transform 1 0 1252 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2882
timestamp 1682952543
transform 1 0 1268 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1682952543
transform 1 0 1284 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2884
timestamp 1682952543
transform 1 0 1292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1682952543
transform 1 0 1108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1682952543
transform 1 0 1132 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2939
timestamp 1682952543
transform 1 0 1140 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2876
timestamp 1682952543
transform 1 0 1300 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1682952543
transform 1 0 1356 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2840
timestamp 1682952543
transform 1 0 1340 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2885
timestamp 1682952543
transform 1 0 1308 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1682952543
transform 1 0 1332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2887
timestamp 1682952543
transform 1 0 1340 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2877
timestamp 1682952543
transform 1 0 1348 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2888
timestamp 1682952543
transform 1 0 1356 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2889
timestamp 1682952543
transform 1 0 1372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1682952543
transform 1 0 1196 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1682952543
transform 1 0 1244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3003
timestamp 1682952543
transform 1 0 1260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1682952543
transform 1 0 1284 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3005
timestamp 1682952543
transform 1 0 1300 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3006
timestamp 1682952543
transform 1 0 1324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1682952543
transform 1 0 1332 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1682952543
transform 1 0 1348 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1682952543
transform 1 0 1364 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2940
timestamp 1682952543
transform 1 0 1244 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2984
timestamp 1682952543
transform 1 0 1252 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3024
timestamp 1682952543
transform 1 0 1148 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3025
timestamp 1682952543
transform 1 0 1180 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3026
timestamp 1682952543
transform 1 0 1228 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1682952543
transform 1 0 1292 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1682952543
transform 1 0 1316 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1682952543
transform 1 0 1332 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3027
timestamp 1682952543
transform 1 0 1260 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1682952543
transform 1 0 1324 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3028
timestamp 1682952543
transform 1 0 1300 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1682952543
transform 1 0 1388 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2878
timestamp 1682952543
transform 1 0 1380 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2879
timestamp 1682952543
transform 1 0 1404 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2890
timestamp 1682952543
transform 1 0 1468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1682952543
transform 1 0 1484 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3010
timestamp 1682952543
transform 1 0 1380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1682952543
transform 1 0 1388 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1682952543
transform 1 0 1420 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2944
timestamp 1682952543
transform 1 0 1380 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1682952543
transform 1 0 1420 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2986
timestamp 1682952543
transform 1 0 1484 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1682952543
transform 1 0 1556 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1682952543
transform 1 0 1548 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2892
timestamp 1682952543
transform 1 0 1508 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1682952543
transform 1 0 1524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2894
timestamp 1682952543
transform 1 0 1540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1682952543
transform 1 0 1548 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1682952543
transform 1 0 1564 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2880
timestamp 1682952543
transform 1 0 1572 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2897
timestamp 1682952543
transform 1 0 1580 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1682952543
transform 1 0 1588 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2899
timestamp 1682952543
transform 1 0 1612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2900
timestamp 1682952543
transform 1 0 1620 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1682952543
transform 1 0 1500 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1682952543
transform 1 0 1508 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2904
timestamp 1682952543
transform 1 0 1524 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3015
timestamp 1682952543
transform 1 0 1532 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2905
timestamp 1682952543
transform 1 0 1540 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3016
timestamp 1682952543
transform 1 0 1548 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1682952543
transform 1 0 1572 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2946
timestamp 1682952543
transform 1 0 1516 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2906
timestamp 1682952543
transform 1 0 1580 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3018
timestamp 1682952543
transform 1 0 1588 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1682952543
transform 1 0 1604 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2907
timestamp 1682952543
transform 1 0 1612 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3020
timestamp 1682952543
transform 1 0 1628 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2947
timestamp 1682952543
transform 1 0 1588 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1682952543
transform 1 0 1508 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1682952543
transform 1 0 1548 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3029
timestamp 1682952543
transform 1 0 1532 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3007
timestamp 1682952543
transform 1 0 1564 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3008
timestamp 1682952543
transform 1 0 1580 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3030
timestamp 1682952543
transform 1 0 1572 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2842
timestamp 1682952543
transform 1 0 1740 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2843
timestamp 1682952543
transform 1 0 1820 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2901
timestamp 1682952543
transform 1 0 1724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1682952543
transform 1 0 1636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1682952543
transform 1 0 1644 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2908
timestamp 1682952543
transform 1 0 1652 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2802
timestamp 1682952543
transform 1 0 1860 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2902
timestamp 1682952543
transform 1 0 1820 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1682952543
transform 1 0 1836 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1682952543
transform 1 0 1844 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2881
timestamp 1682952543
transform 1 0 1852 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2905
timestamp 1682952543
transform 1 0 1860 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2906
timestamp 1682952543
transform 1 0 1876 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2803
timestamp 1682952543
transform 1 0 1980 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2804
timestamp 1682952543
transform 1 0 2012 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2805
timestamp 1682952543
transform 1 0 2044 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1682952543
transform 1 0 1884 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1682952543
transform 1 0 1900 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3023
timestamp 1682952543
transform 1 0 1676 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3024
timestamp 1682952543
transform 1 0 1740 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1682952543
transform 1 0 1780 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3026
timestamp 1682952543
transform 1 0 1836 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1682952543
transform 1 0 1852 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2948
timestamp 1682952543
transform 1 0 1636 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2949
timestamp 1682952543
transform 1 0 1676 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3031
timestamp 1682952543
transform 1 0 1716 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1682952543
transform 1 0 1860 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3028
timestamp 1682952543
transform 1 0 1868 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2910
timestamp 1682952543
transform 1 0 1876 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_2907
timestamp 1682952543
transform 1 0 1900 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2846
timestamp 1682952543
transform 1 0 1996 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2847
timestamp 1682952543
transform 1 0 2036 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2908
timestamp 1682952543
transform 1 0 1996 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2778
timestamp 1682952543
transform 1 0 2196 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2779
timestamp 1682952543
transform 1 0 2284 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2806
timestamp 1682952543
transform 1 0 2172 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2807
timestamp 1682952543
transform 1 0 2220 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2808
timestamp 1682952543
transform 1 0 2276 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1682952543
transform 1 0 2164 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2882
timestamp 1682952543
transform 1 0 2140 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2909
timestamp 1682952543
transform 1 0 2164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1682952543
transform 1 0 1884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1682952543
transform 1 0 1924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3031
timestamp 1682952543
transform 1 0 1980 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1682952543
transform 1 0 2020 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1682952543
transform 1 0 2076 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1682952543
transform 1 0 2084 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1682952543
transform 1 0 2140 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2950
timestamp 1682952543
transform 1 0 1860 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2989
timestamp 1682952543
transform 1 0 1836 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3009
timestamp 1682952543
transform 1 0 1828 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_2951
timestamp 1682952543
transform 1 0 1884 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1682952543
transform 1 0 1924 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1682952543
transform 1 0 1948 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1682952543
transform 1 0 1932 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1682952543
transform 1 0 2020 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2955
timestamp 1682952543
transform 1 0 2068 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3010
timestamp 1682952543
transform 1 0 2116 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1682952543
transform 1 0 2100 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3033
timestamp 1682952543
transform 1 0 2124 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3034
timestamp 1682952543
transform 1 0 2156 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2849
timestamp 1682952543
transform 1 0 2188 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2910
timestamp 1682952543
transform 1 0 2188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2911
timestamp 1682952543
transform 1 0 2276 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1682952543
transform 1 0 2236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3037
timestamp 1682952543
transform 1 0 2276 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2956
timestamp 1682952543
transform 1 0 2276 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3011
timestamp 1682952543
transform 1 0 2236 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1682952543
transform 1 0 2212 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3036
timestamp 1682952543
transform 1 0 2244 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_2850
timestamp 1682952543
transform 1 0 2292 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2780
timestamp 1682952543
transform 1 0 2332 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_2912
timestamp 1682952543
transform 1 0 2292 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2883
timestamp 1682952543
transform 1 0 2308 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2781
timestamp 1682952543
transform 1 0 2388 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2782
timestamp 1682952543
transform 1 0 2444 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2783
timestamp 1682952543
transform 1 0 2484 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1682952543
transform 1 0 2372 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2810
timestamp 1682952543
transform 1 0 2404 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2811
timestamp 1682952543
transform 1 0 2428 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2851
timestamp 1682952543
transform 1 0 2348 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2852
timestamp 1682952543
transform 1 0 2364 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2913
timestamp 1682952543
transform 1 0 2316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2914
timestamp 1682952543
transform 1 0 2332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2915
timestamp 1682952543
transform 1 0 2340 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2916
timestamp 1682952543
transform 1 0 2364 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1682952543
transform 1 0 2300 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1682952543
transform 1 0 2308 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2911
timestamp 1682952543
transform 1 0 2316 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3040
timestamp 1682952543
transform 1 0 2324 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1682952543
transform 1 0 2292 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2991
timestamp 1682952543
transform 1 0 2292 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1682952543
transform 1 0 2404 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1682952543
transform 1 0 2524 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2917
timestamp 1682952543
transform 1 0 2372 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2918
timestamp 1682952543
transform 1 0 2396 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1682952543
transform 1 0 2412 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3041
timestamp 1682952543
transform 1 0 2348 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2957
timestamp 1682952543
transform 1 0 2332 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1682952543
transform 1 0 2372 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2884
timestamp 1682952543
transform 1 0 2420 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2920
timestamp 1682952543
transform 1 0 2428 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2885
timestamp 1682952543
transform 1 0 2444 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2921
timestamp 1682952543
transform 1 0 2524 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1682952543
transform 1 0 2388 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1682952543
transform 1 0 2404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3106
timestamp 1682952543
transform 1 0 2364 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1682952543
transform 1 0 2372 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2958
timestamp 1682952543
transform 1 0 2388 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2913
timestamp 1682952543
transform 1 0 2412 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3044
timestamp 1682952543
transform 1 0 2420 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1682952543
transform 1 0 2436 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1682952543
transform 1 0 2444 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2992
timestamp 1682952543
transform 1 0 2348 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1682952543
transform 1 0 2372 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1682952543
transform 1 0 2396 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1682952543
transform 1 0 2340 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1682952543
transform 1 0 2460 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3047
timestamp 1682952543
transform 1 0 2500 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2959
timestamp 1682952543
transform 1 0 2500 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2784
timestamp 1682952543
transform 1 0 2596 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2855
timestamp 1682952543
transform 1 0 2548 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2856
timestamp 1682952543
transform 1 0 2612 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2922
timestamp 1682952543
transform 1 0 2548 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2785
timestamp 1682952543
transform 1 0 2660 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2857
timestamp 1682952543
transform 1 0 2716 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2923
timestamp 1682952543
transform 1 0 2716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3048
timestamp 1682952543
transform 1 0 2572 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1682952543
transform 1 0 2628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1682952543
transform 1 0 2636 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3051
timestamp 1682952543
transform 1 0 2692 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2995
timestamp 1682952543
transform 1 0 2572 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1682952543
transform 1 0 2716 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1682952543
transform 1 0 2812 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2841
timestamp 1682952543
transform 1 0 2828 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1682952543
transform 1 0 2812 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2886
timestamp 1682952543
transform 1 0 2828 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1682952543
transform 1 0 2844 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2925
timestamp 1682952543
transform 1 0 2836 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2926
timestamp 1682952543
transform 1 0 2844 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2927
timestamp 1682952543
transform 1 0 2852 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1682952543
transform 1 0 2732 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3053
timestamp 1682952543
transform 1 0 2764 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2996
timestamp 1682952543
transform 1 0 2692 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1682952543
transform 1 0 2812 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2997
timestamp 1682952543
transform 1 0 2764 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1682952543
transform 1 0 2836 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1682952543
transform 1 0 2868 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2928
timestamp 1682952543
transform 1 0 2876 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3054
timestamp 1682952543
transform 1 0 2868 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2917
timestamp 1682952543
transform 1 0 2876 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3108
timestamp 1682952543
transform 1 0 2868 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3013
timestamp 1682952543
transform 1 0 2868 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_2929
timestamp 1682952543
transform 1 0 2892 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3055
timestamp 1682952543
transform 1 0 2900 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1682952543
transform 1 0 2900 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2918
timestamp 1682952543
transform 1 0 2924 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_2930
timestamp 1682952543
transform 1 0 2956 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3056
timestamp 1682952543
transform 1 0 2932 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3110
timestamp 1682952543
transform 1 0 2916 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1682952543
transform 1 0 2924 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3112
timestamp 1682952543
transform 1 0 2948 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1682952543
transform 1 0 2924 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_2998
timestamp 1682952543
transform 1 0 2940 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1682952543
transform 1 0 3004 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2931
timestamp 1682952543
transform 1 0 3004 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2919
timestamp 1682952543
transform 1 0 3020 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1682952543
transform 1 0 3052 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2889
timestamp 1682952543
transform 1 0 3068 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3057
timestamp 1682952543
transform 1 0 3028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1682952543
transform 1 0 3052 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3059
timestamp 1682952543
transform 1 0 3068 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3113
timestamp 1682952543
transform 1 0 3028 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1682952543
transform 1 0 3036 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2961
timestamp 1682952543
transform 1 0 3052 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3115
timestamp 1682952543
transform 1 0 3060 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2999
timestamp 1682952543
transform 1 0 3036 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3128
timestamp 1682952543
transform 1 0 3052 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_2786
timestamp 1682952543
transform 1 0 3116 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1682952543
transform 1 0 3100 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2861
timestamp 1682952543
transform 1 0 3084 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2842
timestamp 1682952543
transform 1 0 3100 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2932
timestamp 1682952543
transform 1 0 3076 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2933
timestamp 1682952543
transform 1 0 3084 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2890
timestamp 1682952543
transform 1 0 3108 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1682952543
transform 1 0 3180 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2813
timestamp 1682952543
transform 1 0 3188 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2862
timestamp 1682952543
transform 1 0 3156 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2863
timestamp 1682952543
transform 1 0 3172 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2934
timestamp 1682952543
transform 1 0 3116 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2935
timestamp 1682952543
transform 1 0 3132 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2936
timestamp 1682952543
transform 1 0 3148 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3060
timestamp 1682952543
transform 1 0 3092 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1682952543
transform 1 0 3100 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2962
timestamp 1682952543
transform 1 0 3100 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3062
timestamp 1682952543
transform 1 0 3124 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3063
timestamp 1682952543
transform 1 0 3140 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3000
timestamp 1682952543
transform 1 0 3124 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_2937
timestamp 1682952543
transform 1 0 3164 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2891
timestamp 1682952543
transform 1 0 3172 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2938
timestamp 1682952543
transform 1 0 3188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3064
timestamp 1682952543
transform 1 0 3156 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3065
timestamp 1682952543
transform 1 0 3172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2939
timestamp 1682952543
transform 1 0 3196 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1682952543
transform 1 0 3204 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2963
timestamp 1682952543
transform 1 0 3196 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3001
timestamp 1682952543
transform 1 0 3204 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1682952543
transform 1 0 3196 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3116
timestamp 1682952543
transform 1 0 3212 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2814
timestamp 1682952543
transform 1 0 3236 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1682952543
transform 1 0 3228 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3038
timestamp 1682952543
transform 1 0 3220 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3067
timestamp 1682952543
transform 1 0 3244 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1682952543
transform 1 0 3252 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2964
timestamp 1682952543
transform 1 0 3252 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2815
timestamp 1682952543
transform 1 0 3260 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2843
timestamp 1682952543
transform 1 0 3260 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2940
timestamp 1682952543
transform 1 0 3268 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2788
timestamp 1682952543
transform 1 0 3300 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2816
timestamp 1682952543
transform 1 0 3292 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1682952543
transform 1 0 3300 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2941
timestamp 1682952543
transform 1 0 3292 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1682952543
transform 1 0 3300 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2920
timestamp 1682952543
transform 1 0 3308 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3117
timestamp 1682952543
transform 1 0 3292 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3118
timestamp 1682952543
transform 1 0 3300 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_2942
timestamp 1682952543
transform 1 0 3332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3070
timestamp 1682952543
transform 1 0 3324 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2789
timestamp 1682952543
transform 1 0 3348 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1682952543
transform 1 0 3364 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2817
timestamp 1682952543
transform 1 0 3380 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2943
timestamp 1682952543
transform 1 0 3348 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2944
timestamp 1682952543
transform 1 0 3364 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2945
timestamp 1682952543
transform 1 0 3372 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2921
timestamp 1682952543
transform 1 0 3340 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3071
timestamp 1682952543
transform 1 0 3356 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2922
timestamp 1682952543
transform 1 0 3364 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3072
timestamp 1682952543
transform 1 0 3380 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2946
timestamp 1682952543
transform 1 0 3388 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2965
timestamp 1682952543
transform 1 0 3380 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_2844
timestamp 1682952543
transform 1 0 3420 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_2892
timestamp 1682952543
transform 1 0 3444 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1682952543
transform 1 0 3468 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2947
timestamp 1682952543
transform 1 0 3460 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3073
timestamp 1682952543
transform 1 0 3420 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3074
timestamp 1682952543
transform 1 0 3444 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2966
timestamp 1682952543
transform 1 0 3404 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2967
timestamp 1682952543
transform 1 0 3420 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3119
timestamp 1682952543
transform 1 0 3428 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3075
timestamp 1682952543
transform 1 0 3468 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3076
timestamp 1682952543
transform 1 0 3492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1682952543
transform 1 0 3452 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3129
timestamp 1682952543
transform 1 0 3436 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_2968
timestamp 1682952543
transform 1 0 3468 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3121
timestamp 1682952543
transform 1 0 3476 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1682952543
transform 1 0 3492 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3002
timestamp 1682952543
transform 1 0 3468 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_2948
timestamp 1682952543
transform 1 0 3516 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2969
timestamp 1682952543
transform 1 0 3508 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3130
timestamp 1682952543
transform 1 0 3508 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_2819
timestamp 1682952543
transform 1 0 3532 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2790
timestamp 1682952543
transform 1 0 3588 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_2845
timestamp 1682952543
transform 1 0 3556 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_2867
timestamp 1682952543
transform 1 0 3564 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1682952543
transform 1 0 3636 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_2820
timestamp 1682952543
transform 1 0 3628 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2868
timestamp 1682952543
transform 1 0 3612 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2949
timestamp 1682952543
transform 1 0 3532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2950
timestamp 1682952543
transform 1 0 3540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1682952543
transform 1 0 3564 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1682952543
transform 1 0 3588 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2953
timestamp 1682952543
transform 1 0 3596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2954
timestamp 1682952543
transform 1 0 3604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1682952543
transform 1 0 3524 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2923
timestamp 1682952543
transform 1 0 3532 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3078
timestamp 1682952543
transform 1 0 3556 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3079
timestamp 1682952543
transform 1 0 3564 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1682952543
transform 1 0 3580 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2970
timestamp 1682952543
transform 1 0 3556 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_2955
timestamp 1682952543
transform 1 0 3636 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3081
timestamp 1682952543
transform 1 0 3636 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2821
timestamp 1682952543
transform 1 0 3660 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2846
timestamp 1682952543
transform 1 0 3660 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_2822
timestamp 1682952543
transform 1 0 3700 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_2893
timestamp 1682952543
transform 1 0 3660 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2956
timestamp 1682952543
transform 1 0 3668 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2894
timestamp 1682952543
transform 1 0 3676 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2957
timestamp 1682952543
transform 1 0 3684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1682952543
transform 1 0 3700 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1682952543
transform 1 0 3716 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1682952543
transform 1 0 3724 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3082
timestamp 1682952543
transform 1 0 3660 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3123
timestamp 1682952543
transform 1 0 3612 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2971
timestamp 1682952543
transform 1 0 3636 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1682952543
transform 1 0 3652 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3131
timestamp 1682952543
transform 1 0 3628 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_3014
timestamp 1682952543
transform 1 0 3644 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_3083
timestamp 1682952543
transform 1 0 3676 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1682952543
transform 1 0 3692 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3085
timestamp 1682952543
transform 1 0 3708 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1682952543
transform 1 0 3716 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3003
timestamp 1682952543
transform 1 0 3708 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1682952543
transform 1 0 3716 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_2823
timestamp 1682952543
transform 1 0 3748 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2847
timestamp 1682952543
transform 1 0 3748 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1682952543
transform 1 0 3764 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1682952543
transform 1 0 3780 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2824
timestamp 1682952543
transform 1 0 3812 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2848
timestamp 1682952543
transform 1 0 3828 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2963
timestamp 1682952543
transform 1 0 3812 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3087
timestamp 1682952543
transform 1 0 3772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3088
timestamp 1682952543
transform 1 0 3788 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3089
timestamp 1682952543
transform 1 0 3796 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2973
timestamp 1682952543
transform 1 0 3788 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3124
timestamp 1682952543
transform 1 0 3796 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2974
timestamp 1682952543
transform 1 0 3804 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3004
timestamp 1682952543
transform 1 0 3796 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1682952543
transform 1 0 3796 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_3090
timestamp 1682952543
transform 1 0 3828 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1682952543
transform 1 0 3836 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3005
timestamp 1682952543
transform 1 0 3828 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1682952543
transform 1 0 3844 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2849
timestamp 1682952543
transform 1 0 3852 0 1 2945
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1682952543
transform 1 0 3844 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2924
timestamp 1682952543
transform 1 0 3844 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3092
timestamp 1682952543
transform 1 0 3852 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2792
timestamp 1682952543
transform 1 0 3876 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_2965
timestamp 1682952543
transform 1 0 3876 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1682952543
transform 1 0 3884 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2925
timestamp 1682952543
transform 1 0 3892 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_2870
timestamp 1682952543
transform 1 0 3924 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_2850
timestamp 1682952543
transform 1 0 3932 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_2895
timestamp 1682952543
transform 1 0 3908 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3094
timestamp 1682952543
transform 1 0 3908 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1682952543
transform 1 0 3940 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2825
timestamp 1682952543
transform 1 0 3996 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_2967
timestamp 1682952543
transform 1 0 3972 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1682952543
transform 1 0 3996 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3095
timestamp 1682952543
transform 1 0 3948 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1682952543
transform 1 0 3956 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1682952543
transform 1 0 3964 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3098
timestamp 1682952543
transform 1 0 3972 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1682952543
transform 1 0 3988 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2975
timestamp 1682952543
transform 1 0 3972 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3100
timestamp 1682952543
transform 1 0 4012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1682952543
transform 1 0 4020 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_2871
timestamp 1682952543
transform 1 0 4052 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_2896
timestamp 1682952543
transform 1 0 4044 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_2970
timestamp 1682952543
transform 1 0 4052 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3101
timestamp 1682952543
transform 1 0 4028 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3102
timestamp 1682952543
transform 1 0 4044 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_2976
timestamp 1682952543
transform 1 0 4028 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3125
timestamp 1682952543
transform 1 0 4068 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_2897
timestamp 1682952543
transform 1 0 4076 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3103
timestamp 1682952543
transform 1 0 4076 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1682952543
transform 1 0 4092 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3126
timestamp 1682952543
transform 1 0 4108 0 1 2915
box -2 -2 2 2
use M2_M1  M2_M1_3132
timestamp 1682952543
transform 1 0 4100 0 1 2905
box -2 -2 2 2
use M3_M2  M3_M2_2898
timestamp 1682952543
transform 1 0 4140 0 1 2935
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_24
timestamp 1682952543
transform 1 0 24 0 1 2870
box -10 -3 10 3
use FILL  FILL_778
timestamp 1682952543
transform 1 0 72 0 -1 2970
box -8 -3 16 105
use FILL  FILL_779
timestamp 1682952543
transform 1 0 80 0 -1 2970
box -8 -3 16 105
use FILL  FILL_780
timestamp 1682952543
transform 1 0 88 0 -1 2970
box -8 -3 16 105
use FILL  FILL_781
timestamp 1682952543
transform 1 0 96 0 -1 2970
box -8 -3 16 105
use FILL  FILL_782
timestamp 1682952543
transform 1 0 104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_783
timestamp 1682952543
transform 1 0 112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_784
timestamp 1682952543
transform 1 0 120 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_190
timestamp 1682952543
transform -1 0 144 0 -1 2970
box -9 -3 26 105
use FILL  FILL_785
timestamp 1682952543
transform 1 0 144 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_88
timestamp 1682952543
transform -1 0 192 0 -1 2970
box -8 -3 46 105
use FILL  FILL_786
timestamp 1682952543
transform 1 0 192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_814
timestamp 1682952543
transform 1 0 200 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_188
timestamp 1682952543
transform 1 0 208 0 -1 2970
box -8 -3 104 105
use FILL  FILL_815
timestamp 1682952543
transform 1 0 304 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_100
timestamp 1682952543
transform 1 0 312 0 -1 2970
box -8 -3 46 105
use INVX2  INVX2_201
timestamp 1682952543
transform 1 0 352 0 -1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_189
timestamp 1682952543
transform 1 0 368 0 -1 2970
box -8 -3 104 105
use OAI22X1  OAI22X1_174
timestamp 1682952543
transform -1 0 504 0 -1 2970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_190
timestamp 1682952543
transform 1 0 504 0 -1 2970
box -8 -3 104 105
use M3_M2  M3_M2_3039
timestamp 1682952543
transform 1 0 620 0 1 2875
box -3 -3 3 3
use BUFX2  BUFX2_16
timestamp 1682952543
transform -1 0 624 0 -1 2970
box -5 -3 28 105
use NOR2X1  NOR2X1_28
timestamp 1682952543
transform 1 0 624 0 -1 2970
box -8 -3 32 105
use OAI22X1  OAI22X1_175
timestamp 1682952543
transform 1 0 648 0 -1 2970
box -8 -3 46 105
use NOR2X1  NOR2X1_29
timestamp 1682952543
transform 1 0 688 0 -1 2970
box -8 -3 32 105
use FILL  FILL_816
timestamp 1682952543
transform 1 0 712 0 -1 2970
box -8 -3 16 105
use FILL  FILL_817
timestamp 1682952543
transform 1 0 720 0 -1 2970
box -8 -3 16 105
use FILL  FILL_818
timestamp 1682952543
transform 1 0 728 0 -1 2970
box -8 -3 16 105
use FILL  FILL_819
timestamp 1682952543
transform 1 0 736 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_191
timestamp 1682952543
transform -1 0 840 0 -1 2970
box -8 -3 104 105
use FILL  FILL_820
timestamp 1682952543
transform 1 0 840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_821
timestamp 1682952543
transform 1 0 848 0 -1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_30
timestamp 1682952543
transform 1 0 856 0 -1 2970
box -8 -3 32 105
use INVX2  INVX2_202
timestamp 1682952543
transform 1 0 880 0 -1 2970
box -9 -3 26 105
use M3_M2  M3_M2_3040
timestamp 1682952543
transform 1 0 956 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_192
timestamp 1682952543
transform 1 0 896 0 -1 2970
box -8 -3 104 105
use FILL  FILL_822
timestamp 1682952543
transform 1 0 992 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3041
timestamp 1682952543
transform 1 0 1036 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_193
timestamp 1682952543
transform 1 0 1000 0 -1 2970
box -8 -3 104 105
use FILL  FILL_823
timestamp 1682952543
transform 1 0 1096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_824
timestamp 1682952543
transform 1 0 1104 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_101
timestamp 1682952543
transform 1 0 1112 0 -1 2970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_194
timestamp 1682952543
transform 1 0 1152 0 -1 2970
box -8 -3 104 105
use M3_M2  M3_M2_3042
timestamp 1682952543
transform 1 0 1276 0 1 2875
box -3 -3 3 3
use OAI22X1  OAI22X1_176
timestamp 1682952543
transform -1 0 1288 0 -1 2970
box -8 -3 46 105
use M3_M2  M3_M2_3043
timestamp 1682952543
transform 1 0 1308 0 1 2875
box -3 -3 3 3
use OAI22X1  OAI22X1_177
timestamp 1682952543
transform -1 0 1328 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_102
timestamp 1682952543
transform 1 0 1328 0 -1 2970
box -8 -3 46 105
use INVX2  INVX2_203
timestamp 1682952543
transform 1 0 1368 0 -1 2970
box -9 -3 26 105
use M3_M2  M3_M2_3044
timestamp 1682952543
transform 1 0 1444 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_195
timestamp 1682952543
transform -1 0 1480 0 -1 2970
box -8 -3 104 105
use M3_M2  M3_M2_3045
timestamp 1682952543
transform 1 0 1500 0 1 2875
box -3 -3 3 3
use BUFX2  BUFX2_17
timestamp 1682952543
transform -1 0 1504 0 -1 2970
box -5 -3 28 105
use OAI22X1  OAI22X1_178
timestamp 1682952543
transform 1 0 1504 0 -1 2970
box -8 -3 46 105
use OAI22X1  OAI22X1_179
timestamp 1682952543
transform 1 0 1544 0 -1 2970
box -8 -3 46 105
use AOI22X1  AOI22X1_103
timestamp 1682952543
transform 1 0 1584 0 -1 2970
box -8 -3 46 105
use INVX2  INVX2_205
timestamp 1682952543
transform 1 0 1624 0 -1 2970
box -9 -3 26 105
use M3_M2  M3_M2_3046
timestamp 1682952543
transform 1 0 1700 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_203
timestamp 1682952543
transform -1 0 1736 0 -1 2970
box -8 -3 104 105
use M3_M2  M3_M2_3047
timestamp 1682952543
transform 1 0 1748 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_204
timestamp 1682952543
transform -1 0 1832 0 -1 2970
box -8 -3 104 105
use AOI22X1  AOI22X1_110
timestamp 1682952543
transform 1 0 1832 0 -1 2970
box -8 -3 46 105
use INVX2  INVX2_220
timestamp 1682952543
transform 1 0 1872 0 -1 2970
box -9 -3 26 105
use M3_M2  M3_M2_3048
timestamp 1682952543
transform 1 0 1956 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_205
timestamp 1682952543
transform 1 0 1888 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_206
timestamp 1682952543
transform 1 0 1984 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_207
timestamp 1682952543
transform -1 0 2176 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_208
timestamp 1682952543
transform 1 0 2176 0 -1 2970
box -8 -3 104 105
use NAND2X1  NAND2X1_36
timestamp 1682952543
transform 1 0 2272 0 -1 2970
box -8 -3 32 105
use OAI22X1  OAI22X1_182
timestamp 1682952543
transform 1 0 2296 0 -1 2970
box -8 -3 46 105
use OAI21X1  OAI21X1_41
timestamp 1682952543
transform 1 0 2336 0 -1 2970
box -8 -3 34 105
use OAI21X1  OAI21X1_42
timestamp 1682952543
transform -1 0 2400 0 -1 2970
box -8 -3 34 105
use AOI22X1  AOI22X1_111
timestamp 1682952543
transform 1 0 2400 0 -1 2970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_209
timestamp 1682952543
transform -1 0 2536 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_210
timestamp 1682952543
transform 1 0 2536 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_211
timestamp 1682952543
transform -1 0 2728 0 -1 2970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_212
timestamp 1682952543
transform -1 0 2824 0 -1 2970
box -8 -3 104 105
use NOR2X1  NOR2X1_33
timestamp 1682952543
transform 1 0 2824 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_37
timestamp 1682952543
transform 1 0 2848 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_38
timestamp 1682952543
transform 1 0 2872 0 -1 2970
box -8 -3 32 105
use NAND2X1  NAND2X1_39
timestamp 1682952543
transform 1 0 2896 0 -1 2970
box -8 -3 32 105
use NAND3X1  NAND3X1_3
timestamp 1682952543
transform 1 0 2920 0 -1 2970
box -8 -3 40 105
use XOR2X1  XOR2X1_1
timestamp 1682952543
transform 1 0 2952 0 -1 2970
box -8 -3 64 105
use NAND2X1  NAND2X1_40
timestamp 1682952543
transform 1 0 3008 0 -1 2970
box -8 -3 32 105
use NAND3X1  NAND3X1_4
timestamp 1682952543
transform -1 0 3064 0 -1 2970
box -8 -3 40 105
use M3_M2  M3_M2_3049
timestamp 1682952543
transform 1 0 3084 0 1 2875
box -3 -3 3 3
use INVX2  INVX2_221
timestamp 1682952543
transform -1 0 3080 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_222
timestamp 1682952543
transform 1 0 3080 0 -1 2970
box -9 -3 26 105
use AOI21X1  AOI21X1_0
timestamp 1682952543
transform -1 0 3128 0 -1 2970
box -7 -3 39 105
use INVX2  INVX2_223
timestamp 1682952543
transform 1 0 3128 0 -1 2970
box -9 -3 26 105
use INVX2  INVX2_224
timestamp 1682952543
transform 1 0 3144 0 -1 2970
box -9 -3 26 105
use OAI21X1  OAI21X1_43
timestamp 1682952543
transform 1 0 3160 0 -1 2970
box -8 -3 34 105
use M3_M2  M3_M2_3050
timestamp 1682952543
transform 1 0 3204 0 1 2875
box -3 -3 3 3
use FILL  FILL_847
timestamp 1682952543
transform 1 0 3192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_848
timestamp 1682952543
transform 1 0 3200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_849
timestamp 1682952543
transform 1 0 3208 0 -1 2970
box -8 -3 16 105
use AOI21X1  AOI21X1_1
timestamp 1682952543
transform 1 0 3216 0 -1 2970
box -7 -3 39 105
use FILL  FILL_851
timestamp 1682952543
transform 1 0 3248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_853
timestamp 1682952543
transform 1 0 3256 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_44
timestamp 1682952543
transform 1 0 3264 0 -1 2970
box -8 -3 34 105
use NAND2X1  NAND2X1_41
timestamp 1682952543
transform -1 0 3320 0 -1 2970
box -8 -3 32 105
use FILL  FILL_857
timestamp 1682952543
transform 1 0 3320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_859
timestamp 1682952543
transform 1 0 3328 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_114
timestamp 1682952543
transform 1 0 3336 0 -1 2970
box -8 -3 46 105
use FILL  FILL_861
timestamp 1682952543
transform 1 0 3376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_863
timestamp 1682952543
transform 1 0 3384 0 -1 2970
box -8 -3 16 105
use AOI21X1  AOI21X1_2
timestamp 1682952543
transform 1 0 3392 0 -1 2970
box -7 -3 39 105
use NAND3X1  NAND3X1_5
timestamp 1682952543
transform -1 0 3456 0 -1 2970
box -8 -3 40 105
use INVX2  INVX2_226
timestamp 1682952543
transform 1 0 3456 0 -1 2970
box -9 -3 26 105
use NAND3X1  NAND3X1_6
timestamp 1682952543
transform -1 0 3504 0 -1 2970
box -8 -3 40 105
use FILL  FILL_873
timestamp 1682952543
transform 1 0 3504 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_227
timestamp 1682952543
transform 1 0 3512 0 -1 2970
box -9 -3 26 105
use AOI21X1  AOI21X1_3
timestamp 1682952543
transform 1 0 3528 0 -1 2970
box -7 -3 39 105
use AOI22X1  AOI22X1_116
timestamp 1682952543
transform -1 0 3600 0 -1 2970
box -8 -3 46 105
use AND2X1  AND2X1_0
timestamp 1682952543
transform 1 0 3600 0 -1 2970
box -8 -3 40 105
use AOI21X1  AOI21X1_4
timestamp 1682952543
transform 1 0 3632 0 -1 2970
box -7 -3 39 105
use INVX2  INVX2_228
timestamp 1682952543
transform 1 0 3664 0 -1 2970
box -9 -3 26 105
use OAI22X1  OAI22X1_183
timestamp 1682952543
transform -1 0 3720 0 -1 2970
box -8 -3 46 105
use NAND2X1  NAND2X1_42
timestamp 1682952543
transform 1 0 3720 0 -1 2970
box -8 -3 32 105
use AOI21X1  AOI21X1_5
timestamp 1682952543
transform -1 0 3776 0 -1 2970
box -7 -3 39 105
use NAND2X1  NAND2X1_43
timestamp 1682952543
transform 1 0 3776 0 -1 2970
box -8 -3 32 105
use AOI21X1  AOI21X1_6
timestamp 1682952543
transform 1 0 3800 0 -1 2970
box -7 -3 39 105
use INVX2  INVX2_229
timestamp 1682952543
transform -1 0 3848 0 -1 2970
box -9 -3 26 105
use FILL  FILL_874
timestamp 1682952543
transform 1 0 3848 0 -1 2970
box -8 -3 16 105
use AOI21X1  AOI21X1_7
timestamp 1682952543
transform -1 0 3888 0 -1 2970
box -7 -3 39 105
use FILL  FILL_875
timestamp 1682952543
transform 1 0 3888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_876
timestamp 1682952543
transform 1 0 3896 0 -1 2970
box -8 -3 16 105
use AOI21X1  AOI21X1_8
timestamp 1682952543
transform 1 0 3904 0 -1 2970
box -7 -3 39 105
use FILL  FILL_878
timestamp 1682952543
transform 1 0 3936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_879
timestamp 1682952543
transform 1 0 3944 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_230
timestamp 1682952543
transform 1 0 3952 0 -1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_117
timestamp 1682952543
transform 1 0 3968 0 -1 2970
box -8 -3 46 105
use FILL  FILL_880
timestamp 1682952543
transform 1 0 4008 0 -1 2970
box -8 -3 16 105
use FILL  FILL_881
timestamp 1682952543
transform 1 0 4016 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_118
timestamp 1682952543
transform 1 0 4024 0 -1 2970
box -8 -3 46 105
use FILL  FILL_882
timestamp 1682952543
transform 1 0 4064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_883
timestamp 1682952543
transform 1 0 4072 0 -1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1682952543
transform 1 0 4080 0 -1 2970
box -8 -3 40 105
use FILL  FILL_884
timestamp 1682952543
transform 1 0 4112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_885
timestamp 1682952543
transform 1 0 4120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_886
timestamp 1682952543
transform 1 0 4128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_887
timestamp 1682952543
transform 1 0 4136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_888
timestamp 1682952543
transform 1 0 4144 0 -1 2970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_25
timestamp 1682952543
transform 1 0 4201 0 1 2870
box -10 -3 10 3
use M3_M2  M3_M2_3051
timestamp 1682952543
transform 1 0 188 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1682952543
transform 1 0 132 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1682952543
transform 1 0 172 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3067
timestamp 1682952543
transform 1 0 220 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1682952543
transform 1 0 316 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3068
timestamp 1682952543
transform 1 0 332 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1682952543
transform 1 0 316 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1682952543
transform 1 0 284 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1682952543
transform 1 0 324 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3161
timestamp 1682952543
transform 1 0 132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1682952543
transform 1 0 164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3163
timestamp 1682952543
transform 1 0 172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1682952543
transform 1 0 188 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3165
timestamp 1682952543
transform 1 0 204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1682952543
transform 1 0 220 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3167
timestamp 1682952543
transform 1 0 284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1682952543
transform 1 0 316 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3169
timestamp 1682952543
transform 1 0 324 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1682952543
transform 1 0 84 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3230
timestamp 1682952543
transform 1 0 172 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3304
timestamp 1682952543
transform 1 0 180 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1682952543
transform 1 0 196 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3247
timestamp 1682952543
transform 1 0 164 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1682952543
transform 1 0 84 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1682952543
transform 1 0 204 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3306
timestamp 1682952543
transform 1 0 212 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3307
timestamp 1682952543
transform 1 0 220 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3308
timestamp 1682952543
transform 1 0 236 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3248
timestamp 1682952543
transform 1 0 212 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3232
timestamp 1682952543
transform 1 0 324 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1682952543
transform 1 0 236 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1682952543
transform 1 0 260 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1682952543
transform 1 0 348 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3104
timestamp 1682952543
transform 1 0 428 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1682952543
transform 1 0 356 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1682952543
transform 1 0 372 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1682952543
transform 1 0 492 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1682952543
transform 1 0 556 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1682952543
transform 1 0 612 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1682952543
transform 1 0 588 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3105
timestamp 1682952543
transform 1 0 516 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1682952543
transform 1 0 548 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1682952543
transform 1 0 572 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3055
timestamp 1682952543
transform 1 0 644 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1682952543
transform 1 0 628 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3108
timestamp 1682952543
transform 1 0 652 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3151
timestamp 1682952543
transform 1 0 612 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1682952543
transform 1 0 628 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3170
timestamp 1682952543
transform 1 0 332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1682952543
transform 1 0 356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3172
timestamp 1682952543
transform 1 0 372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1682952543
transform 1 0 412 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3174
timestamp 1682952543
transform 1 0 468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3175
timestamp 1682952543
transform 1 0 484 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1682952543
transform 1 0 500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3177
timestamp 1682952543
transform 1 0 508 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1682952543
transform 1 0 572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1682952543
transform 1 0 604 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1682952543
transform 1 0 612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3181
timestamp 1682952543
transform 1 0 628 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1682952543
transform 1 0 644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3183
timestamp 1682952543
transform 1 0 652 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1682952543
transform 1 0 340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3310
timestamp 1682952543
transform 1 0 348 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3311
timestamp 1682952543
transform 1 0 364 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3312
timestamp 1682952543
transform 1 0 372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1682952543
transform 1 0 388 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3294
timestamp 1682952543
transform 1 0 364 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1682952543
transform 1 0 452 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3314
timestamp 1682952543
transform 1 0 476 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3315
timestamp 1682952543
transform 1 0 492 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3249
timestamp 1682952543
transform 1 0 476 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3316
timestamp 1682952543
transform 1 0 524 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3317
timestamp 1682952543
transform 1 0 612 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3318
timestamp 1682952543
transform 1 0 636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3319
timestamp 1682952543
transform 1 0 644 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3250
timestamp 1682952543
transform 1 0 508 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3251
timestamp 1682952543
transform 1 0 588 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1682952543
transform 1 0 604 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3253
timestamp 1682952543
transform 1 0 636 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3295
timestamp 1682952543
transform 1 0 540 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3296
timestamp 1682952543
transform 1 0 564 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3297
timestamp 1682952543
transform 1 0 612 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3153
timestamp 1682952543
transform 1 0 660 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3184
timestamp 1682952543
transform 1 0 660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1682952543
transform 1 0 676 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1682952543
transform 1 0 692 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3320
timestamp 1682952543
transform 1 0 668 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3234
timestamp 1682952543
transform 1 0 676 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3321
timestamp 1682952543
transform 1 0 684 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3254
timestamp 1682952543
transform 1 0 668 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3298
timestamp 1682952543
transform 1 0 684 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3071
timestamp 1682952543
transform 1 0 764 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1682952543
transform 1 0 732 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1682952543
transform 1 0 756 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1682952543
transform 1 0 764 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3187
timestamp 1682952543
transform 1 0 732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1682952543
transform 1 0 748 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3197
timestamp 1682952543
transform 1 0 756 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3189
timestamp 1682952543
transform 1 0 764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3322
timestamp 1682952543
transform 1 0 740 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1682952543
transform 1 0 756 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3324
timestamp 1682952543
transform 1 0 764 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3198
timestamp 1682952543
transform 1 0 788 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3325
timestamp 1682952543
transform 1 0 788 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3056
timestamp 1682952543
transform 1 0 804 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3190
timestamp 1682952543
transform 1 0 796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3191
timestamp 1682952543
transform 1 0 804 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3235
timestamp 1682952543
transform 1 0 812 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1682952543
transform 1 0 852 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1682952543
transform 1 0 852 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1682952543
transform 1 0 836 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1682952543
transform 1 0 868 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3192
timestamp 1682952543
transform 1 0 836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1682952543
transform 1 0 852 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3236
timestamp 1682952543
transform 1 0 836 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1682952543
transform 1 0 860 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3326
timestamp 1682952543
transform 1 0 860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1682952543
transform 1 0 868 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3255
timestamp 1682952543
transform 1 0 860 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3328
timestamp 1682952543
transform 1 0 900 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1682952543
transform 1 0 916 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3299
timestamp 1682952543
transform 1 0 916 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3057
timestamp 1682952543
transform 1 0 940 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3329
timestamp 1682952543
transform 1 0 932 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3112
timestamp 1682952543
transform 1 0 948 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3256
timestamp 1682952543
transform 1 0 940 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1682952543
transform 1 0 964 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3194
timestamp 1682952543
transform 1 0 964 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1682952543
transform 1 0 972 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3113
timestamp 1682952543
transform 1 0 1020 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1682952543
transform 1 0 1036 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1682952543
transform 1 0 1028 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3200
timestamp 1682952543
transform 1 0 1012 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3196
timestamp 1682952543
transform 1 0 1020 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3330
timestamp 1682952543
transform 1 0 1004 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3197
timestamp 1682952543
transform 1 0 1036 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3073
timestamp 1682952543
transform 1 0 1060 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1682952543
transform 1 0 1076 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1682952543
transform 1 0 1092 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3198
timestamp 1682952543
transform 1 0 1076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1682952543
transform 1 0 1092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3331
timestamp 1682952543
transform 1 0 1060 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1682952543
transform 1 0 1068 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3333
timestamp 1682952543
transform 1 0 1084 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3334
timestamp 1682952543
transform 1 0 1092 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3300
timestamp 1682952543
transform 1 0 1076 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1682952543
transform 1 0 1108 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1682952543
transform 1 0 1124 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3200
timestamp 1682952543
transform 1 0 1108 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1682952543
transform 1 0 1124 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3201
timestamp 1682952543
transform 1 0 1132 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3059
timestamp 1682952543
transform 1 0 1164 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3074
timestamp 1682952543
transform 1 0 1164 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1682952543
transform 1 0 1156 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3140
timestamp 1682952543
transform 1 0 1148 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3202
timestamp 1682952543
transform 1 0 1140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1682952543
transform 1 0 1108 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1682952543
transform 1 0 1116 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1682952543
transform 1 0 1140 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3257
timestamp 1682952543
transform 1 0 1140 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3203
timestamp 1682952543
transform 1 0 1156 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3161
timestamp 1682952543
transform 1 0 1172 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3338
timestamp 1682952543
transform 1 0 1172 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3087
timestamp 1682952543
transform 1 0 1268 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1682952543
transform 1 0 1196 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1682952543
transform 1 0 1212 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3117
timestamp 1682952543
transform 1 0 1252 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3162
timestamp 1682952543
transform 1 0 1196 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3163
timestamp 1682952543
transform 1 0 1236 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3164
timestamp 1682952543
transform 1 0 1284 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3204
timestamp 1682952543
transform 1 0 1196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1682952543
transform 1 0 1204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1682952543
transform 1 0 1236 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3202
timestamp 1682952543
transform 1 0 1284 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3339
timestamp 1682952543
transform 1 0 1284 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3258
timestamp 1682952543
transform 1 0 1204 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3259
timestamp 1682952543
transform 1 0 1244 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1682952543
transform 1 0 1268 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3060
timestamp 1682952543
transform 1 0 1300 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1682952543
transform 1 0 1300 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3340
timestamp 1682952543
transform 1 0 1300 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3061
timestamp 1682952543
transform 1 0 1340 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3207
timestamp 1682952543
transform 1 0 1316 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3204
timestamp 1682952543
transform 1 0 1324 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3208
timestamp 1682952543
transform 1 0 1332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3209
timestamp 1682952543
transform 1 0 1348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1682952543
transform 1 0 1324 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3342
timestamp 1682952543
transform 1 0 1340 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3261
timestamp 1682952543
transform 1 0 1324 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3088
timestamp 1682952543
transform 1 0 1420 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3205
timestamp 1682952543
transform 1 0 1396 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3210
timestamp 1682952543
transform 1 0 1428 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3343
timestamp 1682952543
transform 1 0 1460 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3089
timestamp 1682952543
transform 1 0 1492 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3211
timestamp 1682952543
transform 1 0 1492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1682952543
transform 1 0 1500 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3262
timestamp 1682952543
transform 1 0 1500 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3301
timestamp 1682952543
transform 1 0 1500 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1682952543
transform 1 0 1596 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3075
timestamp 1682952543
transform 1 0 1564 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3090
timestamp 1682952543
transform 1 0 1548 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3213
timestamp 1682952543
transform 1 0 1516 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3206
timestamp 1682952543
transform 1 0 1524 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3118
timestamp 1682952543
transform 1 0 1580 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1682952543
transform 1 0 1660 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3091
timestamp 1682952543
transform 1 0 1628 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3119
timestamp 1682952543
transform 1 0 1636 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3120
timestamp 1682952543
transform 1 0 1668 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1682952543
transform 1 0 1564 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3166
timestamp 1682952543
transform 1 0 1588 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1682952543
transform 1 0 1612 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3214
timestamp 1682952543
transform 1 0 1532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1682952543
transform 1 0 1548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3216
timestamp 1682952543
transform 1 0 1556 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1682952543
transform 1 0 1564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1682952543
transform 1 0 1580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1682952543
transform 1 0 1596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3344
timestamp 1682952543
transform 1 0 1516 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3345
timestamp 1682952543
transform 1 0 1524 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3346
timestamp 1682952543
transform 1 0 1540 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3207
timestamp 1682952543
transform 1 0 1604 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3220
timestamp 1682952543
transform 1 0 1612 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1682952543
transform 1 0 1628 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1682952543
transform 1 0 1644 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3237
timestamp 1682952543
transform 1 0 1564 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3347
timestamp 1682952543
transform 1 0 1572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1682952543
transform 1 0 1588 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3238
timestamp 1682952543
transform 1 0 1596 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3349
timestamp 1682952543
transform 1 0 1604 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1682952543
transform 1 0 1620 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3263
timestamp 1682952543
transform 1 0 1588 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1682952543
transform 1 0 1620 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1682952543
transform 1 0 1652 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3223
timestamp 1682952543
transform 1 0 1660 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1682952543
transform 1 0 1668 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3351
timestamp 1682952543
transform 1 0 1652 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3265
timestamp 1682952543
transform 1 0 1644 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3352
timestamp 1682952543
transform 1 0 1676 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3302
timestamp 1682952543
transform 1 0 1668 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3077
timestamp 1682952543
transform 1 0 1732 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1682952543
transform 1 0 1740 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1682952543
transform 1 0 1780 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3225
timestamp 1682952543
transform 1 0 1740 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3209
timestamp 1682952543
transform 1 0 1764 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3226
timestamp 1682952543
transform 1 0 1780 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1682952543
transform 1 0 1764 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3266
timestamp 1682952543
transform 1 0 1684 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3267
timestamp 1682952543
transform 1 0 1740 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1682952543
transform 1 0 1692 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3304
timestamp 1682952543
transform 1 0 1772 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1682952543
transform 1 0 1796 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3064
timestamp 1682952543
transform 1 0 1836 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1682952543
transform 1 0 1860 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3121
timestamp 1682952543
transform 1 0 1804 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1682952543
transform 1 0 1796 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3227
timestamp 1682952543
transform 1 0 1796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3228
timestamp 1682952543
transform 1 0 1812 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3210
timestamp 1682952543
transform 1 0 1820 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1682952543
transform 1 0 1868 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3066
timestamp 1682952543
transform 1 0 1884 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3229
timestamp 1682952543
transform 1 0 1828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1682952543
transform 1 0 1836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3231
timestamp 1682952543
transform 1 0 1852 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3354
timestamp 1682952543
transform 1 0 1796 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1682952543
transform 1 0 1804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3356
timestamp 1682952543
transform 1 0 1820 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3211
timestamp 1682952543
transform 1 0 1860 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3232
timestamp 1682952543
transform 1 0 1868 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3212
timestamp 1682952543
transform 1 0 1876 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3357
timestamp 1682952543
transform 1 0 1844 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3358
timestamp 1682952543
transform 1 0 1860 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1682952543
transform 1 0 1876 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3268
timestamp 1682952543
transform 1 0 1836 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3305
timestamp 1682952543
transform 1 0 1836 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3233
timestamp 1682952543
transform 1 0 1892 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3234
timestamp 1682952543
transform 1 0 1900 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1682952543
transform 1 0 1924 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3122
timestamp 1682952543
transform 1 0 1940 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3236
timestamp 1682952543
transform 1 0 1940 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3360
timestamp 1682952543
transform 1 0 1932 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3269
timestamp 1682952543
transform 1 0 1932 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1682952543
transform 1 0 2036 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3213
timestamp 1682952543
transform 1 0 1972 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3237
timestamp 1682952543
transform 1 0 2004 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1682952543
transform 1 0 1948 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1682952543
transform 1 0 1972 0 1 2807
box -2 -2 2 2
use M3_M2  M3_M2_3172
timestamp 1682952543
transform 1 0 2060 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3238
timestamp 1682952543
transform 1 0 2060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3239
timestamp 1682952543
transform 1 0 2076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1682952543
transform 1 0 2100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1682952543
transform 1 0 2100 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3173
timestamp 1682952543
transform 1 0 2132 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1682952543
transform 1 0 2220 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3241
timestamp 1682952543
transform 1 0 2132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1682952543
transform 1 0 2140 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1682952543
transform 1 0 2172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3363
timestamp 1682952543
transform 1 0 2124 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3270
timestamp 1682952543
transform 1 0 2124 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3306
timestamp 1682952543
transform 1 0 2108 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1682952543
transform 1 0 2220 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3299
timestamp 1682952543
transform 1 0 2220 0 1 2807
box -2 -2 2 2
use M3_M2  M3_M2_3271
timestamp 1682952543
transform 1 0 2148 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1682952543
transform 1 0 2220 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1682952543
transform 1 0 2204 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1682952543
transform 1 0 2308 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1682952543
transform 1 0 2348 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3141
timestamp 1682952543
transform 1 0 2348 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3244
timestamp 1682952543
transform 1 0 2292 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3245
timestamp 1682952543
transform 1 0 2324 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3246
timestamp 1682952543
transform 1 0 2332 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1682952543
transform 1 0 2340 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3364
timestamp 1682952543
transform 1 0 2244 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3239
timestamp 1682952543
transform 1 0 2292 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3365
timestamp 1682952543
transform 1 0 2332 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3125
timestamp 1682952543
transform 1 0 2388 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3142
timestamp 1682952543
transform 1 0 2388 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1682952543
transform 1 0 2372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1682952543
transform 1 0 2380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3366
timestamp 1682952543
transform 1 0 2348 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3176
timestamp 1682952543
transform 1 0 2404 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1682952543
transform 1 0 2508 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1682952543
transform 1 0 2452 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3215
timestamp 1682952543
transform 1 0 2404 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3250
timestamp 1682952543
transform 1 0 2412 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3216
timestamp 1682952543
transform 1 0 2420 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1682952543
transform 1 0 2572 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3178
timestamp 1682952543
transform 1 0 2548 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3251
timestamp 1682952543
transform 1 0 2436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1682952543
transform 1 0 2444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1682952543
transform 1 0 2508 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3254
timestamp 1682952543
transform 1 0 2548 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1682952543
transform 1 0 2596 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3240
timestamp 1682952543
transform 1 0 2396 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3367
timestamp 1682952543
transform 1 0 2412 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3368
timestamp 1682952543
transform 1 0 2420 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3241
timestamp 1682952543
transform 1 0 2436 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3300
timestamp 1682952543
transform 1 0 2444 0 1 2807
box -2 -2 2 2
use M2_M1  M2_M1_3408
timestamp 1682952543
transform 1 0 2428 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3369
timestamp 1682952543
transform 1 0 2532 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3273
timestamp 1682952543
transform 1 0 2516 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3274
timestamp 1682952543
transform 1 0 2532 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3370
timestamp 1682952543
transform 1 0 2628 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3275
timestamp 1682952543
transform 1 0 2628 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3079
timestamp 1682952543
transform 1 0 2684 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1682952543
transform 1 0 2676 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3128
timestamp 1682952543
transform 1 0 2772 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3256
timestamp 1682952543
transform 1 0 2684 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1682952543
transform 1 0 2732 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1682952543
transform 1 0 2772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1682952543
transform 1 0 2828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3260
timestamp 1682952543
transform 1 0 2844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3371
timestamp 1682952543
transform 1 0 2652 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3276
timestamp 1682952543
transform 1 0 2652 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3372
timestamp 1682952543
transform 1 0 2748 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1682952543
transform 1 0 2836 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1682952543
transform 1 0 2860 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3277
timestamp 1682952543
transform 1 0 2748 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1682952543
transform 1 0 2796 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1682952543
transform 1 0 2836 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1682952543
transform 1 0 2852 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3143
timestamp 1682952543
transform 1 0 2876 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3242
timestamp 1682952543
transform 1 0 2892 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3409
timestamp 1682952543
transform 1 0 2892 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1682952543
transform 1 0 2908 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3375
timestamp 1682952543
transform 1 0 2916 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3281
timestamp 1682952543
transform 1 0 2908 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3410
timestamp 1682952543
transform 1 0 2916 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1682952543
transform 1 0 2940 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3179
timestamp 1682952543
transform 1 0 2956 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3243
timestamp 1682952543
transform 1 0 2948 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3376
timestamp 1682952543
transform 1 0 2956 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3092
timestamp 1682952543
transform 1 0 2972 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3133
timestamp 1682952543
transform 1 0 2980 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1682952543
transform 1 0 2972 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3244
timestamp 1682952543
transform 1 0 2972 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_3134
timestamp 1682952543
transform 1 0 2996 0 1 2835
box -2 -2 2 2
use M3_M2  M3_M2_3180
timestamp 1682952543
transform 1 0 2996 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1682952543
transform 1 0 2988 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1682952543
transform 1 0 3044 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3093
timestamp 1682952543
transform 1 0 3020 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1682952543
transform 1 0 3036 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3129
timestamp 1682952543
transform 1 0 3028 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3135
timestamp 1682952543
transform 1 0 3036 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3144
timestamp 1682952543
transform 1 0 3012 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1682952543
transform 1 0 3020 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3217
timestamp 1682952543
transform 1 0 3020 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1682952543
transform 1 0 3084 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1682952543
transform 1 0 3068 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3136
timestamp 1682952543
transform 1 0 3084 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3146
timestamp 1682952543
transform 1 0 3044 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3147
timestamp 1682952543
transform 1 0 3068 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1682952543
transform 1 0 3028 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3245
timestamp 1682952543
transform 1 0 3012 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3218
timestamp 1682952543
transform 1 0 3052 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3148
timestamp 1682952543
transform 1 0 3092 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1682952543
transform 1 0 3060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3266
timestamp 1682952543
transform 1 0 3076 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3377
timestamp 1682952543
transform 1 0 3052 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3219
timestamp 1682952543
transform 1 0 3084 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3096
timestamp 1682952543
transform 1 0 3124 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3137
timestamp 1682952543
transform 1 0 3124 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3149
timestamp 1682952543
transform 1 0 3116 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1682952543
transform 1 0 3140 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3220
timestamp 1682952543
transform 1 0 3124 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3267
timestamp 1682952543
transform 1 0 3132 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3378
timestamp 1682952543
transform 1 0 3156 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3283
timestamp 1682952543
transform 1 0 3156 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3097
timestamp 1682952543
transform 1 0 3308 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3131
timestamp 1682952543
transform 1 0 3292 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3132
timestamp 1682952543
transform 1 0 3316 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1682952543
transform 1 0 3348 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1682952543
transform 1 0 3228 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3182
timestamp 1682952543
transform 1 0 3244 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3268
timestamp 1682952543
transform 1 0 3180 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1682952543
transform 1 0 3188 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3270
timestamp 1682952543
transform 1 0 3204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3271
timestamp 1682952543
transform 1 0 3228 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3272
timestamp 1682952543
transform 1 0 3236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1682952543
transform 1 0 3244 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1682952543
transform 1 0 3196 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3221
timestamp 1682952543
transform 1 0 3268 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1682952543
transform 1 0 3356 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3184
timestamp 1682952543
transform 1 0 3380 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3274
timestamp 1682952543
transform 1 0 3348 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1682952543
transform 1 0 3228 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3284
timestamp 1682952543
transform 1 0 3228 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3222
timestamp 1682952543
transform 1 0 3356 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3275
timestamp 1682952543
transform 1 0 3364 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3223
timestamp 1682952543
transform 1 0 3372 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3381
timestamp 1682952543
transform 1 0 3340 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3301
timestamp 1682952543
transform 1 0 3348 0 1 2807
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1682952543
transform 1 0 3332 0 1 2795
box -2 -2 2 2
use M2_M1  M2_M1_3382
timestamp 1682952543
transform 1 0 3372 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1682952543
transform 1 0 3380 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3134
timestamp 1682952543
transform 1 0 3388 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1682952543
transform 1 0 3396 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3276
timestamp 1682952543
transform 1 0 3388 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3224
timestamp 1682952543
transform 1 0 3396 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3277
timestamp 1682952543
transform 1 0 3420 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3135
timestamp 1682952543
transform 1 0 3436 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3151
timestamp 1682952543
transform 1 0 3436 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1682952543
transform 1 0 3444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1682952543
transform 1 0 3444 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3081
timestamp 1682952543
transform 1 0 3460 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3098
timestamp 1682952543
transform 1 0 3460 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1682952543
transform 1 0 3468 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3152
timestamp 1682952543
transform 1 0 3460 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3186
timestamp 1682952543
transform 1 0 3476 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3153
timestamp 1682952543
transform 1 0 3484 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3279
timestamp 1682952543
transform 1 0 3468 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3225
timestamp 1682952543
transform 1 0 3484 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1682952543
transform 1 0 3508 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3138
timestamp 1682952543
transform 1 0 3508 0 1 2835
box -2 -2 2 2
use M3_M2  M3_M2_3187
timestamp 1682952543
transform 1 0 3508 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3280
timestamp 1682952543
transform 1 0 3500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1682952543
transform 1 0 3500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3281
timestamp 1682952543
transform 1 0 3540 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3386
timestamp 1682952543
transform 1 0 3532 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3387
timestamp 1682952543
transform 1 0 3540 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3285
timestamp 1682952543
transform 1 0 3540 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1682952543
transform 1 0 3532 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1682952543
transform 1 0 3564 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3154
timestamp 1682952543
transform 1 0 3572 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3226
timestamp 1682952543
transform 1 0 3572 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3302
timestamp 1682952543
transform 1 0 3564 0 1 2807
box -2 -2 2 2
use M3_M2  M3_M2_3286
timestamp 1682952543
transform 1 0 3580 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1682952543
transform 1 0 3604 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1682952543
transform 1 0 3596 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3282
timestamp 1682952543
transform 1 0 3604 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3309
timestamp 1682952543
transform 1 0 3604 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3388
timestamp 1682952543
transform 1 0 3612 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1682952543
transform 1 0 3620 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3246
timestamp 1682952543
transform 1 0 3628 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1682952543
transform 1 0 3668 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1682952543
transform 1 0 3700 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3155
timestamp 1682952543
transform 1 0 3668 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3190
timestamp 1682952543
transform 1 0 3676 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3283
timestamp 1682952543
transform 1 0 3644 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1682952543
transform 1 0 3652 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3390
timestamp 1682952543
transform 1 0 3636 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3285
timestamp 1682952543
transform 1 0 3700 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1682952543
transform 1 0 3668 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1682952543
transform 1 0 3676 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1682952543
transform 1 0 3684 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1682952543
transform 1 0 3676 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3310
timestamp 1682952543
transform 1 0 3668 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3413
timestamp 1682952543
transform 1 0 3708 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3311
timestamp 1682952543
transform 1 0 3708 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3100
timestamp 1682952543
transform 1 0 3740 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3286
timestamp 1682952543
transform 1 0 3724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1682952543
transform 1 0 3740 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1682952543
transform 1 0 3756 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1682952543
transform 1 0 3764 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1682952543
transform 1 0 3764 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3396
timestamp 1682952543
transform 1 0 3780 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3287
timestamp 1682952543
transform 1 0 3756 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3414
timestamp 1682952543
transform 1 0 3764 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3288
timestamp 1682952543
transform 1 0 3780 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1682952543
transform 1 0 3764 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3289
timestamp 1682952543
transform 1 0 3796 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3191
timestamp 1682952543
transform 1 0 3812 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1682952543
transform 1 0 3844 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3290
timestamp 1682952543
transform 1 0 3836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1682952543
transform 1 0 3804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1682952543
transform 1 0 3812 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1682952543
transform 1 0 3828 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1682952543
transform 1 0 3852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1682952543
transform 1 0 3884 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1682952543
transform 1 0 3876 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3082
timestamp 1682952543
transform 1 0 3940 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1682952543
transform 1 0 3932 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3193
timestamp 1682952543
transform 1 0 3924 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3140
timestamp 1682952543
transform 1 0 3972 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3156
timestamp 1682952543
transform 1 0 3940 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3292
timestamp 1682952543
transform 1 0 3924 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1682952543
transform 1 0 3908 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3194
timestamp 1682952543
transform 1 0 3956 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3157
timestamp 1682952543
transform 1 0 3972 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3293
timestamp 1682952543
transform 1 0 3956 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3228
timestamp 1682952543
transform 1 0 3964 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3402
timestamp 1682952543
transform 1 0 3940 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3403
timestamp 1682952543
transform 1 0 3948 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3141
timestamp 1682952543
transform 1 0 3988 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3139
timestamp 1682952543
transform 1 0 3996 0 1 2835
box -2 -2 2 2
use M3_M2  M3_M2_3142
timestamp 1682952543
transform 1 0 4012 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3158
timestamp 1682952543
transform 1 0 3980 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3195
timestamp 1682952543
transform 1 0 4004 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3159
timestamp 1682952543
transform 1 0 4012 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1682952543
transform 1 0 4004 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1682952543
transform 1 0 3980 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3229
timestamp 1682952543
transform 1 0 4012 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3295
timestamp 1682952543
transform 1 0 4020 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3083
timestamp 1682952543
transform 1 0 4028 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1682952543
transform 1 0 4068 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1682952543
transform 1 0 4060 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3160
timestamp 1682952543
transform 1 0 4068 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_3296
timestamp 1682952543
transform 1 0 4060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1682952543
transform 1 0 4044 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1682952543
transform 1 0 4052 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3289
timestamp 1682952543
transform 1 0 4044 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3196
timestamp 1682952543
transform 1 0 4076 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3297
timestamp 1682952543
transform 1 0 4076 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3144
timestamp 1682952543
transform 1 0 4092 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3416
timestamp 1682952543
transform 1 0 4132 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3290
timestamp 1682952543
transform 1 0 4220 0 1 2795
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_26
timestamp 1682952543
transform 1 0 48 0 1 2770
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_213
timestamp 1682952543
transform 1 0 72 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_231
timestamp 1682952543
transform -1 0 184 0 1 2770
box -9 -3 26 105
use M3_M2  M3_M2_3313
timestamp 1682952543
transform 1 0 228 0 1 2775
box -3 -3 3 3
use AOI22X1  AOI22X1_119
timestamp 1682952543
transform 1 0 184 0 1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3314
timestamp 1682952543
transform 1 0 276 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3315
timestamp 1682952543
transform 1 0 292 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_215
timestamp 1682952543
transform 1 0 224 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_233
timestamp 1682952543
transform -1 0 336 0 1 2770
box -9 -3 26 105
use AOI22X1  AOI22X1_121
timestamp 1682952543
transform -1 0 376 0 1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3316
timestamp 1682952543
transform 1 0 420 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1682952543
transform 1 0 436 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_216
timestamp 1682952543
transform 1 0 376 0 1 2770
box -8 -3 104 105
use M3_M2  M3_M2_3318
timestamp 1682952543
transform 1 0 484 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1682952543
transform 1 0 516 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_184
timestamp 1682952543
transform -1 0 512 0 1 2770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_217
timestamp 1682952543
transform 1 0 512 0 1 2770
box -8 -3 104 105
use AOI22X1  AOI22X1_122
timestamp 1682952543
transform 1 0 608 0 1 2770
box -8 -3 46 105
use INVX2  INVX2_234
timestamp 1682952543
transform -1 0 664 0 1 2770
box -9 -3 26 105
use M3_M2  M3_M2_3320
timestamp 1682952543
transform 1 0 676 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3321
timestamp 1682952543
transform 1 0 692 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_185
timestamp 1682952543
transform 1 0 664 0 1 2770
box -8 -3 46 105
use FILL  FILL_889
timestamp 1682952543
transform 1 0 704 0 1 2770
box -8 -3 16 105
use FILL  FILL_890
timestamp 1682952543
transform 1 0 712 0 1 2770
box -8 -3 16 105
use FILL  FILL_891
timestamp 1682952543
transform 1 0 720 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3322
timestamp 1682952543
transform 1 0 748 0 1 2775
box -3 -3 3 3
use AOI22X1  AOI22X1_123
timestamp 1682952543
transform -1 0 768 0 1 2770
box -8 -3 46 105
use INVX2  INVX2_235
timestamp 1682952543
transform 1 0 768 0 1 2770
box -9 -3 26 105
use FILL  FILL_892
timestamp 1682952543
transform 1 0 784 0 1 2770
box -8 -3 16 105
use FILL  FILL_893
timestamp 1682952543
transform 1 0 792 0 1 2770
box -8 -3 16 105
use FILL  FILL_894
timestamp 1682952543
transform 1 0 800 0 1 2770
box -8 -3 16 105
use FILL  FILL_901
timestamp 1682952543
transform 1 0 808 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_129
timestamp 1682952543
transform 1 0 816 0 1 2770
box -8 -3 46 105
use FILL  FILL_903
timestamp 1682952543
transform 1 0 856 0 1 2770
box -8 -3 16 105
use FILL  FILL_904
timestamp 1682952543
transform 1 0 864 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_240
timestamp 1682952543
transform 1 0 872 0 1 2770
box -9 -3 26 105
use FILL  FILL_905
timestamp 1682952543
transform 1 0 888 0 1 2770
box -8 -3 16 105
use FILL  FILL_906
timestamp 1682952543
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_907
timestamp 1682952543
transform 1 0 904 0 1 2770
box -8 -3 16 105
use FILL  FILL_908
timestamp 1682952543
transform 1 0 912 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_35
timestamp 1682952543
transform 1 0 920 0 1 2770
box -8 -3 32 105
use FILL  FILL_909
timestamp 1682952543
transform 1 0 944 0 1 2770
box -8 -3 16 105
use FILL  FILL_912
timestamp 1682952543
transform 1 0 952 0 1 2770
box -8 -3 16 105
use FILL  FILL_914
timestamp 1682952543
transform 1 0 960 0 1 2770
box -8 -3 16 105
use FILL  FILL_916
timestamp 1682952543
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_918
timestamp 1682952543
transform 1 0 976 0 1 2770
box -8 -3 16 105
use BUFX2  BUFX2_18
timestamp 1682952543
transform 1 0 984 0 1 2770
box -5 -3 28 105
use FILL  FILL_919
timestamp 1682952543
transform 1 0 1008 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_241
timestamp 1682952543
transform -1 0 1032 0 1 2770
box -9 -3 26 105
use FILL  FILL_920
timestamp 1682952543
transform 1 0 1032 0 1 2770
box -8 -3 16 105
use FILL  FILL_921
timestamp 1682952543
transform 1 0 1040 0 1 2770
box -8 -3 16 105
use FILL  FILL_922
timestamp 1682952543
transform 1 0 1048 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3323
timestamp 1682952543
transform 1 0 1076 0 1 2775
box -3 -3 3 3
use AOI22X1  AOI22X1_130
timestamp 1682952543
transform 1 0 1056 0 1 2770
box -8 -3 46 105
use FILL  FILL_923
timestamp 1682952543
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_131
timestamp 1682952543
transform 1 0 1104 0 1 2770
box -8 -3 46 105
use FILL  FILL_924
timestamp 1682952543
transform 1 0 1144 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_242
timestamp 1682952543
transform 1 0 1152 0 1 2770
box -9 -3 26 105
use FILL  FILL_925
timestamp 1682952543
transform 1 0 1168 0 1 2770
box -8 -3 16 105
use FILL  FILL_926
timestamp 1682952543
transform 1 0 1176 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_243
timestamp 1682952543
transform 1 0 1184 0 1 2770
box -9 -3 26 105
use M3_M2  M3_M2_3324
timestamp 1682952543
transform 1 0 1300 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_221
timestamp 1682952543
transform -1 0 1296 0 1 2770
box -8 -3 104 105
use FILL  FILL_937
timestamp 1682952543
transform 1 0 1296 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3325
timestamp 1682952543
transform 1 0 1316 0 1 2775
box -3 -3 3 3
use FILL  FILL_938
timestamp 1682952543
transform 1 0 1304 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_133
timestamp 1682952543
transform 1 0 1312 0 1 2770
box -8 -3 46 105
use FILL  FILL_939
timestamp 1682952543
transform 1 0 1352 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3326
timestamp 1682952543
transform 1 0 1372 0 1 2775
box -3 -3 3 3
use FILL  FILL_940
timestamp 1682952543
transform 1 0 1360 0 1 2770
box -8 -3 16 105
use FILL  FILL_941
timestamp 1682952543
transform 1 0 1368 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_222
timestamp 1682952543
transform -1 0 1472 0 1 2770
box -8 -3 104 105
use FILL  FILL_942
timestamp 1682952543
transform 1 0 1472 0 1 2770
box -8 -3 16 105
use FILL  FILL_943
timestamp 1682952543
transform 1 0 1480 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_244
timestamp 1682952543
transform -1 0 1504 0 1 2770
box -9 -3 26 105
use FILL  FILL_944
timestamp 1682952543
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_134
timestamp 1682952543
transform 1 0 1512 0 1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3327
timestamp 1682952543
transform 1 0 1572 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_188
timestamp 1682952543
transform 1 0 1552 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_135
timestamp 1682952543
transform 1 0 1592 0 1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_189
timestamp 1682952543
transform -1 0 1672 0 1 2770
box -8 -3 46 105
use FILL  FILL_945
timestamp 1682952543
transform 1 0 1672 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_223
timestamp 1682952543
transform -1 0 1776 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_245
timestamp 1682952543
transform -1 0 1792 0 1 2770
box -9 -3 26 105
use AOI22X1  AOI22X1_136
timestamp 1682952543
transform -1 0 1832 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_137
timestamp 1682952543
transform 1 0 1832 0 1 2770
box -8 -3 46 105
use INVX2  INVX2_246
timestamp 1682952543
transform 1 0 1872 0 1 2770
box -9 -3 26 105
use FILL  FILL_946
timestamp 1682952543
transform 1 0 1888 0 1 2770
box -8 -3 16 105
use FILL  FILL_947
timestamp 1682952543
transform 1 0 1896 0 1 2770
box -8 -3 16 105
use AND2X2  AND2X2_11
timestamp 1682952543
transform -1 0 1936 0 1 2770
box -8 -3 40 105
use FILL  FILL_948
timestamp 1682952543
transform 1 0 1936 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_247
timestamp 1682952543
transform 1 0 1944 0 1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_224
timestamp 1682952543
transform 1 0 1960 0 1 2770
box -8 -3 104 105
use FILL  FILL_949
timestamp 1682952543
transform 1 0 2056 0 1 2770
box -8 -3 16 105
use AND2X2  AND2X2_16
timestamp 1682952543
transform 1 0 2064 0 1 2770
box -8 -3 40 105
use INVX2  INVX2_251
timestamp 1682952543
transform 1 0 2096 0 1 2770
box -9 -3 26 105
use NOR2X1  NOR2X1_38
timestamp 1682952543
transform 1 0 2112 0 1 2770
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_228
timestamp 1682952543
transform -1 0 2232 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_229
timestamp 1682952543
transform 1 0 2232 0 1 2770
box -8 -3 104 105
use M3_M2  M3_M2_3328
timestamp 1682952543
transform 1 0 2356 0 1 2775
box -3 -3 3 3
use NAND2X1  NAND2X1_44
timestamp 1682952543
transform 1 0 2328 0 1 2770
box -8 -3 32 105
use INVX2  INVX2_252
timestamp 1682952543
transform 1 0 2352 0 1 2770
box -9 -3 26 105
use NAND2X1  NAND2X1_45
timestamp 1682952543
transform 1 0 2368 0 1 2770
box -8 -3 32 105
use INVX2  INVX2_253
timestamp 1682952543
transform -1 0 2408 0 1 2770
box -9 -3 26 105
use NOR2X1  NOR2X1_39
timestamp 1682952543
transform -1 0 2432 0 1 2770
box -8 -3 32 105
use INVX2  INVX2_254
timestamp 1682952543
transform -1 0 2448 0 1 2770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_230
timestamp 1682952543
transform -1 0 2544 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_231
timestamp 1682952543
transform -1 0 2640 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_232
timestamp 1682952543
transform 1 0 2640 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_233
timestamp 1682952543
transform 1 0 2736 0 1 2770
box -8 -3 104 105
use OAI21X1  OAI21X1_45
timestamp 1682952543
transform 1 0 2832 0 1 2770
box -8 -3 34 105
use FILL  FILL_988
timestamp 1682952543
transform 1 0 2864 0 1 2770
box -8 -3 16 105
use FILL  FILL_989
timestamp 1682952543
transform 1 0 2872 0 1 2770
box -8 -3 16 105
use FILL  FILL_990
timestamp 1682952543
transform 1 0 2880 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_43
timestamp 1682952543
transform 1 0 2888 0 1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_44
timestamp 1682952543
transform 1 0 2912 0 1 2770
box -8 -3 32 105
use FILL  FILL_991
timestamp 1682952543
transform 1 0 2936 0 1 2770
box -8 -3 16 105
use FILL  FILL_992
timestamp 1682952543
transform 1 0 2944 0 1 2770
box -8 -3 16 105
use FILL  FILL_993
timestamp 1682952543
transform 1 0 2952 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_12
timestamp 1682952543
transform 1 0 2960 0 1 2770
box -8 -3 40 105
use FILL  FILL_994
timestamp 1682952543
transform 1 0 2992 0 1 2770
box -8 -3 16 105
use FILL  FILL_997
timestamp 1682952543
transform 1 0 3000 0 1 2770
box -8 -3 16 105
use FILL  FILL_999
timestamp 1682952543
transform 1 0 3008 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_13
timestamp 1682952543
transform 1 0 3016 0 1 2770
box -8 -3 40 105
use INVX2  INVX2_261
timestamp 1682952543
transform 1 0 3048 0 1 2770
box -9 -3 26 105
use NAND3X1  NAND3X1_14
timestamp 1682952543
transform 1 0 3064 0 1 2770
box -8 -3 40 105
use FILL  FILL_1001
timestamp 1682952543
transform 1 0 3096 0 1 2770
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1682952543
transform 1 0 3104 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_16
timestamp 1682952543
transform -1 0 3144 0 1 2770
box -8 -3 40 105
use FILL  FILL_1008
timestamp 1682952543
transform 1 0 3144 0 1 2770
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1682952543
transform 1 0 3152 0 1 2770
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1682952543
transform 1 0 3160 0 1 2770
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1682952543
transform 1 0 3168 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_263
timestamp 1682952543
transform 1 0 3176 0 1 2770
box -9 -3 26 105
use AND2X2  AND2X2_17
timestamp 1682952543
transform 1 0 3192 0 1 2770
box -8 -3 40 105
use M3_M2  M3_M2_3329
timestamp 1682952543
transform 1 0 3372 0 1 2775
box -3 -3 3 3
use FAX1  FAX1_7
timestamp 1682952543
transform 1 0 3224 0 1 2770
box -5 -3 126 105
use INVX2  INVX2_264
timestamp 1682952543
transform 1 0 3344 0 1 2770
box -9 -3 26 105
use INVX2  INVX2_265
timestamp 1682952543
transform -1 0 3376 0 1 2770
box -9 -3 26 105
use FILL  FILL_1017
timestamp 1682952543
transform 1 0 3376 0 1 2770
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1682952543
transform 1 0 3384 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_47
timestamp 1682952543
transform 1 0 3392 0 1 2770
box -8 -3 34 105
use FILL  FILL_1019
timestamp 1682952543
transform 1 0 3424 0 1 2770
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1682952543
transform 1 0 3432 0 1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_46
timestamp 1682952543
transform 1 0 3440 0 1 2770
box -8 -3 32 105
use FILL  FILL_1021
timestamp 1682952543
transform 1 0 3464 0 1 2770
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1682952543
transform 1 0 3472 0 1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_49
timestamp 1682952543
transform -1 0 3504 0 1 2770
box -8 -3 32 105
use FILL  FILL_1032
timestamp 1682952543
transform 1 0 3504 0 1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_50
timestamp 1682952543
transform -1 0 3536 0 1 2770
box -8 -3 32 105
use OAI21X1  OAI21X1_48
timestamp 1682952543
transform 1 0 3536 0 1 2770
box -8 -3 34 105
use NAND2X1  NAND2X1_51
timestamp 1682952543
transform -1 0 3592 0 1 2770
box -8 -3 32 105
use FILL  FILL_1033
timestamp 1682952543
transform 1 0 3592 0 1 2770
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1682952543
transform 1 0 3600 0 1 2770
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1682952543
transform 1 0 3608 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_266
timestamp 1682952543
transform 1 0 3616 0 1 2770
box -9 -3 26 105
use FILL  FILL_1036
timestamp 1682952543
transform 1 0 3632 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3330
timestamp 1682952543
transform 1 0 3676 0 1 2775
box -3 -3 3 3
use OAI21X1  OAI21X1_49
timestamp 1682952543
transform 1 0 3640 0 1 2770
box -8 -3 34 105
use OR2X1  OR2X1_0
timestamp 1682952543
transform 1 0 3672 0 1 2770
box -8 -3 40 105
use FILL  FILL_1043
timestamp 1682952543
transform 1 0 3704 0 1 2770
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1682952543
transform 1 0 3712 0 1 2770
box -8 -3 16 105
use AOI21X1  AOI21X1_9
timestamp 1682952543
transform -1 0 3752 0 1 2770
box -7 -3 39 105
use FILL  FILL_1045
timestamp 1682952543
transform 1 0 3752 0 1 2770
box -8 -3 16 105
use AOI21X1  AOI21X1_10
timestamp 1682952543
transform -1 0 3792 0 1 2770
box -7 -3 39 105
use FILL  FILL_1046
timestamp 1682952543
transform 1 0 3792 0 1 2770
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1682952543
transform 1 0 3800 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_191
timestamp 1682952543
transform 1 0 3808 0 1 2770
box -8 -3 46 105
use FILL  FILL_1048
timestamp 1682952543
transform 1 0 3848 0 1 2770
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1682952543
transform 1 0 3856 0 1 2770
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1682952543
transform 1 0 3864 0 1 2770
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1682952543
transform 1 0 3872 0 1 2770
box -8 -3 16 105
use AOI21X1  AOI21X1_11
timestamp 1682952543
transform 1 0 3880 0 1 2770
box -7 -3 39 105
use OAI21X1  OAI21X1_50
timestamp 1682952543
transform 1 0 3912 0 1 2770
box -8 -3 34 105
use OAI21X1  OAI21X1_51
timestamp 1682952543
transform 1 0 3944 0 1 2770
box -8 -3 34 105
use FILL  FILL_1054
timestamp 1682952543
transform 1 0 3976 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3331
timestamp 1682952543
transform 1 0 4012 0 1 2775
box -3 -3 3 3
use NAND3X1  NAND3X1_18
timestamp 1682952543
transform -1 0 4016 0 1 2770
box -8 -3 40 105
use FILL  FILL_1055
timestamp 1682952543
transform 1 0 4016 0 1 2770
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1682952543
transform 1 0 4024 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_268
timestamp 1682952543
transform -1 0 4048 0 1 2770
box -9 -3 26 105
use NAND2X1  NAND2X1_52
timestamp 1682952543
transform 1 0 4048 0 1 2770
box -8 -3 32 105
use FILL  FILL_1063
timestamp 1682952543
transform 1 0 4072 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3332
timestamp 1682952543
transform 1 0 4100 0 1 2775
box -3 -3 3 3
use NAND2X1  NAND2X1_53
timestamp 1682952543
transform -1 0 4104 0 1 2770
box -8 -3 32 105
use FILL  FILL_1064
timestamp 1682952543
transform 1 0 4104 0 1 2770
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1682952543
transform 1 0 4112 0 1 2770
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1682952543
transform 1 0 4120 0 1 2770
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1682952543
transform 1 0 4128 0 1 2770
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1682952543
transform 1 0 4136 0 1 2770
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1682952543
transform 1 0 4144 0 1 2770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_27
timestamp 1682952543
transform 1 0 4177 0 1 2770
box -10 -3 10 3
use M2_M1  M2_M1_3434
timestamp 1682952543
transform 1 0 84 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3415
timestamp 1682952543
transform 1 0 164 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1682952543
transform 1 0 196 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3435
timestamp 1682952543
transform 1 0 196 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3416
timestamp 1682952543
transform 1 0 204 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3436
timestamp 1682952543
transform 1 0 212 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1682952543
transform 1 0 220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1682952543
transform 1 0 132 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1682952543
transform 1 0 164 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1682952543
transform 1 0 172 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3525
timestamp 1682952543
transform 1 0 180 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3526
timestamp 1682952543
transform 1 0 188 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3527
timestamp 1682952543
transform 1 0 204 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3460
timestamp 1682952543
transform 1 0 180 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3543
timestamp 1682952543
transform 1 0 188 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1682952543
transform 1 0 156 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1682952543
transform 1 0 268 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1682952543
transform 1 0 260 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3387
timestamp 1682952543
transform 1 0 244 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1682952543
transform 1 0 372 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1682952543
transform 1 0 332 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3438
timestamp 1682952543
transform 1 0 244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1682952543
transform 1 0 260 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1682952543
transform 1 0 276 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3417
timestamp 1682952543
transform 1 0 284 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3441
timestamp 1682952543
transform 1 0 300 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3418
timestamp 1682952543
transform 1 0 308 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1682952543
transform 1 0 404 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1682952543
transform 1 0 420 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1682952543
transform 1 0 444 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1682952543
transform 1 0 388 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3442
timestamp 1682952543
transform 1 0 316 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3443
timestamp 1682952543
transform 1 0 332 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3444
timestamp 1682952543
transform 1 0 340 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1682952543
transform 1 0 356 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3446
timestamp 1682952543
transform 1 0 364 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1682952543
transform 1 0 252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1682952543
transform 1 0 276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3530
timestamp 1682952543
transform 1 0 284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1682952543
transform 1 0 292 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3439
timestamp 1682952543
transform 1 0 300 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3532
timestamp 1682952543
transform 1 0 308 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3533
timestamp 1682952543
transform 1 0 324 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1682952543
transform 1 0 332 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3461
timestamp 1682952543
transform 1 0 252 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1682952543
transform 1 0 276 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1682952543
transform 1 0 292 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3503
timestamp 1682952543
transform 1 0 268 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1682952543
transform 1 0 244 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1682952543
transform 1 0 340 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3535
timestamp 1682952543
transform 1 0 348 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3441
timestamp 1682952543
transform 1 0 356 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3419
timestamp 1682952543
transform 1 0 380 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3447
timestamp 1682952543
transform 1 0 388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3448
timestamp 1682952543
transform 1 0 404 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3420
timestamp 1682952543
transform 1 0 412 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3389
timestamp 1682952543
transform 1 0 476 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1682952543
transform 1 0 524 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3449
timestamp 1682952543
transform 1 0 420 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3450
timestamp 1682952543
transform 1 0 428 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1682952543
transform 1 0 444 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1682952543
transform 1 0 460 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1682952543
transform 1 0 476 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3536
timestamp 1682952543
transform 1 0 364 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3464
timestamp 1682952543
transform 1 0 324 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3537
timestamp 1682952543
transform 1 0 380 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1682952543
transform 1 0 396 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3539
timestamp 1682952543
transform 1 0 420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3540
timestamp 1682952543
transform 1 0 436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1682952543
transform 1 0 452 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3465
timestamp 1682952543
transform 1 0 364 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1682952543
transform 1 0 380 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1682952543
transform 1 0 396 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3504
timestamp 1682952543
transform 1 0 332 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3544
timestamp 1682952543
transform 1 0 356 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3442
timestamp 1682952543
transform 1 0 460 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3542
timestamp 1682952543
transform 1 0 524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1682952543
transform 1 0 556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1682952543
transform 1 0 564 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3545
timestamp 1682952543
transform 1 0 572 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3468
timestamp 1682952543
transform 1 0 436 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1682952543
transform 1 0 420 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3506
timestamp 1682952543
transform 1 0 452 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1682952543
transform 1 0 524 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1682952543
transform 1 0 564 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3507
timestamp 1682952543
transform 1 0 556 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3563
timestamp 1682952543
transform 1 0 556 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_3454
timestamp 1682952543
transform 1 0 596 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3455
timestamp 1682952543
transform 1 0 604 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1682952543
transform 1 0 620 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3391
timestamp 1682952543
transform 1 0 644 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1682952543
transform 1 0 724 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3457
timestamp 1682952543
transform 1 0 644 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1682952543
transform 1 0 612 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3547
timestamp 1682952543
transform 1 0 628 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3548
timestamp 1682952543
transform 1 0 692 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3508
timestamp 1682952543
transform 1 0 620 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1682952543
transform 1 0 596 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3546
timestamp 1682952543
transform 1 0 612 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3443
timestamp 1682952543
transform 1 0 708 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3549
timestamp 1682952543
transform 1 0 724 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1682952543
transform 1 0 732 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1682952543
transform 1 0 740 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3471
timestamp 1682952543
transform 1 0 692 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1682952543
transform 1 0 732 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1682952543
transform 1 0 724 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3336
timestamp 1682952543
transform 1 0 804 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_3420
timestamp 1682952543
transform 1 0 804 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3458
timestamp 1682952543
transform 1 0 764 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3459
timestamp 1682952543
transform 1 0 772 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1682952543
transform 1 0 788 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3421
timestamp 1682952543
transform 1 0 796 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3552
timestamp 1682952543
transform 1 0 780 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3553
timestamp 1682952543
transform 1 0 796 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3473
timestamp 1682952543
transform 1 0 796 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3510
timestamp 1682952543
transform 1 0 772 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3547
timestamp 1682952543
transform 1 0 788 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3564
timestamp 1682952543
transform 1 0 796 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1682952543
transform 1 0 828 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3461
timestamp 1682952543
transform 1 0 820 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3565
timestamp 1682952543
transform 1 0 812 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_3462
timestamp 1682952543
transform 1 0 836 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3394
timestamp 1682952543
transform 1 0 860 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3463
timestamp 1682952543
transform 1 0 860 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3444
timestamp 1682952543
transform 1 0 860 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3337
timestamp 1682952543
transform 1 0 948 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1682952543
transform 1 0 948 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3421
timestamp 1682952543
transform 1 0 948 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3554
timestamp 1682952543
transform 1 0 900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1682952543
transform 1 0 940 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3395
timestamp 1682952543
transform 1 0 964 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3548
timestamp 1682952543
transform 1 0 956 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3396
timestamp 1682952543
transform 1 0 980 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3417
timestamp 1682952543
transform 1 0 1004 0 1 2755
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1682952543
transform 1 0 1012 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3418
timestamp 1682952543
transform 1 0 1028 0 1 2755
box -2 -2 2 2
use M3_M2  M3_M2_3397
timestamp 1682952543
transform 1 0 1028 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3422
timestamp 1682952543
transform 1 0 1036 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3556
timestamp 1682952543
transform 1 0 1028 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1682952543
transform 1 0 1036 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1682952543
transform 1 0 1052 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3474
timestamp 1682952543
transform 1 0 1052 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3511
timestamp 1682952543
transform 1 0 1036 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3465
timestamp 1682952543
transform 1 0 1068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1682952543
transform 1 0 1076 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3445
timestamp 1682952543
transform 1 0 1076 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3559
timestamp 1682952543
transform 1 0 1084 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3512
timestamp 1682952543
transform 1 0 1068 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3475
timestamp 1682952543
transform 1 0 1084 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3467
timestamp 1682952543
transform 1 0 1108 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3338
timestamp 1682952543
transform 1 0 1140 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1682952543
transform 1 0 1132 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3423
timestamp 1682952543
transform 1 0 1140 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1682952543
transform 1 0 1172 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3468
timestamp 1682952543
transform 1 0 1164 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3469
timestamp 1682952543
transform 1 0 1172 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3560
timestamp 1682952543
transform 1 0 1140 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1682952543
transform 1 0 1156 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1682952543
transform 1 0 1204 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3446
timestamp 1682952543
transform 1 0 1196 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1682952543
transform 1 0 1252 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3471
timestamp 1682952543
transform 1 0 1244 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3562
timestamp 1682952543
transform 1 0 1236 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3563
timestamp 1682952543
transform 1 0 1252 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3363
timestamp 1682952543
transform 1 0 1276 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3447
timestamp 1682952543
transform 1 0 1284 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1682952543
transform 1 0 1292 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3472
timestamp 1682952543
transform 1 0 1292 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3473
timestamp 1682952543
transform 1 0 1300 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3448
timestamp 1682952543
transform 1 0 1300 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1682952543
transform 1 0 1316 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_3474
timestamp 1682952543
transform 1 0 1316 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3340
timestamp 1682952543
transform 1 0 1332 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1682952543
transform 1 0 1340 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3424
timestamp 1682952543
transform 1 0 1332 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3475
timestamp 1682952543
transform 1 0 1356 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3425
timestamp 1682952543
transform 1 0 1364 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3564
timestamp 1682952543
transform 1 0 1324 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3565
timestamp 1682952543
transform 1 0 1332 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3449
timestamp 1682952543
transform 1 0 1340 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3566
timestamp 1682952543
transform 1 0 1348 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3513
timestamp 1682952543
transform 1 0 1332 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3514
timestamp 1682952543
transform 1 0 1348 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1682952543
transform 1 0 1380 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3567
timestamp 1682952543
transform 1 0 1372 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3341
timestamp 1682952543
transform 1 0 1412 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3426
timestamp 1682952543
transform 1 0 1396 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3476
timestamp 1682952543
transform 1 0 1404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1682952543
transform 1 0 1412 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1682952543
transform 1 0 1396 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3476
timestamp 1682952543
transform 1 0 1396 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3515
timestamp 1682952543
transform 1 0 1388 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3342
timestamp 1682952543
transform 1 0 1436 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_3569
timestamp 1682952543
transform 1 0 1428 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1682952543
transform 1 0 1436 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3549
timestamp 1682952543
transform 1 0 1436 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1682952543
transform 1 0 1460 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3368
timestamp 1682952543
transform 1 0 1556 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3478
timestamp 1682952543
transform 1 0 1452 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1682952543
transform 1 0 1468 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3369
timestamp 1682952543
transform 1 0 1604 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1682952543
transform 1 0 1628 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3371
timestamp 1682952543
transform 1 0 1684 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1682952543
transform 1 0 1652 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3399
timestamp 1682952543
transform 1 0 1668 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3480
timestamp 1682952543
transform 1 0 1580 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3481
timestamp 1682952543
transform 1 0 1668 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1682952543
transform 1 0 1684 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1682952543
transform 1 0 1492 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3572
timestamp 1682952543
transform 1 0 1548 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3573
timestamp 1682952543
transform 1 0 1556 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1682952543
transform 1 0 1572 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3516
timestamp 1682952543
transform 1 0 1468 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1682952543
transform 1 0 1492 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3566
timestamp 1682952543
transform 1 0 1452 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3567
timestamp 1682952543
transform 1 0 1484 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1682952543
transform 1 0 1508 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3450
timestamp 1682952543
transform 1 0 1580 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3575
timestamp 1682952543
transform 1 0 1588 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3576
timestamp 1682952543
transform 1 0 1636 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3577
timestamp 1682952543
transform 1 0 1684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1682952543
transform 1 0 1700 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3477
timestamp 1682952543
transform 1 0 1636 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3478
timestamp 1682952543
transform 1 0 1684 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3479
timestamp 1682952543
transform 1 0 1700 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3518
timestamp 1682952543
transform 1 0 1668 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3569
timestamp 1682952543
transform 1 0 1588 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3400
timestamp 1682952543
transform 1 0 1724 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3483
timestamp 1682952543
transform 1 0 1724 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1682952543
transform 1 0 1748 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1682952543
transform 1 0 1756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1682952543
transform 1 0 1732 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3480
timestamp 1682952543
transform 1 0 1732 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3451
timestamp 1682952543
transform 1 0 1756 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3634
timestamp 1682952543
transform 1 0 1756 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3550
timestamp 1682952543
transform 1 0 1764 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3343
timestamp 1682952543
transform 1 0 1796 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3372
timestamp 1682952543
transform 1 0 1828 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3344
timestamp 1682952543
transform 1 0 1932 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1682952543
transform 1 0 1924 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3486
timestamp 1682952543
transform 1 0 1836 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3427
timestamp 1682952543
transform 1 0 1900 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3487
timestamp 1682952543
transform 1 0 1924 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3401
timestamp 1682952543
transform 1 0 1948 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3580
timestamp 1682952543
transform 1 0 1788 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1682952543
transform 1 0 1804 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3582
timestamp 1682952543
transform 1 0 1812 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3583
timestamp 1682952543
transform 1 0 1828 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1682952543
transform 1 0 1844 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3585
timestamp 1682952543
transform 1 0 1892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1682952543
transform 1 0 1780 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3481
timestamp 1682952543
transform 1 0 1812 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1682952543
transform 1 0 1788 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1682952543
transform 1 0 1940 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3586
timestamp 1682952543
transform 1 0 1956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3636
timestamp 1682952543
transform 1 0 1940 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3519
timestamp 1682952543
transform 1 0 1884 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3520
timestamp 1682952543
transform 1 0 1940 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3637
timestamp 1682952543
transform 1 0 1964 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3638
timestamp 1682952543
transform 1 0 1972 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1682952543
transform 1 0 1948 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3551
timestamp 1682952543
transform 1 0 1924 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1682952543
transform 1 0 1964 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3402
timestamp 1682952543
transform 1 0 1988 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3453
timestamp 1682952543
transform 1 0 1996 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3587
timestamp 1682952543
transform 1 0 2012 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1682952543
transform 1 0 1996 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3482
timestamp 1682952543
transform 1 0 2004 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3640
timestamp 1682952543
transform 1 0 2020 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1682952543
transform 1 0 2004 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3345
timestamp 1682952543
transform 1 0 2076 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1682952543
transform 1 0 2068 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3375
timestamp 1682952543
transform 1 0 2084 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3422
timestamp 1682952543
transform 1 0 2076 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1682952543
transform 1 0 2068 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3483
timestamp 1682952543
transform 1 0 2068 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3571
timestamp 1682952543
transform 1 0 2068 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_3588
timestamp 1682952543
transform 1 0 2092 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3346
timestamp 1682952543
transform 1 0 2108 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1682952543
transform 1 0 2100 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1682952543
transform 1 0 2140 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1682952543
transform 1 0 2172 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3404
timestamp 1682952543
transform 1 0 2196 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3489
timestamp 1682952543
transform 1 0 2196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1682952543
transform 1 0 2156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3348
timestamp 1682952543
transform 1 0 2252 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3405
timestamp 1682952543
transform 1 0 2228 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3490
timestamp 1682952543
transform 1 0 2228 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3590
timestamp 1682952543
transform 1 0 2252 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3522
timestamp 1682952543
transform 1 0 2252 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3552
timestamp 1682952543
transform 1 0 2276 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_3423
timestamp 1682952543
transform 1 0 2324 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1682952543
transform 1 0 2316 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3591
timestamp 1682952543
transform 1 0 2324 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3553
timestamp 1682952543
transform 1 0 2316 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3406
timestamp 1682952543
transform 1 0 2340 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3492
timestamp 1682952543
transform 1 0 2340 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3592
timestamp 1682952543
transform 1 0 2348 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3485
timestamp 1682952543
transform 1 0 2332 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1682952543
transform 1 0 2348 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3554
timestamp 1682952543
transform 1 0 2340 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_3493
timestamp 1682952543
transform 1 0 2372 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3486
timestamp 1682952543
transform 1 0 2372 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3494
timestamp 1682952543
transform 1 0 2396 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3524
timestamp 1682952543
transform 1 0 2388 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3376
timestamp 1682952543
transform 1 0 2476 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3495
timestamp 1682952543
transform 1 0 2516 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1682952543
transform 1 0 2420 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1682952543
transform 1 0 2436 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1682952543
transform 1 0 2476 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3596
timestamp 1682952543
transform 1 0 2532 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1682952543
transform 1 0 2540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1682952543
transform 1 0 2548 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3487
timestamp 1682952543
transform 1 0 2420 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3641
timestamp 1682952543
transform 1 0 2428 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3653
timestamp 1682952543
transform 1 0 2412 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3525
timestamp 1682952543
transform 1 0 2428 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1682952543
transform 1 0 2532 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1682952543
transform 1 0 2548 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3407
timestamp 1682952543
transform 1 0 2636 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3496
timestamp 1682952543
transform 1 0 2636 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1682952543
transform 1 0 2612 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3489
timestamp 1682952543
transform 1 0 2612 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1682952543
transform 1 0 2756 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3377
timestamp 1682952543
transform 1 0 2692 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3378
timestamp 1682952543
transform 1 0 2748 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1682952543
transform 1 0 2668 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3497
timestamp 1682952543
transform 1 0 2668 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3428
timestamp 1682952543
transform 1 0 2692 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3498
timestamp 1682952543
transform 1 0 2756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3600
timestamp 1682952543
transform 1 0 2692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1682952543
transform 1 0 2756 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3499
timestamp 1682952543
transform 1 0 2772 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3490
timestamp 1682952543
transform 1 0 2772 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3424
timestamp 1682952543
transform 1 0 2804 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3429
timestamp 1682952543
transform 1 0 2804 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3602
timestamp 1682952543
transform 1 0 2804 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3555
timestamp 1682952543
transform 1 0 2804 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1682952543
transform 1 0 2828 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3603
timestamp 1682952543
transform 1 0 2820 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3491
timestamp 1682952543
transform 1 0 2820 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3642
timestamp 1682952543
transform 1 0 2828 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1682952543
transform 1 0 2828 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1682952543
transform 1 0 2844 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3492
timestamp 1682952543
transform 1 0 2844 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3655
timestamp 1682952543
transform 1 0 2852 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3431
timestamp 1682952543
transform 1 0 2868 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3605
timestamp 1682952543
transform 1 0 2868 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1682952543
transform 1 0 2868 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3527
timestamp 1682952543
transform 1 0 2868 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3500
timestamp 1682952543
transform 1 0 2892 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1682952543
transform 1 0 2884 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3493
timestamp 1682952543
transform 1 0 2884 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3425
timestamp 1682952543
transform 1 0 2908 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3501
timestamp 1682952543
transform 1 0 2908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1682952543
transform 1 0 2916 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3454
timestamp 1682952543
transform 1 0 2916 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3503
timestamp 1682952543
transform 1 0 2932 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3607
timestamp 1682952543
transform 1 0 2924 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3528
timestamp 1682952543
transform 1 0 2932 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3608
timestamp 1682952543
transform 1 0 2940 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1682952543
transform 1 0 2964 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3504
timestamp 1682952543
transform 1 0 2972 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3505
timestamp 1682952543
transform 1 0 2980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1682952543
transform 1 0 2988 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3455
timestamp 1682952543
transform 1 0 2964 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3494
timestamp 1682952543
transform 1 0 2972 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1682952543
transform 1 0 2988 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3609
timestamp 1682952543
transform 1 0 3028 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3495
timestamp 1682952543
transform 1 0 3036 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3656
timestamp 1682952543
transform 1 0 3036 0 1 2705
box -2 -2 2 2
use M2_M1  M2_M1_3610
timestamp 1682952543
transform 1 0 3044 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1682952543
transform 1 0 3044 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1682952543
transform 1 0 3060 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3496
timestamp 1682952543
transform 1 0 3084 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3657
timestamp 1682952543
transform 1 0 3084 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3556
timestamp 1682952543
transform 1 0 3100 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3456
timestamp 1682952543
transform 1 0 3116 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3612
timestamp 1682952543
transform 1 0 3132 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3645
timestamp 1682952543
transform 1 0 3116 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1682952543
transform 1 0 3124 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3530
timestamp 1682952543
transform 1 0 3124 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3647
timestamp 1682952543
transform 1 0 3148 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3379
timestamp 1682952543
transform 1 0 3188 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3613
timestamp 1682952543
transform 1 0 3180 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3497
timestamp 1682952543
transform 1 0 3180 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1682952543
transform 1 0 3212 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3381
timestamp 1682952543
transform 1 0 3236 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3507
timestamp 1682952543
transform 1 0 3212 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1682952543
transform 1 0 3204 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1682952543
transform 1 0 3204 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3531
timestamp 1682952543
transform 1 0 3204 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3409
timestamp 1682952543
transform 1 0 3276 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3615
timestamp 1682952543
transform 1 0 3236 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3616
timestamp 1682952543
transform 1 0 3260 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3617
timestamp 1682952543
transform 1 0 3268 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3498
timestamp 1682952543
transform 1 0 3236 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1682952543
transform 1 0 3212 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3558
timestamp 1682952543
transform 1 0 3260 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_3649
timestamp 1682952543
transform 1 0 3276 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3532
timestamp 1682952543
transform 1 0 3276 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1682952543
transform 1 0 3308 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3618
timestamp 1682952543
transform 1 0 3300 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1682952543
transform 1 0 3316 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3350
timestamp 1682952543
transform 1 0 3332 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_3509
timestamp 1682952543
transform 1 0 3332 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3351
timestamp 1682952543
transform 1 0 3348 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_3427
timestamp 1682952543
transform 1 0 3444 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3432
timestamp 1682952543
transform 1 0 3396 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3619
timestamp 1682952543
transform 1 0 3348 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1682952543
transform 1 0 3356 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3457
timestamp 1682952543
transform 1 0 3372 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1682952543
transform 1 0 3348 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3534
timestamp 1682952543
transform 1 0 3412 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3510
timestamp 1682952543
transform 1 0 3460 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3499
timestamp 1682952543
transform 1 0 3460 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3352
timestamp 1682952543
transform 1 0 3492 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_3419
timestamp 1682952543
transform 1 0 3492 0 1 2755
box -2 -2 2 2
use M3_M2  M3_M2_3410
timestamp 1682952543
transform 1 0 3484 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3353
timestamp 1682952543
transform 1 0 3516 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_3428
timestamp 1682952543
transform 1 0 3604 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3411
timestamp 1682952543
transform 1 0 3612 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3621
timestamp 1682952543
transform 1 0 3500 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1682952543
transform 1 0 3508 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1682952543
transform 1 0 3516 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3535
timestamp 1682952543
transform 1 0 3492 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1682952543
transform 1 0 3516 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1682952543
transform 1 0 3524 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1682952543
transform 1 0 3508 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3560
timestamp 1682952543
transform 1 0 3540 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3383
timestamp 1682952543
transform 1 0 3644 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3511
timestamp 1682952543
transform 1 0 3644 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3412
timestamp 1682952543
transform 1 0 3660 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3624
timestamp 1682952543
transform 1 0 3652 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3501
timestamp 1682952543
transform 1 0 3644 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_3429
timestamp 1682952543
transform 1 0 3780 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3384
timestamp 1682952543
transform 1 0 3916 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3430
timestamp 1682952543
transform 1 0 3804 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3413
timestamp 1682952543
transform 1 0 3812 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3414
timestamp 1682952543
transform 1 0 3908 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_3512
timestamp 1682952543
transform 1 0 3668 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1682952543
transform 1 0 3676 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3433
timestamp 1682952543
transform 1 0 3692 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1682952543
transform 1 0 3788 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3514
timestamp 1682952543
transform 1 0 3796 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3435
timestamp 1682952543
transform 1 0 3804 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3436
timestamp 1682952543
transform 1 0 3860 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3431
timestamp 1682952543
transform 1 0 3940 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3515
timestamp 1682952543
transform 1 0 3908 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1682952543
transform 1 0 3916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3517
timestamp 1682952543
transform 1 0 3924 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1682952543
transform 1 0 3940 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3458
timestamp 1682952543
transform 1 0 3668 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_3625
timestamp 1682952543
transform 1 0 3684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3626
timestamp 1682952543
transform 1 0 3692 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3627
timestamp 1682952543
transform 1 0 3892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1682952543
transform 1 0 3900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3629
timestamp 1682952543
transform 1 0 3916 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3537
timestamp 1682952543
transform 1 0 3684 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1682952543
transform 1 0 3732 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3539
timestamp 1682952543
transform 1 0 3788 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3540
timestamp 1682952543
transform 1 0 3900 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3572
timestamp 1682952543
transform 1 0 3772 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3459
timestamp 1682952543
transform 1 0 3924 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3437
timestamp 1682952543
transform 1 0 3948 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3630
timestamp 1682952543
transform 1 0 3948 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1682952543
transform 1 0 3956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1682952543
transform 1 0 3980 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3438
timestamp 1682952543
transform 1 0 3996 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_3519
timestamp 1682952543
transform 1 0 4004 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3385
timestamp 1682952543
transform 1 0 4020 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3632
timestamp 1682952543
transform 1 0 4012 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3386
timestamp 1682952543
transform 1 0 4052 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_3433
timestamp 1682952543
transform 1 0 4132 0 1 2745
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1682952543
transform 1 0 4028 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3650
timestamp 1682952543
transform 1 0 4020 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3541
timestamp 1682952543
transform 1 0 4020 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_3521
timestamp 1682952543
transform 1 0 4140 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_3633
timestamp 1682952543
transform 1 0 4044 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3502
timestamp 1682952543
transform 1 0 4044 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1682952543
transform 1 0 4148 0 1 2705
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_28
timestamp 1682952543
transform 1 0 24 0 1 2670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_214
timestamp 1682952543
transform 1 0 72 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_232
timestamp 1682952543
transform -1 0 184 0 -1 2770
box -9 -3 26 105
use AOI22X1  AOI22X1_120
timestamp 1682952543
transform 1 0 184 0 -1 2770
box -8 -3 46 105
use FILL  FILL_895
timestamp 1682952543
transform 1 0 224 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_124
timestamp 1682952543
transform -1 0 272 0 -1 2770
box -8 -3 46 105
use INVX2  INVX2_236
timestamp 1682952543
transform 1 0 272 0 -1 2770
box -9 -3 26 105
use AOI22X1  AOI22X1_125
timestamp 1682952543
transform 1 0 288 0 -1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_126
timestamp 1682952543
transform 1 0 328 0 -1 2770
box -8 -3 46 105
use INVX2  INVX2_237
timestamp 1682952543
transform 1 0 368 0 -1 2770
box -9 -3 26 105
use OAI22X1  OAI22X1_186
timestamp 1682952543
transform -1 0 424 0 -1 2770
box -8 -3 46 105
use OAI22X1  OAI22X1_187
timestamp 1682952543
transform -1 0 464 0 -1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3573
timestamp 1682952543
transform 1 0 508 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_218
timestamp 1682952543
transform 1 0 464 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_238
timestamp 1682952543
transform -1 0 576 0 -1 2770
box -9 -3 26 105
use FILL  FILL_896
timestamp 1682952543
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_897
timestamp 1682952543
transform 1 0 584 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3574
timestamp 1682952543
transform 1 0 628 0 1 2675
box -3 -3 3 3
use AOI22X1  AOI22X1_127
timestamp 1682952543
transform 1 0 592 0 -1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3575
timestamp 1682952543
transform 1 0 716 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_219
timestamp 1682952543
transform 1 0 632 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_239
timestamp 1682952543
transform -1 0 744 0 -1 2770
box -9 -3 26 105
use FILL  FILL_898
timestamp 1682952543
transform 1 0 744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_899
timestamp 1682952543
transform 1 0 752 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3576
timestamp 1682952543
transform 1 0 772 0 1 2675
box -3 -3 3 3
use AOI22X1  AOI22X1_128
timestamp 1682952543
transform -1 0 800 0 -1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3577
timestamp 1682952543
transform 1 0 812 0 1 2675
box -3 -3 3 3
use FILL  FILL_900
timestamp 1682952543
transform 1 0 800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_902
timestamp 1682952543
transform 1 0 808 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3578
timestamp 1682952543
transform 1 0 828 0 1 2675
box -3 -3 3 3
use NOR2X1  NOR2X1_36
timestamp 1682952543
transform 1 0 816 0 -1 2770
box -8 -3 32 105
use FILL  FILL_910
timestamp 1682952543
transform 1 0 840 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3579
timestamp 1682952543
transform 1 0 876 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3580
timestamp 1682952543
transform 1 0 924 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_220
timestamp 1682952543
transform 1 0 848 0 -1 2770
box -8 -3 104 105
use FILL  FILL_911
timestamp 1682952543
transform 1 0 944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_913
timestamp 1682952543
transform 1 0 952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_915
timestamp 1682952543
transform 1 0 960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_917
timestamp 1682952543
transform 1 0 968 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_37
timestamp 1682952543
transform 1 0 976 0 -1 2770
box -8 -3 32 105
use FILL  FILL_927
timestamp 1682952543
transform 1 0 1000 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3581
timestamp 1682952543
transform 1 0 1020 0 1 2675
box -3 -3 3 3
use FILL  FILL_928
timestamp 1682952543
transform 1 0 1008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_929
timestamp 1682952543
transform 1 0 1016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_930
timestamp 1682952543
transform 1 0 1024 0 -1 2770
box -8 -3 16 105
use AND2X2  AND2X2_9
timestamp 1682952543
transform -1 0 1064 0 -1 2770
box -8 -3 40 105
use FILL  FILL_931
timestamp 1682952543
transform 1 0 1064 0 -1 2770
box -8 -3 16 105
use AND2X2  AND2X2_10
timestamp 1682952543
transform 1 0 1072 0 -1 2770
box -8 -3 40 105
use FILL  FILL_932
timestamp 1682952543
transform 1 0 1104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_933
timestamp 1682952543
transform 1 0 1112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_934
timestamp 1682952543
transform 1 0 1120 0 -1 2770
box -8 -3 16 105
use FILL  FILL_935
timestamp 1682952543
transform 1 0 1128 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_132
timestamp 1682952543
transform 1 0 1136 0 -1 2770
box -8 -3 46 105
use FILL  FILL_936
timestamp 1682952543
transform 1 0 1176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_950
timestamp 1682952543
transform 1 0 1184 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3582
timestamp 1682952543
transform 1 0 1204 0 1 2675
box -3 -3 3 3
use FILL  FILL_951
timestamp 1682952543
transform 1 0 1192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_952
timestamp 1682952543
transform 1 0 1200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_953
timestamp 1682952543
transform 1 0 1208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_954
timestamp 1682952543
transform 1 0 1216 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3583
timestamp 1682952543
transform 1 0 1260 0 1 2675
box -3 -3 3 3
use OAI22X1  OAI22X1_190
timestamp 1682952543
transform -1 0 1264 0 -1 2770
box -8 -3 46 105
use FILL  FILL_955
timestamp 1682952543
transform 1 0 1264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_956
timestamp 1682952543
transform 1 0 1272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_957
timestamp 1682952543
transform 1 0 1280 0 -1 2770
box -8 -3 16 105
use FILL  FILL_958
timestamp 1682952543
transform 1 0 1288 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_248
timestamp 1682952543
transform 1 0 1296 0 -1 2770
box -9 -3 26 105
use FILL  FILL_959
timestamp 1682952543
transform 1 0 1312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_960
timestamp 1682952543
transform 1 0 1320 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_138
timestamp 1682952543
transform -1 0 1368 0 -1 2770
box -8 -3 46 105
use FILL  FILL_961
timestamp 1682952543
transform 1 0 1368 0 -1 2770
box -8 -3 16 105
use AND2X2  AND2X2_12
timestamp 1682952543
transform -1 0 1408 0 -1 2770
box -8 -3 40 105
use INVX2  INVX2_249
timestamp 1682952543
transform 1 0 1408 0 -1 2770
box -9 -3 26 105
use FILL  FILL_962
timestamp 1682952543
transform 1 0 1424 0 -1 2770
box -8 -3 16 105
use BUFX2  BUFX2_19
timestamp 1682952543
transform 1 0 1432 0 -1 2770
box -5 -3 28 105
use M3_M2  M3_M2_3584
timestamp 1682952543
transform 1 0 1508 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_225
timestamp 1682952543
transform 1 0 1456 0 -1 2770
box -8 -3 104 105
use AND2X2  AND2X2_13
timestamp 1682952543
transform -1 0 1584 0 -1 2770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_226
timestamp 1682952543
transform -1 0 1680 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_250
timestamp 1682952543
transform 1 0 1680 0 -1 2770
box -9 -3 26 105
use FILL  FILL_963
timestamp 1682952543
transform 1 0 1696 0 -1 2770
box -8 -3 16 105
use BUFX2  BUFX2_20
timestamp 1682952543
transform 1 0 1704 0 -1 2770
box -5 -3 28 105
use M3_M2  M3_M2_3585
timestamp 1682952543
transform 1 0 1748 0 1 2675
box -3 -3 3 3
use BUFX2  BUFX2_21
timestamp 1682952543
transform 1 0 1728 0 -1 2770
box -5 -3 28 105
use FILL  FILL_964
timestamp 1682952543
transform 1 0 1752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_965
timestamp 1682952543
transform 1 0 1760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_966
timestamp 1682952543
transform 1 0 1768 0 -1 2770
box -8 -3 16 105
use AND2X2  AND2X2_14
timestamp 1682952543
transform 1 0 1776 0 -1 2770
box -8 -3 40 105
use AND2X2  AND2X2_15
timestamp 1682952543
transform -1 0 1840 0 -1 2770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_227
timestamp 1682952543
transform -1 0 1936 0 -1 2770
box -8 -3 104 105
use NAND3X1  NAND3X1_8
timestamp 1682952543
transform -1 0 1968 0 -1 2770
box -8 -3 40 105
use FILL  FILL_967
timestamp 1682952543
transform 1 0 1968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_968
timestamp 1682952543
transform 1 0 1976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_969
timestamp 1682952543
transform 1 0 1984 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3586
timestamp 1682952543
transform 1 0 2020 0 1 2675
box -3 -3 3 3
use NAND3X1  NAND3X1_9
timestamp 1682952543
transform -1 0 2024 0 -1 2770
box -8 -3 40 105
use FILL  FILL_970
timestamp 1682952543
transform 1 0 2024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_971
timestamp 1682952543
transform 1 0 2032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_972
timestamp 1682952543
transform 1 0 2040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_973
timestamp 1682952543
transform 1 0 2048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_974
timestamp 1682952543
transform 1 0 2056 0 -1 2770
box -8 -3 16 105
use FILL  FILL_975
timestamp 1682952543
transform 1 0 2064 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3587
timestamp 1682952543
transform 1 0 2100 0 1 2675
box -3 -3 3 3
use NOR2X1  NOR2X1_40
timestamp 1682952543
transform 1 0 2072 0 -1 2770
box -8 -3 32 105
use FILL  FILL_976
timestamp 1682952543
transform 1 0 2096 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3588
timestamp 1682952543
transform 1 0 2116 0 1 2675
box -3 -3 3 3
use FILL  FILL_977
timestamp 1682952543
transform 1 0 2104 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3589
timestamp 1682952543
transform 1 0 2188 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_234
timestamp 1682952543
transform -1 0 2208 0 -1 2770
box -8 -3 104 105
use FILL  FILL_978
timestamp 1682952543
transform 1 0 2208 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3590
timestamp 1682952543
transform 1 0 2244 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3591
timestamp 1682952543
transform 1 0 2268 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_235
timestamp 1682952543
transform 1 0 2216 0 -1 2770
box -8 -3 104 105
use FILL  FILL_979
timestamp 1682952543
transform 1 0 2312 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_41
timestamp 1682952543
transform 1 0 2320 0 -1 2770
box -8 -3 32 105
use INVX2  INVX2_255
timestamp 1682952543
transform 1 0 2344 0 -1 2770
box -9 -3 26 105
use FILL  FILL_980
timestamp 1682952543
transform 1 0 2360 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3592
timestamp 1682952543
transform 1 0 2388 0 1 2675
box -3 -3 3 3
use OAI21X1  OAI21X1_46
timestamp 1682952543
transform 1 0 2368 0 -1 2770
box -8 -3 34 105
use M3_M2  M3_M2_3593
timestamp 1682952543
transform 1 0 2436 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3594
timestamp 1682952543
transform 1 0 2484 0 1 2675
box -3 -3 3 3
use NAND3X1  NAND3X1_10
timestamp 1682952543
transform -1 0 2432 0 -1 2770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_236
timestamp 1682952543
transform -1 0 2528 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_256
timestamp 1682952543
transform 1 0 2528 0 -1 2770
box -9 -3 26 105
use FILL  FILL_981
timestamp 1682952543
transform 1 0 2544 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_237
timestamp 1682952543
transform -1 0 2648 0 -1 2770
box -8 -3 104 105
use M3_M2  M3_M2_3595
timestamp 1682952543
transform 1 0 2676 0 1 2675
box -3 -3 3 3
use FILL  FILL_982
timestamp 1682952543
transform 1 0 2648 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_238
timestamp 1682952543
transform 1 0 2656 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_257
timestamp 1682952543
transform 1 0 2752 0 -1 2770
box -9 -3 26 105
use FILL  FILL_983
timestamp 1682952543
transform 1 0 2768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_984
timestamp 1682952543
transform 1 0 2776 0 -1 2770
box -8 -3 16 105
use FILL  FILL_985
timestamp 1682952543
transform 1 0 2784 0 -1 2770
box -8 -3 16 105
use FILL  FILL_986
timestamp 1682952543
transform 1 0 2792 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_42
timestamp 1682952543
transform 1 0 2800 0 -1 2770
box -8 -3 32 105
use FILL  FILL_987
timestamp 1682952543
transform 1 0 2824 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_11
timestamp 1682952543
transform 1 0 2832 0 -1 2770
box -8 -3 40 105
use FILL  FILL_995
timestamp 1682952543
transform 1 0 2864 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3596
timestamp 1682952543
transform 1 0 2892 0 1 2675
box -3 -3 3 3
use INVX2  INVX2_258
timestamp 1682952543
transform -1 0 2888 0 -1 2770
box -9 -3 26 105
use NOR2X1  NOR2X1_45
timestamp 1682952543
transform -1 0 2912 0 -1 2770
box -8 -3 32 105
use INVX2  INVX2_259
timestamp 1682952543
transform 1 0 2912 0 -1 2770
box -9 -3 26 105
use M3_M2  M3_M2_3597
timestamp 1682952543
transform 1 0 2948 0 1 2675
box -3 -3 3 3
use INVX2  INVX2_260
timestamp 1682952543
transform 1 0 2928 0 -1 2770
box -9 -3 26 105
use NOR2X1  NOR2X1_46
timestamp 1682952543
transform -1 0 2968 0 -1 2770
box -8 -3 32 105
use NOR2X1  NOR2X1_47
timestamp 1682952543
transform 1 0 2968 0 -1 2770
box -8 -3 32 105
use FILL  FILL_996
timestamp 1682952543
transform 1 0 2992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_998
timestamp 1682952543
transform 1 0 3000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1682952543
transform 1 0 3008 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_262
timestamp 1682952543
transform 1 0 3016 0 -1 2770
box -9 -3 26 105
use FILL  FILL_1002
timestamp 1682952543
transform 1 0 3032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1682952543
transform 1 0 3040 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_15
timestamp 1682952543
transform 1 0 3048 0 -1 2770
box -8 -3 40 105
use FILL  FILL_1004
timestamp 1682952543
transform 1 0 3080 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1682952543
transform 1 0 3088 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1682952543
transform 1 0 3096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1682952543
transform 1 0 3104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1682952543
transform 1 0 3112 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_17
timestamp 1682952543
transform 1 0 3120 0 -1 2770
box -8 -3 40 105
use FILL  FILL_1012
timestamp 1682952543
transform 1 0 3152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1682952543
transform 1 0 3160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1682952543
transform 1 0 3168 0 -1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_47
timestamp 1682952543
transform 1 0 3176 0 -1 2770
box -8 -3 32 105
use FILL  FILL_1022
timestamp 1682952543
transform 1 0 3200 0 -1 2770
box -8 -3 16 105
use XOR2X1  XOR2X1_2
timestamp 1682952543
transform 1 0 3208 0 -1 2770
box -8 -3 64 105
use FILL  FILL_1023
timestamp 1682952543
transform 1 0 3264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1024
timestamp 1682952543
transform 1 0 3272 0 -1 2770
box -8 -3 16 105
use NAND2X1  NAND2X1_48
timestamp 1682952543
transform -1 0 3304 0 -1 2770
box -8 -3 32 105
use FILL  FILL_1025
timestamp 1682952543
transform 1 0 3304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1682952543
transform 1 0 3312 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1682952543
transform 1 0 3320 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1682952543
transform 1 0 3328 0 -1 2770
box -8 -3 16 105
use FAX1  FAX1_8
timestamp 1682952543
transform 1 0 3336 0 -1 2770
box -5 -3 126 105
use FILL  FILL_1029
timestamp 1682952543
transform 1 0 3456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1682952543
transform 1 0 3464 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1682952543
transform 1 0 3472 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1682952543
transform 1 0 3480 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3598
timestamp 1682952543
transform 1 0 3500 0 1 2675
box -3 -3 3 3
use FILL  FILL_1039
timestamp 1682952543
transform 1 0 3488 0 -1 2770
box -8 -3 16 105
use FAX1  FAX1_9
timestamp 1682952543
transform 1 0 3496 0 -1 2770
box -5 -3 126 105
use FILL  FILL_1040
timestamp 1682952543
transform 1 0 3616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1682952543
transform 1 0 3624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1682952543
transform 1 0 3632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1682952543
transform 1 0 3640 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1682952543
transform 1 0 3648 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_267
timestamp 1682952543
transform -1 0 3672 0 -1 2770
box -9 -3 26 105
use M3_M2  M3_M2_3599
timestamp 1682952543
transform 1 0 3724 0 1 2675
box -3 -3 3 3
use FAX1  FAX1_10
timestamp 1682952543
transform 1 0 3672 0 -1 2770
box -5 -3 126 105
use FAX1  FAX1_11
timestamp 1682952543
transform -1 0 3912 0 -1 2770
box -5 -3 126 105
use AOI21X1  AOI21X1_12
timestamp 1682952543
transform 1 0 3912 0 -1 2770
box -7 -3 39 105
use FILL  FILL_1056
timestamp 1682952543
transform 1 0 3944 0 -1 2770
box -8 -3 16 105
use AOI21X1  AOI21X1_13
timestamp 1682952543
transform 1 0 3952 0 -1 2770
box -7 -3 39 105
use FILL  FILL_1057
timestamp 1682952543
transform 1 0 3984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1682952543
transform 1 0 3992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1682952543
transform 1 0 4000 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1682952543
transform 1 0 4008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1682952543
transform 1 0 4016 0 -1 2770
box -8 -3 16 105
use FAX1  FAX1_12
timestamp 1682952543
transform 1 0 4024 0 -1 2770
box -5 -3 126 105
use FILL  FILL_1070
timestamp 1682952543
transform 1 0 4144 0 -1 2770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_29
timestamp 1682952543
transform 1 0 4201 0 1 2670
box -10 -3 10 3
use M3_M2  M3_M2_3667
timestamp 1682952543
transform 1 0 108 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3691
timestamp 1682952543
transform 1 0 116 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3679
timestamp 1682952543
transform 1 0 92 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1682952543
transform 1 0 116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3796
timestamp 1682952543
transform 1 0 76 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1682952543
transform 1 0 100 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3762
timestamp 1682952543
transform 1 0 108 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3786
timestamp 1682952543
transform 1 0 116 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3600
timestamp 1682952543
transform 1 0 212 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1682952543
transform 1 0 156 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1682952543
transform 1 0 204 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3681
timestamp 1682952543
transform 1 0 148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3682
timestamp 1682952543
transform 1 0 156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1682952543
transform 1 0 140 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3763
timestamp 1682952543
transform 1 0 148 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3736
timestamp 1682952543
transform 1 0 172 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3683
timestamp 1682952543
transform 1 0 196 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3737
timestamp 1682952543
transform 1 0 204 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3635
timestamp 1682952543
transform 1 0 356 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1682952543
transform 1 0 372 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1682952543
transform 1 0 316 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3695
timestamp 1682952543
transform 1 0 348 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3684
timestamp 1682952543
transform 1 0 252 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3685
timestamp 1682952543
transform 1 0 292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1682952543
transform 1 0 348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1682952543
transform 1 0 356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1682952543
transform 1 0 372 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3799
timestamp 1682952543
transform 1 0 172 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3764
timestamp 1682952543
transform 1 0 236 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3787
timestamp 1682952543
transform 1 0 172 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1682952543
transform 1 0 380 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3689
timestamp 1682952543
transform 1 0 388 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3800
timestamp 1682952543
transform 1 0 268 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3765
timestamp 1682952543
transform 1 0 348 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_3801
timestamp 1682952543
transform 1 0 356 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3802
timestamp 1682952543
transform 1 0 380 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3803
timestamp 1682952543
transform 1 0 388 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3788
timestamp 1682952543
transform 1 0 268 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3789
timestamp 1682952543
transform 1 0 300 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1682952543
transform 1 0 508 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1682952543
transform 1 0 420 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3696
timestamp 1682952543
transform 1 0 404 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1682952543
transform 1 0 444 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3690
timestamp 1682952543
transform 1 0 404 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1682952543
transform 1 0 444 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3739
timestamp 1682952543
transform 1 0 492 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3602
timestamp 1682952543
transform 1 0 540 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3636
timestamp 1682952543
transform 1 0 556 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1682952543
transform 1 0 548 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3692
timestamp 1682952543
transform 1 0 500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1682952543
transform 1 0 516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1682952543
transform 1 0 532 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3740
timestamp 1682952543
transform 1 0 540 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3695
timestamp 1682952543
transform 1 0 548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3696
timestamp 1682952543
transform 1 0 556 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1682952543
transform 1 0 420 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3805
timestamp 1682952543
transform 1 0 508 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3806
timestamp 1682952543
transform 1 0 524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1682952543
transform 1 0 540 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3790
timestamp 1682952543
transform 1 0 404 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3791
timestamp 1682952543
transform 1 0 420 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1682952543
transform 1 0 524 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1682952543
transform 1 0 532 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3699
timestamp 1682952543
transform 1 0 612 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3664
timestamp 1682952543
transform 1 0 620 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3741
timestamp 1682952543
transform 1 0 580 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3697
timestamp 1682952543
transform 1 0 588 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3742
timestamp 1682952543
transform 1 0 604 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3808
timestamp 1682952543
transform 1 0 572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1682952543
transform 1 0 580 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3810
timestamp 1682952543
transform 1 0 596 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3698
timestamp 1682952543
transform 1 0 620 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3766
timestamp 1682952543
transform 1 0 620 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1682952543
transform 1 0 636 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3700
timestamp 1682952543
transform 1 0 652 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3699
timestamp 1682952543
transform 1 0 652 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3743
timestamp 1682952543
transform 1 0 660 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3637
timestamp 1682952543
transform 1 0 676 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3700
timestamp 1682952543
transform 1 0 668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3811
timestamp 1682952543
transform 1 0 660 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3701
timestamp 1682952543
transform 1 0 716 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3701
timestamp 1682952543
transform 1 0 716 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3824
timestamp 1682952543
transform 1 0 700 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3793
timestamp 1682952543
transform 1 0 724 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_3877
timestamp 1682952543
transform 1 0 732 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3615
timestamp 1682952543
transform 1 0 756 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_3812
timestamp 1682952543
transform 1 0 756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3813
timestamp 1682952543
transform 1 0 764 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3702
timestamp 1682952543
transform 1 0 780 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3814
timestamp 1682952543
transform 1 0 788 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3616
timestamp 1682952543
transform 1 0 836 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3638
timestamp 1682952543
transform 1 0 852 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1682952543
transform 1 0 828 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3702
timestamp 1682952543
transform 1 0 828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3703
timestamp 1682952543
transform 1 0 836 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3744
timestamp 1682952543
transform 1 0 844 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3704
timestamp 1682952543
transform 1 0 852 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3815
timestamp 1682952543
transform 1 0 844 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3767
timestamp 1682952543
transform 1 0 852 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1682952543
transform 1 0 844 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1682952543
transform 1 0 836 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3603
timestamp 1682952543
transform 1 0 868 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3745
timestamp 1682952543
transform 1 0 868 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3768
timestamp 1682952543
transform 1 0 868 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_3878
timestamp 1682952543
transform 1 0 868 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3746
timestamp 1682952543
transform 1 0 900 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3816
timestamp 1682952543
transform 1 0 900 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3639
timestamp 1682952543
transform 1 0 924 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3817
timestamp 1682952543
transform 1 0 916 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3604
timestamp 1682952543
transform 1 0 948 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1682952543
transform 1 0 940 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3705
timestamp 1682952543
transform 1 0 948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3706
timestamp 1682952543
transform 1 0 956 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3769
timestamp 1682952543
transform 1 0 948 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3617
timestamp 1682952543
transform 1 0 972 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3748
timestamp 1682952543
transform 1 0 972 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3707
timestamp 1682952543
transform 1 0 980 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1682952543
transform 1 0 972 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3795
timestamp 1682952543
transform 1 0 972 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1682952543
transform 1 0 988 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3826
timestamp 1682952543
transform 1 0 988 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3640
timestamp 1682952543
transform 1 0 1012 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3641
timestamp 1682952543
transform 1 0 1028 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3665
timestamp 1682952543
transform 1 0 1012 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3771
timestamp 1682952543
transform 1 0 1004 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_3708
timestamp 1682952543
transform 1 0 1020 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1682952543
transform 1 0 1036 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3772
timestamp 1682952543
transform 1 0 1020 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3749
timestamp 1682952543
transform 1 0 1060 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3819
timestamp 1682952543
transform 1 0 1060 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3796
timestamp 1682952543
transform 1 0 1052 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3827
timestamp 1682952543
transform 1 0 1044 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1682952543
transform 1 0 1084 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3619
timestamp 1682952543
transform 1 0 1108 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1682952543
transform 1 0 1140 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1682952543
transform 1 0 1156 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1682952543
transform 1 0 1076 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1682952543
transform 1 0 1164 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3710
timestamp 1682952543
transform 1 0 1124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1682952543
transform 1 0 1164 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3712
timestamp 1682952543
transform 1 0 1172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1682952543
transform 1 0 1076 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3773
timestamp 1682952543
transform 1 0 1108 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3774
timestamp 1682952543
transform 1 0 1124 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_3821
timestamp 1682952543
transform 1 0 1164 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3775
timestamp 1682952543
transform 1 0 1172 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3797
timestamp 1682952543
transform 1 0 1140 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3798
timestamp 1682952543
transform 1 0 1156 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3644
timestamp 1682952543
transform 1 0 1212 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3822
timestamp 1682952543
transform 1 0 1212 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3605
timestamp 1682952543
transform 1 0 1244 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_3713
timestamp 1682952543
transform 1 0 1228 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1682952543
transform 1 0 1244 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1682952543
transform 1 0 1236 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3799
timestamp 1682952543
transform 1 0 1228 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3828
timestamp 1682952543
transform 1 0 1260 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3622
timestamp 1682952543
transform 1 0 1292 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1682952543
transform 1 0 1316 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_3715
timestamp 1682952543
transform 1 0 1292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1682952543
transform 1 0 1324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1682952543
transform 1 0 1388 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3776
timestamp 1682952543
transform 1 0 1340 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_3824
timestamp 1682952543
transform 1 0 1372 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3606
timestamp 1682952543
transform 1 0 1420 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1682952543
transform 1 0 1404 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3645
timestamp 1682952543
transform 1 0 1436 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3718
timestamp 1682952543
transform 1 0 1428 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3646
timestamp 1682952543
transform 1 0 1476 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3647
timestamp 1682952543
transform 1 0 1524 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1682952543
transform 1 0 1516 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3719
timestamp 1682952543
transform 1 0 1452 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1682952543
transform 1 0 1476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1682952543
transform 1 0 1500 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3722
timestamp 1682952543
transform 1 0 1508 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1682952543
transform 1 0 1524 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3825
timestamp 1682952543
transform 1 0 1444 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3826
timestamp 1682952543
transform 1 0 1468 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3800
timestamp 1682952543
transform 1 0 1420 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3801
timestamp 1682952543
transform 1 0 1444 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1682952543
transform 1 0 1404 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1682952543
transform 1 0 1436 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3648
timestamp 1682952543
transform 1 0 1636 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3724
timestamp 1682952543
transform 1 0 1572 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3750
timestamp 1682952543
transform 1 0 1580 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3751
timestamp 1682952543
transform 1 0 1596 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3725
timestamp 1682952543
transform 1 0 1628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3726
timestamp 1682952543
transform 1 0 1636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3827
timestamp 1682952543
transform 1 0 1492 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3828
timestamp 1682952543
transform 1 0 1516 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3829
timestamp 1682952543
transform 1 0 1532 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3830
timestamp 1682952543
transform 1 0 1548 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3802
timestamp 1682952543
transform 1 0 1596 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1682952543
transform 1 0 1548 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1682952543
transform 1 0 1652 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_3831
timestamp 1682952543
transform 1 0 1660 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3803
timestamp 1682952543
transform 1 0 1660 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3649
timestamp 1682952543
transform 1 0 1692 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3607
timestamp 1682952543
transform 1 0 1764 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3672
timestamp 1682952543
transform 1 0 1756 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3727
timestamp 1682952543
transform 1 0 1700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3832
timestamp 1682952543
transform 1 0 1676 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3833
timestamp 1682952543
transform 1 0 1676 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3625
timestamp 1682952543
transform 1 0 1780 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1682952543
transform 1 0 1788 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1682952543
transform 1 0 1780 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3728
timestamp 1682952543
transform 1 0 1772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1682952543
transform 1 0 1780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1682952543
transform 1 0 1796 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3752
timestamp 1682952543
transform 1 0 1804 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3731
timestamp 1682952543
transform 1 0 1812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1682952543
transform 1 0 1828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3833
timestamp 1682952543
transform 1 0 1804 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3650
timestamp 1682952543
transform 1 0 1844 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3666
timestamp 1682952543
transform 1 0 1844 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3834
timestamp 1682952543
transform 1 0 1836 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3834
timestamp 1682952543
transform 1 0 1828 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3626
timestamp 1682952543
transform 1 0 1876 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1682952543
transform 1 0 1860 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3658
timestamp 1682952543
transform 1 0 1860 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_3674
timestamp 1682952543
transform 1 0 1868 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1682952543
transform 1 0 1908 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3667
timestamp 1682952543
transform 1 0 1876 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3668
timestamp 1682952543
transform 1 0 1884 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1682952543
transform 1 0 1868 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3704
timestamp 1682952543
transform 1 0 1900 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3669
timestamp 1682952543
transform 1 0 1908 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1682952543
transform 1 0 1900 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3627
timestamp 1682952543
transform 1 0 1924 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_3659
timestamp 1682952543
transform 1 0 1924 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_3652
timestamp 1682952543
transform 1 0 1948 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1682952543
transform 1 0 1956 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3660
timestamp 1682952543
transform 1 0 1964 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_3670
timestamp 1682952543
transform 1 0 1932 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3705
timestamp 1682952543
transform 1 0 1948 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3671
timestamp 1682952543
transform 1 0 1956 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1682952543
transform 1 0 1948 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3753
timestamp 1682952543
transform 1 0 1956 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3804
timestamp 1682952543
transform 1 0 1956 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3628
timestamp 1682952543
transform 1 0 1996 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3608
timestamp 1682952543
transform 1 0 2036 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3653
timestamp 1682952543
transform 1 0 1988 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1682952543
transform 1 0 2004 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1682952543
transform 1 0 2028 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3661
timestamp 1682952543
transform 1 0 1988 0 1 2635
box -2 -2 2 2
use M3_M2  M3_M2_3677
timestamp 1682952543
transform 1 0 1996 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3672
timestamp 1682952543
transform 1 0 1980 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3805
timestamp 1682952543
transform 1 0 1972 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1682952543
transform 1 0 2020 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3662
timestamp 1682952543
transform 1 0 2028 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_3673
timestamp 1682952543
transform 1 0 2004 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3706
timestamp 1682952543
transform 1 0 2012 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3674
timestamp 1682952543
transform 1 0 2028 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3707
timestamp 1682952543
transform 1 0 2036 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3675
timestamp 1682952543
transform 1 0 2052 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1682952543
transform 1 0 1996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3737
timestamp 1682952543
transform 1 0 2012 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3835
timestamp 1682952543
transform 1 0 2012 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1682952543
transform 1 0 2036 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3806
timestamp 1682952543
transform 1 0 2028 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_3836
timestamp 1682952543
transform 1 0 2060 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3807
timestamp 1682952543
transform 1 0 2052 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3835
timestamp 1682952543
transform 1 0 2060 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1682952543
transform 1 0 2084 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_3879
timestamp 1682952543
transform 1 0 2076 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3629
timestamp 1682952543
transform 1 0 2108 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1682952543
transform 1 0 2100 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1682952543
transform 1 0 2092 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3739
timestamp 1682952543
transform 1 0 2092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3837
timestamp 1682952543
transform 1 0 2092 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3709
timestamp 1682952543
transform 1 0 2116 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3838
timestamp 1682952543
transform 1 0 2108 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1682952543
transform 1 0 2124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1682952543
transform 1 0 2124 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3658
timestamp 1682952543
transform 1 0 2156 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1682952543
transform 1 0 2156 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1682952543
transform 1 0 2164 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3741
timestamp 1682952543
transform 1 0 2140 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1682952543
transform 1 0 2156 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3836
timestamp 1682952543
transform 1 0 2148 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_3840
timestamp 1682952543
transform 1 0 2164 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3630
timestamp 1682952543
transform 1 0 2180 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_3743
timestamp 1682952543
transform 1 0 2180 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3609
timestamp 1682952543
transform 1 0 2204 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3711
timestamp 1682952543
transform 1 0 2212 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3744
timestamp 1682952543
transform 1 0 2220 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1682952543
transform 1 0 2212 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3712
timestamp 1682952543
transform 1 0 2260 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3745
timestamp 1682952543
transform 1 0 2236 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1682952543
transform 1 0 2252 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3837
timestamp 1682952543
transform 1 0 2236 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_3842
timestamp 1682952543
transform 1 0 2260 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3680
timestamp 1682952543
transform 1 0 2276 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3747
timestamp 1682952543
transform 1 0 2276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3748
timestamp 1682952543
transform 1 0 2292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3749
timestamp 1682952543
transform 1 0 2300 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3777
timestamp 1682952543
transform 1 0 2300 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1682952543
transform 1 0 2356 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1682952543
transform 1 0 2380 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1682952543
transform 1 0 2396 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3750
timestamp 1682952543
transform 1 0 2332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3751
timestamp 1682952543
transform 1 0 2348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1682952543
transform 1 0 2356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3753
timestamp 1682952543
transform 1 0 2364 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3754
timestamp 1682952543
transform 1 0 2380 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3843
timestamp 1682952543
transform 1 0 2340 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3778
timestamp 1682952543
transform 1 0 2364 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1682952543
transform 1 0 2340 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_3844
timestamp 1682952543
transform 1 0 2388 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1682952543
transform 1 0 2396 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3839
timestamp 1682952543
transform 1 0 2388 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1682952543
transform 1 0 2492 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1682952543
transform 1 0 2476 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3755
timestamp 1682952543
transform 1 0 2412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1682952543
transform 1 0 2420 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1682952543
transform 1 0 2476 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1682952543
transform 1 0 2412 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1682952543
transform 1 0 2500 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3631
timestamp 1682952543
transform 1 0 2540 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3717
timestamp 1682952543
transform 1 0 2556 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3611
timestamp 1682952543
transform 1 0 2660 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3659
timestamp 1682952543
transform 1 0 2684 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1682952543
transform 1 0 2716 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1682952543
transform 1 0 2724 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3718
timestamp 1682952543
transform 1 0 2620 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3719
timestamp 1682952543
transform 1 0 2668 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1682952543
transform 1 0 2740 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3720
timestamp 1682952543
transform 1 0 2732 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3758
timestamp 1682952543
transform 1 0 2548 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3759
timestamp 1682952543
transform 1 0 2604 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3760
timestamp 1682952543
transform 1 0 2620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3761
timestamp 1682952543
transform 1 0 2628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1682952543
transform 1 0 2668 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1682952543
transform 1 0 2524 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3849
timestamp 1682952543
transform 1 0 2612 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3840
timestamp 1682952543
transform 1 0 2556 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3754
timestamp 1682952543
transform 1 0 2724 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3763
timestamp 1682952543
transform 1 0 2732 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1682952543
transform 1 0 2740 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1682952543
transform 1 0 2708 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1682952543
transform 1 0 2724 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3779
timestamp 1682952543
transform 1 0 2740 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1682952543
transform 1 0 2732 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3612
timestamp 1682952543
transform 1 0 2756 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1682952543
transform 1 0 2756 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1682952543
transform 1 0 2780 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3755
timestamp 1682952543
transform 1 0 2764 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3765
timestamp 1682952543
transform 1 0 2772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3766
timestamp 1682952543
transform 1 0 2780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1682952543
transform 1 0 2756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3853
timestamp 1682952543
transform 1 0 2764 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3808
timestamp 1682952543
transform 1 0 2764 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3842
timestamp 1682952543
transform 1 0 2756 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1682952543
transform 1 0 2796 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3721
timestamp 1682952543
transform 1 0 2796 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3663
timestamp 1682952543
transform 1 0 2836 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1682952543
transform 1 0 2820 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3722
timestamp 1682952543
transform 1 0 2836 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3677
timestamp 1682952543
transform 1 0 2844 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3723
timestamp 1682952543
transform 1 0 2860 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3767
timestamp 1682952543
transform 1 0 2812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1682952543
transform 1 0 2828 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3769
timestamp 1682952543
transform 1 0 2852 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3770
timestamp 1682952543
transform 1 0 2860 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1682952543
transform 1 0 2788 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1682952543
transform 1 0 2804 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1682952543
transform 1 0 2796 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3809
timestamp 1682952543
transform 1 0 2804 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3843
timestamp 1682952543
transform 1 0 2804 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3780
timestamp 1682952543
transform 1 0 2836 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_3856
timestamp 1682952543
transform 1 0 2868 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3844
timestamp 1682952543
transform 1 0 2868 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1682952543
transform 1 0 2884 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3756
timestamp 1682952543
transform 1 0 2876 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1682952543
transform 1 0 2940 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1682952543
transform 1 0 2908 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3757
timestamp 1682952543
transform 1 0 2916 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3857
timestamp 1682952543
transform 1 0 2884 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3810
timestamp 1682952543
transform 1 0 2884 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3613
timestamp 1682952543
transform 1 0 3004 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1682952543
transform 1 0 2956 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1682952543
transform 1 0 2988 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3663
timestamp 1682952543
transform 1 0 2972 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1682952543
transform 1 0 3044 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_3678
timestamp 1682952543
transform 1 0 2956 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_3771
timestamp 1682952543
transform 1 0 2948 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1682952543
transform 1 0 2932 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1682952543
transform 1 0 2940 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3811
timestamp 1682952543
transform 1 0 2932 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3845
timestamp 1682952543
transform 1 0 2892 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1682952543
transform 1 0 2916 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1682952543
transform 1 0 2996 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3772
timestamp 1682952543
transform 1 0 2996 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3773
timestamp 1682952543
transform 1 0 3052 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3860
timestamp 1682952543
transform 1 0 2972 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3812
timestamp 1682952543
transform 1 0 2956 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1682952543
transform 1 0 2972 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1682952543
transform 1 0 2956 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1682952543
transform 1 0 3060 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3726
timestamp 1682952543
transform 1 0 3124 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1682952543
transform 1 0 3156 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3774
timestamp 1682952543
transform 1 0 3124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3775
timestamp 1682952543
transform 1 0 3156 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1682952543
transform 1 0 3164 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1682952543
transform 1 0 3196 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1682952543
transform 1 0 3076 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3781
timestamp 1682952543
transform 1 0 3140 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3814
timestamp 1682952543
transform 1 0 3076 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1682952543
transform 1 0 3292 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3665
timestamp 1682952543
transform 1 0 3308 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1682952543
transform 1 0 3316 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1682952543
transform 1 0 3476 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1682952543
transform 1 0 3404 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1682952543
transform 1 0 3428 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3778
timestamp 1682952543
transform 1 0 3268 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1682952543
transform 1 0 3292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3780
timestamp 1682952543
transform 1 0 3300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1682952543
transform 1 0 3308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1682952543
transform 1 0 3244 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3863
timestamp 1682952543
transform 1 0 3260 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3815
timestamp 1682952543
transform 1 0 3244 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3782
timestamp 1682952543
transform 1 0 3268 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3758
timestamp 1682952543
transform 1 0 3396 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3782
timestamp 1682952543
transform 1 0 3412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3783
timestamp 1682952543
transform 1 0 3420 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3784
timestamp 1682952543
transform 1 0 3428 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1682952543
transform 1 0 3292 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1682952543
transform 1 0 3404 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1682952543
transform 1 0 3412 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3816
timestamp 1682952543
transform 1 0 3292 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3817
timestamp 1682952543
transform 1 0 3324 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_3881
timestamp 1682952543
transform 1 0 3396 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3818
timestamp 1682952543
transform 1 0 3500 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_3882
timestamp 1682952543
transform 1 0 3516 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3849
timestamp 1682952543
transform 1 0 3476 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3730
timestamp 1682952543
transform 1 0 3532 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3785
timestamp 1682952543
transform 1 0 3540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3867
timestamp 1682952543
transform 1 0 3532 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3731
timestamp 1682952543
transform 1 0 3564 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3786
timestamp 1682952543
transform 1 0 3556 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1682952543
transform 1 0 3564 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3868
timestamp 1682952543
transform 1 0 3548 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3883
timestamp 1682952543
transform 1 0 3652 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3732
timestamp 1682952543
transform 1 0 3684 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3869
timestamp 1682952543
transform 1 0 3684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1682952543
transform 1 0 3724 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3789
timestamp 1682952543
transform 1 0 3780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3790
timestamp 1682952543
transform 1 0 3788 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3870
timestamp 1682952543
transform 1 0 3700 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3783
timestamp 1682952543
transform 1 0 3772 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3784
timestamp 1682952543
transform 1 0 3788 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1682952543
transform 1 0 3892 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1682952543
transform 1 0 4004 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1682952543
transform 1 0 3956 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3690
timestamp 1682952543
transform 1 0 4028 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1682952543
transform 1 0 3812 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3734
timestamp 1682952543
transform 1 0 3908 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3735
timestamp 1682952543
transform 1 0 3932 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_3791
timestamp 1682952543
transform 1 0 3812 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3759
timestamp 1682952543
transform 1 0 3900 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3760
timestamp 1682952543
transform 1 0 3916 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3792
timestamp 1682952543
transform 1 0 3924 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3793
timestamp 1682952543
transform 1 0 3932 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3761
timestamp 1682952543
transform 1 0 4100 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_3794
timestamp 1682952543
transform 1 0 4132 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1682952543
transform 1 0 4148 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_3871
timestamp 1682952543
transform 1 0 3796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3872
timestamp 1682952543
transform 1 0 3908 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3873
timestamp 1682952543
transform 1 0 3916 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3819
timestamp 1682952543
transform 1 0 3700 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3820
timestamp 1682952543
transform 1 0 3788 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3785
timestamp 1682952543
transform 1 0 4028 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_3874
timestamp 1682952543
transform 1 0 4036 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1682952543
transform 1 0 4148 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1682952543
transform 1 0 4220 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_3884
timestamp 1682952543
transform 1 0 3900 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3821
timestamp 1682952543
transform 1 0 3916 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3822
timestamp 1682952543
transform 1 0 3964 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_3885
timestamp 1682952543
transform 1 0 4020 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3850
timestamp 1682952543
transform 1 0 3796 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1682952543
transform 1 0 3860 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_3886
timestamp 1682952543
transform 1 0 4044 0 1 2595
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_30
timestamp 1682952543
transform 1 0 48 0 1 2570
box -10 -3 10 3
use BUFX2  BUFX2_22
timestamp 1682952543
transform -1 0 96 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_23
timestamp 1682952543
transform -1 0 120 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_24
timestamp 1682952543
transform 1 0 120 0 1 2570
box -5 -3 28 105
use INVX2  INVX2_269
timestamp 1682952543
transform -1 0 160 0 1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_239
timestamp 1682952543
transform 1 0 160 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_240
timestamp 1682952543
transform 1 0 256 0 1 2570
box -8 -3 104 105
use AOI22X1  AOI22X1_139
timestamp 1682952543
transform 1 0 352 0 1 2570
box -8 -3 46 105
use INVX2  INVX2_270
timestamp 1682952543
transform 1 0 392 0 1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_241
timestamp 1682952543
transform 1 0 408 0 1 2570
box -8 -3 104 105
use OAI22X1  OAI22X1_192
timestamp 1682952543
transform -1 0 544 0 1 2570
box -8 -3 46 105
use INVX2  INVX2_271
timestamp 1682952543
transform -1 0 560 0 1 2570
box -9 -3 26 105
use FILL  FILL_1071
timestamp 1682952543
transform 1 0 560 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_140
timestamp 1682952543
transform 1 0 568 0 1 2570
box -8 -3 46 105
use FILL  FILL_1072
timestamp 1682952543
transform 1 0 608 0 1 2570
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1682952543
transform 1 0 616 0 1 2570
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1682952543
transform 1 0 624 0 1 2570
box -8 -3 16 105
use AND2X2  AND2X2_18
timestamp 1682952543
transform -1 0 664 0 1 2570
box -8 -3 40 105
use FILL  FILL_1075
timestamp 1682952543
transform 1 0 664 0 1 2570
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1682952543
transform 1 0 672 0 1 2570
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1682952543
transform 1 0 680 0 1 2570
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1682952543
transform 1 0 688 0 1 2570
box -8 -3 16 105
use AND2X2  AND2X2_19
timestamp 1682952543
transform -1 0 728 0 1 2570
box -8 -3 40 105
use FILL  FILL_1087
timestamp 1682952543
transform 1 0 728 0 1 2570
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1682952543
transform 1 0 736 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3852
timestamp 1682952543
transform 1 0 756 0 1 2575
box -3 -3 3 3
use FILL  FILL_1091
timestamp 1682952543
transform 1 0 744 0 1 2570
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1682952543
transform 1 0 752 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3853
timestamp 1682952543
transform 1 0 780 0 1 2575
box -3 -3 3 3
use NOR2X1  NOR2X1_48
timestamp 1682952543
transform 1 0 760 0 1 2570
box -8 -3 32 105
use FILL  FILL_1095
timestamp 1682952543
transform 1 0 784 0 1 2570
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1682952543
transform 1 0 792 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3854
timestamp 1682952543
transform 1 0 812 0 1 2575
box -3 -3 3 3
use FILL  FILL_1099
timestamp 1682952543
transform 1 0 800 0 1 2570
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1682952543
transform 1 0 808 0 1 2570
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1682952543
transform 1 0 816 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3855
timestamp 1682952543
transform 1 0 868 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_194
timestamp 1682952543
transform 1 0 824 0 1 2570
box -8 -3 46 105
use FILL  FILL_1104
timestamp 1682952543
transform 1 0 864 0 1 2570
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1682952543
transform 1 0 872 0 1 2570
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1682952543
transform 1 0 880 0 1 2570
box -8 -3 16 105
use FILL  FILL_1107
timestamp 1682952543
transform 1 0 888 0 1 2570
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1682952543
transform 1 0 896 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_50
timestamp 1682952543
transform 1 0 904 0 1 2570
box -8 -3 32 105
use FILL  FILL_1115
timestamp 1682952543
transform 1 0 928 0 1 2570
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1682952543
transform 1 0 936 0 1 2570
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1682952543
transform 1 0 944 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_30
timestamp 1682952543
transform 1 0 952 0 1 2570
box -5 -3 28 105
use FILL  FILL_1121
timestamp 1682952543
transform 1 0 976 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3856
timestamp 1682952543
transform 1 0 1012 0 1 2575
box -3 -3 3 3
use BUFX2  BUFX2_31
timestamp 1682952543
transform 1 0 984 0 1 2570
box -5 -3 28 105
use FILL  FILL_1122
timestamp 1682952543
transform 1 0 1008 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3857
timestamp 1682952543
transform 1 0 1044 0 1 2575
box -3 -3 3 3
use AND2X2  AND2X2_20
timestamp 1682952543
transform -1 0 1048 0 1 2570
box -8 -3 40 105
use FILL  FILL_1123
timestamp 1682952543
transform 1 0 1048 0 1 2570
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1682952543
transform 1 0 1056 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3858
timestamp 1682952543
transform 1 0 1092 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_247
timestamp 1682952543
transform 1 0 1064 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_273
timestamp 1682952543
transform 1 0 1160 0 1 2570
box -9 -3 26 105
use FILL  FILL_1125
timestamp 1682952543
transform 1 0 1176 0 1 2570
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1682952543
transform 1 0 1184 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3859
timestamp 1682952543
transform 1 0 1204 0 1 2575
box -3 -3 3 3
use FILL  FILL_1127
timestamp 1682952543
transform 1 0 1192 0 1 2570
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1682952543
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3860
timestamp 1682952543
transform 1 0 1220 0 1 2575
box -3 -3 3 3
use FILL  FILL_1129
timestamp 1682952543
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3861
timestamp 1682952543
transform 1 0 1252 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_195
timestamp 1682952543
transform -1 0 1256 0 1 2570
box -8 -3 46 105
use FILL  FILL_1130
timestamp 1682952543
transform 1 0 1256 0 1 2570
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1682952543
transform 1 0 1264 0 1 2570
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1682952543
transform 1 0 1272 0 1 2570
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1682952543
transform 1 0 1280 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3862
timestamp 1682952543
transform 1 0 1316 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_248
timestamp 1682952543
transform -1 0 1384 0 1 2570
box -8 -3 104 105
use FILL  FILL_1134
timestamp 1682952543
transform 1 0 1384 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_32
timestamp 1682952543
transform 1 0 1392 0 1 2570
box -5 -3 28 105
use FILL  FILL_1135
timestamp 1682952543
transform 1 0 1416 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_33
timestamp 1682952543
transform 1 0 1424 0 1 2570
box -5 -3 28 105
use M3_M2  M3_M2_3863
timestamp 1682952543
transform 1 0 1468 0 1 2575
box -3 -3 3 3
use BUFX2  BUFX2_34
timestamp 1682952543
transform 1 0 1448 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_35
timestamp 1682952543
transform 1 0 1472 0 1 2570
box -5 -3 28 105
use OAI22X1  OAI22X1_196
timestamp 1682952543
transform 1 0 1496 0 1 2570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_249
timestamp 1682952543
transform 1 0 1536 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_274
timestamp 1682952543
transform -1 0 1648 0 1 2570
box -9 -3 26 105
use FILL  FILL_1136
timestamp 1682952543
transform 1 0 1648 0 1 2570
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1682952543
transform 1 0 1656 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3864
timestamp 1682952543
transform 1 0 1732 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3865
timestamp 1682952543
transform 1 0 1764 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_251
timestamp 1682952543
transform 1 0 1664 0 1 2570
box -8 -3 104 105
use FILL  FILL_1174
timestamp 1682952543
transform 1 0 1760 0 1 2570
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1682952543
transform 1 0 1768 0 1 2570
box -8 -3 16 105
use AND2X2  AND2X2_23
timestamp 1682952543
transform -1 0 1808 0 1 2570
box -8 -3 40 105
use AND2X2  AND2X2_24
timestamp 1682952543
transform -1 0 1840 0 1 2570
box -8 -3 40 105
use FILL  FILL_1176
timestamp 1682952543
transform 1 0 1840 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_19
timestamp 1682952543
transform -1 0 1880 0 1 2570
box -8 -3 40 105
use M3_M2  M3_M2_3866
timestamp 1682952543
transform 1 0 1900 0 1 2575
box -3 -3 3 3
use NAND3X1  NAND3X1_20
timestamp 1682952543
transform -1 0 1912 0 1 2570
box -8 -3 40 105
use FILL  FILL_1177
timestamp 1682952543
transform 1 0 1912 0 1 2570
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1682952543
transform 1 0 1920 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_21
timestamp 1682952543
transform -1 0 1960 0 1 2570
box -8 -3 40 105
use FILL  FILL_1179
timestamp 1682952543
transform 1 0 1960 0 1 2570
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1682952543
transform 1 0 1968 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3867
timestamp 1682952543
transform 1 0 1988 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3868
timestamp 1682952543
transform 1 0 2012 0 1 2575
box -3 -3 3 3
use NAND3X1  NAND3X1_22
timestamp 1682952543
transform -1 0 2008 0 1 2570
box -8 -3 40 105
use INVX2  INVX2_278
timestamp 1682952543
transform 1 0 2008 0 1 2570
box -9 -3 26 105
use M3_M2  M3_M2_3869
timestamp 1682952543
transform 1 0 2060 0 1 2575
box -3 -3 3 3
use NAND3X1  NAND3X1_23
timestamp 1682952543
transform 1 0 2024 0 1 2570
box -8 -3 40 105
use FILL  FILL_1181
timestamp 1682952543
transform 1 0 2056 0 1 2570
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1682952543
transform 1 0 2064 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_51
timestamp 1682952543
transform 1 0 2072 0 1 2570
box -8 -3 32 105
use FILL  FILL_1183
timestamp 1682952543
transform 1 0 2096 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3870
timestamp 1682952543
transform 1 0 2116 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_279
timestamp 1682952543
transform 1 0 2104 0 1 2570
box -9 -3 26 105
use FILL  FILL_1184
timestamp 1682952543
transform 1 0 2120 0 1 2570
box -8 -3 16 105
use AND2X2  AND2X2_25
timestamp 1682952543
transform 1 0 2128 0 1 2570
box -8 -3 40 105
use FILL  FILL_1185
timestamp 1682952543
transform 1 0 2160 0 1 2570
box -8 -3 16 105
use AND2X2  AND2X2_26
timestamp 1682952543
transform 1 0 2168 0 1 2570
box -8 -3 40 105
use FILL  FILL_1199
timestamp 1682952543
transform 1 0 2200 0 1 2570
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1682952543
transform 1 0 2208 0 1 2570
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1682952543
transform 1 0 2216 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3871
timestamp 1682952543
transform 1 0 2244 0 1 2575
box -3 -3 3 3
use AND2X2  AND2X2_27
timestamp 1682952543
transform 1 0 2224 0 1 2570
box -8 -3 40 105
use FILL  FILL_1205
timestamp 1682952543
transform 1 0 2256 0 1 2570
box -8 -3 16 105
use AND2X2  AND2X2_29
timestamp 1682952543
transform 1 0 2264 0 1 2570
box -8 -3 40 105
use FILL  FILL_1207
timestamp 1682952543
transform 1 0 2296 0 1 2570
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1682952543
transform 1 0 2304 0 1 2570
box -8 -3 16 105
use AND2X2  AND2X2_30
timestamp 1682952543
transform -1 0 2344 0 1 2570
box -8 -3 40 105
use INVX2  INVX2_284
timestamp 1682952543
transform 1 0 2344 0 1 2570
box -9 -3 26 105
use AND2X2  AND2X2_31
timestamp 1682952543
transform -1 0 2392 0 1 2570
box -8 -3 40 105
use NOR2X1  NOR2X1_52
timestamp 1682952543
transform 1 0 2392 0 1 2570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_255
timestamp 1682952543
transform -1 0 2512 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_256
timestamp 1682952543
transform 1 0 2512 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_285
timestamp 1682952543
transform 1 0 2608 0 1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_257
timestamp 1682952543
transform -1 0 2720 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_286
timestamp 1682952543
transform 1 0 2720 0 1 2570
box -9 -3 26 105
use BUFX2  BUFX2_40
timestamp 1682952543
transform 1 0 2736 0 1 2570
box -5 -3 28 105
use INVX2  INVX2_287
timestamp 1682952543
transform 1 0 2760 0 1 2570
box -9 -3 26 105
use INVX2  INVX2_288
timestamp 1682952543
transform -1 0 2792 0 1 2570
box -9 -3 26 105
use NOR2X1  NOR2X1_53
timestamp 1682952543
transform 1 0 2792 0 1 2570
box -8 -3 32 105
use NAND3X1  NAND3X1_24
timestamp 1682952543
transform 1 0 2816 0 1 2570
box -8 -3 40 105
use INVX2  INVX2_289
timestamp 1682952543
transform -1 0 2864 0 1 2570
box -9 -3 26 105
use FILL  FILL_1209
timestamp 1682952543
transform 1 0 2864 0 1 2570
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1682952543
transform 1 0 2872 0 1 2570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_0
timestamp 1682952543
transform -1 0 2936 0 1 2570
box -8 -3 64 105
use NAND2X1  NAND2X1_54
timestamp 1682952543
transform 1 0 2936 0 1 2570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_258
timestamp 1682952543
transform 1 0 2960 0 1 2570
box -8 -3 104 105
use FILL  FILL_1211
timestamp 1682952543
transform 1 0 3056 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_259
timestamp 1682952543
transform 1 0 3064 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_260
timestamp 1682952543
transform -1 0 3256 0 1 2570
box -8 -3 104 105
use AND2X2  AND2X2_32
timestamp 1682952543
transform 1 0 3256 0 1 2570
box -8 -3 40 105
use FAX1  FAX1_13
timestamp 1682952543
transform 1 0 3288 0 1 2570
box -5 -3 126 105
use FAX1  FAX1_14
timestamp 1682952543
transform 1 0 3408 0 1 2570
box -5 -3 126 105
use FILL  FILL_1212
timestamp 1682952543
transform 1 0 3528 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3872
timestamp 1682952543
transform 1 0 3548 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3873
timestamp 1682952543
transform 1 0 3564 0 1 2575
box -3 -3 3 3
use M3_M2  M3_M2_3874
timestamp 1682952543
transform 1 0 3596 0 1 2575
box -3 -3 3 3
use FILL  FILL_1213
timestamp 1682952543
transform 1 0 3536 0 1 2570
box -8 -3 16 105
use FAX1  FAX1_15
timestamp 1682952543
transform 1 0 3544 0 1 2570
box -5 -3 126 105
use FILL  FILL_1214
timestamp 1682952543
transform 1 0 3664 0 1 2570
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1682952543
transform 1 0 3672 0 1 2570
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1682952543
transform 1 0 3680 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_3875
timestamp 1682952543
transform 1 0 3708 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_261
timestamp 1682952543
transform 1 0 3688 0 1 2570
box -8 -3 104 105
use FILL  FILL_1217
timestamp 1682952543
transform 1 0 3784 0 1 2570
box -8 -3 16 105
use FAX1  FAX1_16
timestamp 1682952543
transform 1 0 3792 0 1 2570
box -5 -3 126 105
use FAX1  FAX1_17
timestamp 1682952543
transform 1 0 3912 0 1 2570
box -5 -3 126 105
use FAX1  FAX1_18
timestamp 1682952543
transform -1 0 4152 0 1 2570
box -5 -3 126 105
use top_level_VIA0  top_level_VIA0_31
timestamp 1682952543
transform 1 0 4177 0 1 2570
box -10 -3 10 3
use M3_M2  M3_M2_3876
timestamp 1682952543
transform 1 0 68 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3877
timestamp 1682952543
transform 1 0 140 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1682952543
transform 1 0 84 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3893
timestamp 1682952543
transform 1 0 84 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1682952543
transform 1 0 172 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3987
timestamp 1682952543
transform 1 0 108 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_3995
timestamp 1682952543
transform 1 0 116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3996
timestamp 1682952543
transform 1 0 164 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4010
timestamp 1682952543
transform 1 0 132 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1682952543
transform 1 0 204 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3895
timestamp 1682952543
transform 1 0 204 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1682952543
transform 1 0 188 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3988
timestamp 1682952543
transform 1 0 204 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_3896
timestamp 1682952543
transform 1 0 300 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1682952543
transform 1 0 228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3999
timestamp 1682952543
transform 1 0 284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1682952543
transform 1 0 348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4001
timestamp 1682952543
transform 1 0 380 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4060
timestamp 1682952543
transform 1 0 188 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3897
timestamp 1682952543
transform 1 0 484 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3897
timestamp 1682952543
transform 1 0 404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1682952543
transform 1 0 436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4003
timestamp 1682952543
transform 1 0 484 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3898
timestamp 1682952543
transform 1 0 508 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1682952543
transform 1 0 604 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1682952543
transform 1 0 596 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3898
timestamp 1682952543
transform 1 0 508 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1682952543
transform 1 0 604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1682952543
transform 1 0 548 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4005
timestamp 1682952543
transform 1 0 596 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4061
timestamp 1682952543
transform 1 0 500 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3989
timestamp 1682952543
transform 1 0 604 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4006
timestamp 1682952543
transform 1 0 620 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3990
timestamp 1682952543
transform 1 0 636 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4011
timestamp 1682952543
transform 1 0 644 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1682952543
transform 1 0 668 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3900
timestamp 1682952543
transform 1 0 668 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3959
timestamp 1682952543
transform 1 0 676 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1682952543
transform 1 0 716 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3901
timestamp 1682952543
transform 1 0 708 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3960
timestamp 1682952543
transform 1 0 716 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4007
timestamp 1682952543
transform 1 0 692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1682952543
transform 1 0 700 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3991
timestamp 1682952543
transform 1 0 708 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4009
timestamp 1682952543
transform 1 0 716 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4012
timestamp 1682952543
transform 1 0 692 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4062
timestamp 1682952543
transform 1 0 716 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_3887
timestamp 1682952543
transform 1 0 732 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1682952543
transform 1 0 740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1682952543
transform 1 0 748 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4078
timestamp 1682952543
transform 1 0 740 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4079
timestamp 1682952543
transform 1 0 772 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3901
timestamp 1682952543
transform 1 0 812 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4010
timestamp 1682952543
transform 1 0 812 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3878
timestamp 1682952543
transform 1 0 836 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4011
timestamp 1682952543
transform 1 0 828 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4063
timestamp 1682952543
transform 1 0 828 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_3904
timestamp 1682952543
transform 1 0 852 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4108
timestamp 1682952543
transform 1 0 852 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_3879
timestamp 1682952543
transform 1 0 876 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1682952543
transform 1 0 876 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3905
timestamp 1682952543
transform 1 0 868 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4064
timestamp 1682952543
transform 1 0 876 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3931
timestamp 1682952543
transform 1 0 900 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4012
timestamp 1682952543
transform 1 0 900 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3880
timestamp 1682952543
transform 1 0 924 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3961
timestamp 1682952543
transform 1 0 924 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4013
timestamp 1682952543
transform 1 0 924 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4013
timestamp 1682952543
transform 1 0 924 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3932
timestamp 1682952543
transform 1 0 940 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3906
timestamp 1682952543
transform 1 0 940 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4014
timestamp 1682952543
transform 1 0 956 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4014
timestamp 1682952543
transform 1 0 948 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1682952543
transform 1 0 980 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3907
timestamp 1682952543
transform 1 0 980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4015
timestamp 1682952543
transform 1 0 988 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4015
timestamp 1682952543
transform 1 0 988 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4080
timestamp 1682952543
transform 1 0 996 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3881
timestamp 1682952543
transform 1 0 1028 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_3888
timestamp 1682952543
transform 1 0 1020 0 1 2545
box -2 -2 2 2
use M3_M2  M3_M2_3962
timestamp 1682952543
transform 1 0 1012 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3908
timestamp 1682952543
transform 1 0 1060 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1682952543
transform 1 0 1068 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3963
timestamp 1682952543
transform 1 0 1092 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4016
timestamp 1682952543
transform 1 0 1028 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4017
timestamp 1682952543
transform 1 0 1036 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3992
timestamp 1682952543
transform 1 0 1044 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4018
timestamp 1682952543
transform 1 0 1052 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3993
timestamp 1682952543
transform 1 0 1060 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4019
timestamp 1682952543
transform 1 0 1078 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3994
timestamp 1682952543
transform 1 0 1084 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4020
timestamp 1682952543
transform 1 0 1092 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4016
timestamp 1682952543
transform 1 0 1052 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4065
timestamp 1682952543
transform 1 0 1060 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3882
timestamp 1682952543
transform 1 0 1108 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_3910
timestamp 1682952543
transform 1 0 1108 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4017
timestamp 1682952543
transform 1 0 1116 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4066
timestamp 1682952543
transform 1 0 1116 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1682952543
transform 1 0 1140 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1682952543
transform 1 0 1236 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3965
timestamp 1682952543
transform 1 0 1204 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3911
timestamp 1682952543
transform 1 0 1228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1682952543
transform 1 0 1140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4022
timestamp 1682952543
transform 1 0 1148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1682952543
transform 1 0 1204 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4018
timestamp 1682952543
transform 1 0 1204 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4081
timestamp 1682952543
transform 1 0 1148 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4024
timestamp 1682952543
transform 1 0 1244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3912
timestamp 1682952543
transform 1 0 1268 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1682952543
transform 1 0 1284 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4019
timestamp 1682952543
transform 1 0 1276 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4082
timestamp 1682952543
transform 1 0 1292 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_3913
timestamp 1682952543
transform 1 0 1308 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4026
timestamp 1682952543
transform 1 0 1308 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4083
timestamp 1682952543
transform 1 0 1308 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_3914
timestamp 1682952543
transform 1 0 1324 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3903
timestamp 1682952543
transform 1 0 1340 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3915
timestamp 1682952543
transform 1 0 1340 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3904
timestamp 1682952543
transform 1 0 1372 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3934
timestamp 1682952543
transform 1 0 1364 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3966
timestamp 1682952543
transform 1 0 1356 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3916
timestamp 1682952543
transform 1 0 1364 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1682952543
transform 1 0 1356 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4084
timestamp 1682952543
transform 1 0 1364 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3935
timestamp 1682952543
transform 1 0 1404 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3917
timestamp 1682952543
transform 1 0 1404 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3883
timestamp 1682952543
transform 1 0 1420 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4028
timestamp 1682952543
transform 1 0 1412 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4020
timestamp 1682952543
transform 1 0 1412 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4085
timestamp 1682952543
transform 1 0 1412 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3967
timestamp 1682952543
transform 1 0 1444 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4029
timestamp 1682952543
transform 1 0 1444 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1682952543
transform 1 0 1452 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4021
timestamp 1682952543
transform 1 0 1452 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3884
timestamp 1682952543
transform 1 0 1468 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3968
timestamp 1682952543
transform 1 0 1476 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3918
timestamp 1682952543
transform 1 0 1484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1682952543
transform 1 0 1492 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1682952543
transform 1 0 1516 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4032
timestamp 1682952543
transform 1 0 1564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4033
timestamp 1682952543
transform 1 0 1572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1682952543
transform 1 0 1580 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4022
timestamp 1682952543
transform 1 0 1564 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1682952543
transform 1 0 1596 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3920
timestamp 1682952543
transform 1 0 1596 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1682952543
transform 1 0 1588 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1682952543
transform 1 0 1628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1682952543
transform 1 0 1620 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4037
timestamp 1682952543
transform 1 0 1636 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4023
timestamp 1682952543
transform 1 0 1620 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_3922
timestamp 1682952543
transform 1 0 1676 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3937
timestamp 1682952543
transform 1 0 1708 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1682952543
transform 1 0 1724 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3923
timestamp 1682952543
transform 1 0 1708 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3969
timestamp 1682952543
transform 1 0 1716 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3924
timestamp 1682952543
transform 1 0 1724 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4038
timestamp 1682952543
transform 1 0 1692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1682952543
transform 1 0 1700 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4040
timestamp 1682952543
transform 1 0 1708 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4024
timestamp 1682952543
transform 1 0 1692 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3970
timestamp 1682952543
transform 1 0 1756 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4041
timestamp 1682952543
transform 1 0 1756 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4042
timestamp 1682952543
transform 1 0 1772 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4025
timestamp 1682952543
transform 1 0 1764 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4086
timestamp 1682952543
transform 1 0 1756 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4087
timestamp 1682952543
transform 1 0 1780 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1682952543
transform 1 0 1876 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1682952543
transform 1 0 1900 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3925
timestamp 1682952543
transform 1 0 1796 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3926
timestamp 1682952543
transform 1 0 1804 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3971
timestamp 1682952543
transform 1 0 1812 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3927
timestamp 1682952543
transform 1 0 1900 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3905
timestamp 1682952543
transform 1 0 1980 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3941
timestamp 1682952543
transform 1 0 1996 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3928
timestamp 1682952543
transform 1 0 1996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1682952543
transform 1 0 1812 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1682952543
transform 1 0 1820 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1682952543
transform 1 0 1852 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4046
timestamp 1682952543
transform 1 0 1916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1682952543
transform 1 0 1964 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4026
timestamp 1682952543
transform 1 0 1812 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4027
timestamp 1682952543
transform 1 0 1852 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3885
timestamp 1682952543
transform 1 0 2060 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1682952543
transform 1 0 2044 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1682952543
transform 1 0 2092 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1682952543
transform 1 0 2028 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3908
timestamp 1682952543
transform 1 0 2124 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3929
timestamp 1682952543
transform 1 0 2028 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3930
timestamp 1682952543
transform 1 0 2116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1682952543
transform 1 0 2124 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1682952543
transform 1 0 2140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3933
timestamp 1682952543
transform 1 0 2148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4048
timestamp 1682952543
transform 1 0 2076 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1682952543
transform 1 0 2108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4050
timestamp 1682952543
transform 1 0 2116 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4051
timestamp 1682952543
transform 1 0 2132 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4052
timestamp 1682952543
transform 1 0 2148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4053
timestamp 1682952543
transform 1 0 2156 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4028
timestamp 1682952543
transform 1 0 2076 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1682952543
transform 1 0 2052 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4089
timestamp 1682952543
transform 1 0 2092 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4090
timestamp 1682952543
transform 1 0 2108 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1682952543
transform 1 0 2140 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4029
timestamp 1682952543
transform 1 0 2156 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1682952543
transform 1 0 2156 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1682952543
transform 1 0 2172 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3934
timestamp 1682952543
transform 1 0 2188 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4093
timestamp 1682952543
transform 1 0 2188 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3943
timestamp 1682952543
transform 1 0 2204 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1682952543
transform 1 0 2228 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3935
timestamp 1682952543
transform 1 0 2220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1682952543
transform 1 0 2220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1682952543
transform 1 0 2236 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4030
timestamp 1682952543
transform 1 0 2236 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3973
timestamp 1682952543
transform 1 0 2260 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4056
timestamp 1682952543
transform 1 0 2260 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1682952543
transform 1 0 2276 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1682952543
transform 1 0 2276 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3886
timestamp 1682952543
transform 1 0 2308 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3974
timestamp 1682952543
transform 1 0 2316 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3937
timestamp 1682952543
transform 1 0 2324 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1682952543
transform 1 0 2300 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4031
timestamp 1682952543
transform 1 0 2300 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4059
timestamp 1682952543
transform 1 0 2324 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3975
timestamp 1682952543
transform 1 0 2340 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4060
timestamp 1682952543
transform 1 0 2340 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4094
timestamp 1682952543
transform 1 0 2332 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3909
timestamp 1682952543
transform 1 0 2372 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3938
timestamp 1682952543
transform 1 0 2372 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3976
timestamp 1682952543
transform 1 0 2380 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1682952543
transform 1 0 2404 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1682952543
transform 1 0 2396 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1682952543
transform 1 0 2412 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3939
timestamp 1682952543
transform 1 0 2404 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1682952543
transform 1 0 2412 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3941
timestamp 1682952543
transform 1 0 2428 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1682952543
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1682952543
transform 1 0 2396 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4032
timestamp 1682952543
transform 1 0 2388 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1682952543
transform 1 0 2380 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_3942
timestamp 1682952543
transform 1 0 2444 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1682952543
transform 1 0 2420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1682952543
transform 1 0 2436 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4033
timestamp 1682952543
transform 1 0 2436 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4096
timestamp 1682952543
transform 1 0 2420 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3977
timestamp 1682952543
transform 1 0 2452 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4097
timestamp 1682952543
transform 1 0 2444 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3911
timestamp 1682952543
transform 1 0 2484 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3943
timestamp 1682952543
transform 1 0 2484 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3978
timestamp 1682952543
transform 1 0 2492 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3887
timestamp 1682952543
transform 1 0 2524 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1682952543
transform 1 0 2532 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3944
timestamp 1682952543
transform 1 0 2516 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3945
timestamp 1682952543
transform 1 0 2524 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1682952543
transform 1 0 2476 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4066
timestamp 1682952543
transform 1 0 2492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1682952543
transform 1 0 2508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4068
timestamp 1682952543
transform 1 0 2524 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4034
timestamp 1682952543
transform 1 0 2524 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3912
timestamp 1682952543
transform 1 0 2556 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4069
timestamp 1682952543
transform 1 0 2548 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3946
timestamp 1682952543
transform 1 0 2556 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3948
timestamp 1682952543
transform 1 0 2596 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3947
timestamp 1682952543
transform 1 0 2596 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1682952543
transform 1 0 2604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4070
timestamp 1682952543
transform 1 0 2572 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1682952543
transform 1 0 2588 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3995
timestamp 1682952543
transform 1 0 2596 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4072
timestamp 1682952543
transform 1 0 2604 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4067
timestamp 1682952543
transform 1 0 2572 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4098
timestamp 1682952543
transform 1 0 2572 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3996
timestamp 1682952543
transform 1 0 2612 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1682952543
transform 1 0 2604 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3913
timestamp 1682952543
transform 1 0 2652 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1682952543
transform 1 0 2628 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3949
timestamp 1682952543
transform 1 0 2628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3950
timestamp 1682952543
transform 1 0 2636 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1682952543
transform 1 0 2652 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3997
timestamp 1682952543
transform 1 0 2636 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_3952
timestamp 1682952543
transform 1 0 2668 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1682952543
transform 1 0 2644 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4074
timestamp 1682952543
transform 1 0 2660 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4036
timestamp 1682952543
transform 1 0 2644 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4068
timestamp 1682952543
transform 1 0 2652 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4037
timestamp 1682952543
transform 1 0 2668 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1682952543
transform 1 0 2660 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3914
timestamp 1682952543
transform 1 0 2676 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1682952543
transform 1 0 2676 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4069
timestamp 1682952543
transform 1 0 2676 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1682952543
transform 1 0 2708 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1682952543
transform 1 0 2772 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1682952543
transform 1 0 2796 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_3953
timestamp 1682952543
transform 1 0 2708 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3979
timestamp 1682952543
transform 1 0 2788 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4075
timestamp 1682952543
transform 1 0 2692 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1682952543
transform 1 0 2732 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3998
timestamp 1682952543
transform 1 0 2780 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4077
timestamp 1682952543
transform 1 0 2788 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4078
timestamp 1682952543
transform 1 0 2796 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4038
timestamp 1682952543
transform 1 0 2692 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1682952543
transform 1 0 2732 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1682952543
transform 1 0 2796 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3891
timestamp 1682952543
transform 1 0 2812 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1682952543
transform 1 0 2812 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3954
timestamp 1682952543
transform 1 0 2812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1682952543
transform 1 0 2828 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4079
timestamp 1682952543
transform 1 0 2820 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3999
timestamp 1682952543
transform 1 0 2828 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4080
timestamp 1682952543
transform 1 0 2836 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3916
timestamp 1682952543
transform 1 0 2884 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3951
timestamp 1682952543
transform 1 0 2868 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3956
timestamp 1682952543
transform 1 0 2852 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1682952543
transform 1 0 2860 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4000
timestamp 1682952543
transform 1 0 2860 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4081
timestamp 1682952543
transform 1 0 2868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_3958
timestamp 1682952543
transform 1 0 2892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1682952543
transform 1 0 2916 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3892
timestamp 1682952543
transform 1 0 2964 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3917
timestamp 1682952543
transform 1 0 2956 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1682952543
transform 1 0 2948 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3889
timestamp 1682952543
transform 1 0 2956 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1682952543
transform 1 0 2948 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3961
timestamp 1682952543
transform 1 0 2964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1682952543
transform 1 0 2988 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1682952543
transform 1 0 3004 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4082
timestamp 1682952543
transform 1 0 2892 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4083
timestamp 1682952543
transform 1 0 2900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1682952543
transform 1 0 2916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4131
timestamp 1682952543
transform 1 0 2884 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4070
timestamp 1682952543
transform 1 0 2876 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4001
timestamp 1682952543
transform 1 0 2932 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4085
timestamp 1682952543
transform 1 0 2940 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4132
timestamp 1682952543
transform 1 0 2916 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4071
timestamp 1682952543
transform 1 0 2908 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1682952543
transform 1 0 2900 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1682952543
transform 1 0 2884 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4102
timestamp 1682952543
transform 1 0 2956 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1682952543
transform 1 0 2948 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_3964
timestamp 1682952543
transform 1 0 3052 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1682952543
transform 1 0 2988 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4087
timestamp 1682952543
transform 1 0 3004 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4002
timestamp 1682952543
transform 1 0 3028 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4088
timestamp 1682952543
transform 1 0 3036 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4040
timestamp 1682952543
transform 1 0 3004 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1682952543
transform 1 0 3036 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4072
timestamp 1682952543
transform 1 0 2988 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4073
timestamp 1682952543
transform 1 0 3044 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4103
timestamp 1682952543
transform 1 0 3020 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1682952543
transform 1 0 3084 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1682952543
transform 1 0 3132 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3918
timestamp 1682952543
transform 1 0 3164 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1682952543
transform 1 0 3188 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3965
timestamp 1682952543
transform 1 0 3108 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1682952543
transform 1 0 3116 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3967
timestamp 1682952543
transform 1 0 3132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1682952543
transform 1 0 3148 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3969
timestamp 1682952543
transform 1 0 3156 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1682952543
transform 1 0 3172 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3971
timestamp 1682952543
transform 1 0 3180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1682952543
transform 1 0 3068 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4090
timestamp 1682952543
transform 1 0 3084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1682952543
transform 1 0 3092 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4092
timestamp 1682952543
transform 1 0 3100 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4042
timestamp 1682952543
transform 1 0 3068 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4003
timestamp 1682952543
transform 1 0 3116 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4093
timestamp 1682952543
transform 1 0 3124 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4004
timestamp 1682952543
transform 1 0 3132 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4094
timestamp 1682952543
transform 1 0 3148 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1682952543
transform 1 0 3164 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4043
timestamp 1682952543
transform 1 0 3116 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1682952543
transform 1 0 3172 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4096
timestamp 1682952543
transform 1 0 3188 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4044
timestamp 1682952543
transform 1 0 3156 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4074
timestamp 1682952543
transform 1 0 3164 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1682952543
transform 1 0 3156 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1682952543
transform 1 0 3172 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_3890
timestamp 1682952543
transform 1 0 3204 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3972
timestamp 1682952543
transform 1 0 3220 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1682952543
transform 1 0 3196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1682952543
transform 1 0 3204 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3920
timestamp 1682952543
transform 1 0 3244 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3921
timestamp 1682952543
transform 1 0 3276 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3973
timestamp 1682952543
transform 1 0 3244 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3980
timestamp 1682952543
transform 1 0 3324 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3974
timestamp 1682952543
transform 1 0 3332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1682952543
transform 1 0 3228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1682952543
transform 1 0 3284 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4101
timestamp 1682952543
transform 1 0 3332 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4045
timestamp 1682952543
transform 1 0 3244 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4046
timestamp 1682952543
transform 1 0 3268 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1682952543
transform 1 0 3252 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1682952543
transform 1 0 3324 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_3955
timestamp 1682952543
transform 1 0 3380 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1682952543
transform 1 0 3500 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3894
timestamp 1682952543
transform 1 0 3516 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3922
timestamp 1682952543
transform 1 0 3412 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3923
timestamp 1682952543
transform 1 0 3436 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3956
timestamp 1682952543
transform 1 0 3412 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3975
timestamp 1682952543
transform 1 0 3380 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3981
timestamp 1682952543
transform 1 0 3396 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3976
timestamp 1682952543
transform 1 0 3420 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4102
timestamp 1682952543
transform 1 0 3380 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1682952543
transform 1 0 3396 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4006
timestamp 1682952543
transform 1 0 3404 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3982
timestamp 1682952543
transform 1 0 3428 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3977
timestamp 1682952543
transform 1 0 3516 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3895
timestamp 1682952543
transform 1 0 3604 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1682952543
transform 1 0 3644 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_3891
timestamp 1682952543
transform 1 0 3556 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3978
timestamp 1682952543
transform 1 0 3540 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4104
timestamp 1682952543
transform 1 0 3412 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1682952543
transform 1 0 3428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1682952543
transform 1 0 3436 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1682952543
transform 1 0 3492 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1682952543
transform 1 0 3532 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4047
timestamp 1682952543
transform 1 0 3396 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1682952543
transform 1 0 3420 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1682952543
transform 1 0 3388 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4114
timestamp 1682952543
transform 1 0 3388 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4049
timestamp 1682952543
transform 1 0 3492 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3983
timestamp 1682952543
transform 1 0 3556 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_3957
timestamp 1682952543
transform 1 0 3660 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3979
timestamp 1682952543
transform 1 0 3644 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3980
timestamp 1682952543
transform 1 0 3660 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1682952543
transform 1 0 3556 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1682952543
transform 1 0 3564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1682952543
transform 1 0 3620 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4050
timestamp 1682952543
transform 1 0 3564 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1682952543
transform 1 0 3548 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1682952543
transform 1 0 3724 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_3981
timestamp 1682952543
transform 1 0 3708 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_3984
timestamp 1682952543
transform 1 0 3740 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3982
timestamp 1682952543
transform 1 0 3756 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1682952543
transform 1 0 3772 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3984
timestamp 1682952543
transform 1 0 3788 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1682952543
transform 1 0 3708 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1682952543
transform 1 0 3724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4114
timestamp 1682952543
transform 1 0 3740 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1682952543
transform 1 0 3748 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1682952543
transform 1 0 3764 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4051
timestamp 1682952543
transform 1 0 3708 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1682952543
transform 1 0 3692 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4007
timestamp 1682952543
transform 1 0 3772 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_3985
timestamp 1682952543
transform 1 0 3796 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_3985
timestamp 1682952543
transform 1 0 3804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4117
timestamp 1682952543
transform 1 0 3780 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1682952543
transform 1 0 3796 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4052
timestamp 1682952543
transform 1 0 3748 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4107
timestamp 1682952543
transform 1 0 3764 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1682952543
transform 1 0 3756 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_3986
timestamp 1682952543
transform 1 0 3860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3987
timestamp 1682952543
transform 1 0 3868 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1682952543
transform 1 0 3884 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1682952543
transform 1 0 3844 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_3986
timestamp 1682952543
transform 1 0 3892 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4120
timestamp 1682952543
transform 1 0 3876 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1682952543
transform 1 0 3892 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4008
timestamp 1682952543
transform 1 0 3900 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4133
timestamp 1682952543
transform 1 0 3804 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4053
timestamp 1682952543
transform 1 0 3836 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4054
timestamp 1682952543
transform 1 0 3860 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4055
timestamp 1682952543
transform 1 0 3884 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1682952543
transform 1 0 3804 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4077
timestamp 1682952543
transform 1 0 3828 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4116
timestamp 1682952543
transform 1 0 3852 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_3989
timestamp 1682952543
transform 1 0 3964 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1682952543
transform 1 0 3972 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1682952543
transform 1 0 3996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1682952543
transform 1 0 4004 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4122
timestamp 1682952543
transform 1 0 3940 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4123
timestamp 1682952543
transform 1 0 3964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1682952543
transform 1 0 3988 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4009
timestamp 1682952543
transform 1 0 3996 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4125
timestamp 1682952543
transform 1 0 4012 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4056
timestamp 1682952543
transform 1 0 3940 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4057
timestamp 1682952543
transform 1 0 3964 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4117
timestamp 1682952543
transform 1 0 3972 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_3892
timestamp 1682952543
transform 1 0 4028 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_3993
timestamp 1682952543
transform 1 0 4044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4126
timestamp 1682952543
transform 1 0 4020 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1682952543
transform 1 0 4028 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4058
timestamp 1682952543
transform 1 0 4012 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_3924
timestamp 1682952543
transform 1 0 4116 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_3925
timestamp 1682952543
transform 1 0 4148 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_3994
timestamp 1682952543
transform 1 0 4140 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4128
timestamp 1682952543
transform 1 0 4052 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1682952543
transform 1 0 4060 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1682952543
transform 1 0 4116 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4059
timestamp 1682952543
transform 1 0 4060 0 1 2515
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_32
timestamp 1682952543
transform 1 0 24 0 1 2470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_242
timestamp 1682952543
transform 1 0 72 0 -1 2570
box -8 -3 104 105
use BUFX2  BUFX2_25
timestamp 1682952543
transform -1 0 192 0 -1 2570
box -5 -3 28 105
use M3_M2  M3_M2_4118
timestamp 1682952543
transform 1 0 252 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_243
timestamp 1682952543
transform 1 0 192 0 -1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_244
timestamp 1682952543
transform 1 0 288 0 -1 2570
box -8 -3 104 105
use FILL  FILL_1076
timestamp 1682952543
transform 1 0 384 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_245
timestamp 1682952543
transform 1 0 392 0 -1 2570
box -8 -3 104 105
use FILL  FILL_1077
timestamp 1682952543
transform 1 0 488 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_246
timestamp 1682952543
transform 1 0 496 0 -1 2570
box -8 -3 104 105
use FILL  FILL_1078
timestamp 1682952543
transform 1 0 592 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_26
timestamp 1682952543
transform -1 0 624 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1079
timestamp 1682952543
transform 1 0 624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1682952543
transform 1 0 632 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4119
timestamp 1682952543
transform 1 0 668 0 1 2475
box -3 -3 3 3
use BUFX2  BUFX2_27
timestamp 1682952543
transform -1 0 664 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1081
timestamp 1682952543
transform 1 0 664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1682952543
transform 1 0 672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1682952543
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_193
timestamp 1682952543
transform 1 0 688 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1088
timestamp 1682952543
transform 1 0 728 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1682952543
transform 1 0 736 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1682952543
transform 1 0 744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1094
timestamp 1682952543
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_49
timestamp 1682952543
transform 1 0 760 0 -1 2570
box -8 -3 32 105
use FILL  FILL_1096
timestamp 1682952543
transform 1 0 784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1682952543
transform 1 0 792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1682952543
transform 1 0 800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1682952543
transform 1 0 808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1682952543
transform 1 0 816 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_272
timestamp 1682952543
transform -1 0 840 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1109
timestamp 1682952543
transform 1 0 840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1682952543
transform 1 0 848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1682952543
transform 1 0 856 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_28
timestamp 1682952543
transform -1 0 888 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1112
timestamp 1682952543
transform 1 0 888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1682952543
transform 1 0 896 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1682952543
transform 1 0 904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1682952543
transform 1 0 912 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_29
timestamp 1682952543
transform 1 0 920 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1120
timestamp 1682952543
transform 1 0 944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1682952543
transform 1 0 952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1682952543
transform 1 0 960 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4120
timestamp 1682952543
transform 1 0 980 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_141
timestamp 1682952543
transform 1 0 968 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1139
timestamp 1682952543
transform 1 0 1008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1682952543
transform 1 0 1016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1682952543
transform 1 0 1024 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_21
timestamp 1682952543
transform -1 0 1064 0 -1 2570
box -8 -3 40 105
use M3_M2  M3_M2_4121
timestamp 1682952543
transform 1 0 1076 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4122
timestamp 1682952543
transform 1 0 1092 0 1 2475
box -3 -3 3 3
use AND2X2  AND2X2_22
timestamp 1682952543
transform 1 0 1064 0 -1 2570
box -8 -3 40 105
use M3_M2  M3_M2_4123
timestamp 1682952543
transform 1 0 1108 0 1 2475
box -3 -3 3 3
use FILL  FILL_1142
timestamp 1682952543
transform 1 0 1096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1682952543
transform 1 0 1104 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_275
timestamp 1682952543
transform 1 0 1112 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1144
timestamp 1682952543
transform 1 0 1128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1682952543
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_250
timestamp 1682952543
transform -1 0 1240 0 -1 2570
box -8 -3 104 105
use FILL  FILL_1146
timestamp 1682952543
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1682952543
transform 1 0 1248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1682952543
transform 1 0 1256 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_142
timestamp 1682952543
transform -1 0 1304 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1149
timestamp 1682952543
transform 1 0 1304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1682952543
transform 1 0 1312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1682952543
transform 1 0 1320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1682952543
transform 1 0 1328 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_36
timestamp 1682952543
transform -1 0 1360 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1153
timestamp 1682952543
transform 1 0 1360 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_37
timestamp 1682952543
transform -1 0 1392 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1154
timestamp 1682952543
transform 1 0 1392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1682952543
transform 1 0 1400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1682952543
transform 1 0 1408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1682952543
transform 1 0 1416 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_38
timestamp 1682952543
transform -1 0 1448 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1158
timestamp 1682952543
transform 1 0 1448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1682952543
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_39
timestamp 1682952543
transform 1 0 1464 0 -1 2570
box -5 -3 28 105
use FILL  FILL_1160
timestamp 1682952543
transform 1 0 1488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1682952543
transform 1 0 1496 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_276
timestamp 1682952543
transform 1 0 1504 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1162
timestamp 1682952543
transform 1 0 1520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1682952543
transform 1 0 1528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1682952543
transform 1 0 1536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1682952543
transform 1 0 1544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1682952543
transform 1 0 1552 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_277
timestamp 1682952543
transform 1 0 1560 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1167
timestamp 1682952543
transform 1 0 1576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1682952543
transform 1 0 1584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1682952543
transform 1 0 1592 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4124
timestamp 1682952543
transform 1 0 1644 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_143
timestamp 1682952543
transform 1 0 1600 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1170
timestamp 1682952543
transform 1 0 1640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1682952543
transform 1 0 1648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1682952543
transform 1 0 1656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1682952543
transform 1 0 1664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1682952543
transform 1 0 1672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1682952543
transform 1 0 1680 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4125
timestamp 1682952543
transform 1 0 1708 0 1 2475
box -3 -3 3 3
use INVX2  INVX2_280
timestamp 1682952543
transform 1 0 1688 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1189
timestamp 1682952543
transform 1 0 1704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1682952543
transform 1 0 1712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1682952543
transform 1 0 1720 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4126
timestamp 1682952543
transform 1 0 1740 0 1 2475
box -3 -3 3 3
use FILL  FILL_1192
timestamp 1682952543
transform 1 0 1728 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4127
timestamp 1682952543
transform 1 0 1780 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_144
timestamp 1682952543
transform 1 0 1736 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1193
timestamp 1682952543
transform 1 0 1776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1682952543
transform 1 0 1784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1682952543
transform 1 0 1792 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_281
timestamp 1682952543
transform 1 0 1800 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_252
timestamp 1682952543
transform -1 0 1912 0 -1 2570
box -8 -3 104 105
use M3_M2  M3_M2_4128
timestamp 1682952543
transform 1 0 1948 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4129
timestamp 1682952543
transform 1 0 1988 0 1 2475
box -3 -3 3 3
use M3_M2  M3_M2_4130
timestamp 1682952543
transform 1 0 2004 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_253
timestamp 1682952543
transform -1 0 2008 0 -1 2570
box -8 -3 104 105
use FILL  FILL_1196
timestamp 1682952543
transform 1 0 2008 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_254
timestamp 1682952543
transform 1 0 2016 0 -1 2570
box -8 -3 104 105
use M3_M2  M3_M2_4131
timestamp 1682952543
transform 1 0 2148 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_145
timestamp 1682952543
transform 1 0 2112 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1197
timestamp 1682952543
transform 1 0 2152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1682952543
transform 1 0 2160 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4132
timestamp 1682952543
transform 1 0 2188 0 1 2475
box -3 -3 3 3
use INVX2  INVX2_282
timestamp 1682952543
transform 1 0 2168 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1202
timestamp 1682952543
transform 1 0 2184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1682952543
transform 1 0 2192 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_283
timestamp 1682952543
transform 1 0 2200 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1204
timestamp 1682952543
transform 1 0 2216 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_28
timestamp 1682952543
transform 1 0 2224 0 -1 2570
box -8 -3 40 105
use FILL  FILL_1206
timestamp 1682952543
transform 1 0 2256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1682952543
transform 1 0 2264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1682952543
transform 1 0 2272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1682952543
transform 1 0 2280 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_33
timestamp 1682952543
transform 1 0 2288 0 -1 2570
box -8 -3 40 105
use FILL  FILL_1221
timestamp 1682952543
transform 1 0 2320 0 -1 2570
box -8 -3 16 105
use AND2X2  AND2X2_34
timestamp 1682952543
transform 1 0 2328 0 -1 2570
box -8 -3 40 105
use FILL  FILL_1222
timestamp 1682952543
transform 1 0 2360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1682952543
transform 1 0 2368 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4133
timestamp 1682952543
transform 1 0 2388 0 1 2475
box -3 -3 3 3
use INVX2  INVX2_290
timestamp 1682952543
transform 1 0 2376 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1224
timestamp 1682952543
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_146
timestamp 1682952543
transform 1 0 2400 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1225
timestamp 1682952543
transform 1 0 2440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1682952543
transform 1 0 2448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1682952543
transform 1 0 2456 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_291
timestamp 1682952543
transform 1 0 2464 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1228
timestamp 1682952543
transform 1 0 2480 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_147
timestamp 1682952543
transform 1 0 2488 0 -1 2570
box -8 -3 46 105
use INVX2  INVX2_292
timestamp 1682952543
transform 1 0 2528 0 -1 2570
box -9 -3 26 105
use FILL  FILL_1229
timestamp 1682952543
transform 1 0 2544 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1682952543
transform 1 0 2552 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1231
timestamp 1682952543
transform 1 0 2560 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_148
timestamp 1682952543
transform 1 0 2568 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1232
timestamp 1682952543
transform 1 0 2608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1682952543
transform 1 0 2616 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4134
timestamp 1682952543
transform 1 0 2668 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_149
timestamp 1682952543
transform -1 0 2664 0 -1 2570
box -8 -3 46 105
use FILL  FILL_1234
timestamp 1682952543
transform 1 0 2664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1682952543
transform 1 0 2672 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4135
timestamp 1682952543
transform 1 0 2700 0 1 2475
box -3 -3 3 3
use INVX2  INVX2_293
timestamp 1682952543
transform 1 0 2680 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_262
timestamp 1682952543
transform 1 0 2696 0 -1 2570
box -8 -3 104 105
use BUFX2  BUFX2_41
timestamp 1682952543
transform 1 0 2792 0 -1 2570
box -5 -3 28 105
use INVX2  INVX2_294
timestamp 1682952543
transform -1 0 2832 0 -1 2570
box -9 -3 26 105
use BUFX2  BUFX2_42
timestamp 1682952543
transform 1 0 2832 0 -1 2570
box -5 -3 28 105
use OAI21X1  OAI21X1_52
timestamp 1682952543
transform 1 0 2856 0 -1 2570
box -8 -3 34 105
use OAI21X1  OAI21X1_53
timestamp 1682952543
transform 1 0 2888 0 -1 2570
box -8 -3 34 105
use AND2X2  AND2X2_35
timestamp 1682952543
transform -1 0 2952 0 -1 2570
box -8 -3 40 105
use OR2X1  OR2X1_1
timestamp 1682952543
transform 1 0 2952 0 -1 2570
box -8 -3 40 105
use INVX2  INVX2_295
timestamp 1682952543
transform 1 0 2984 0 -1 2570
box -9 -3 26 105
use M3_M2  M3_M2_4136
timestamp 1682952543
transform 1 0 3020 0 1 2475
box -3 -3 3 3
use XNOR2X1  XNOR2X1_1
timestamp 1682952543
transform 1 0 3000 0 -1 2570
box -8 -3 64 105
use AND2X2  AND2X2_36
timestamp 1682952543
transform 1 0 3056 0 -1 2570
box -8 -3 40 105
use INVX2  INVX2_296
timestamp 1682952543
transform -1 0 3104 0 -1 2570
box -9 -3 26 105
use AOI22X1  AOI22X1_150
timestamp 1682952543
transform 1 0 3104 0 -1 2570
box -8 -3 46 105
use M3_M2  M3_M2_4137
timestamp 1682952543
transform 1 0 3164 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_151
timestamp 1682952543
transform 1 0 3144 0 -1 2570
box -8 -3 46 105
use INVX2  INVX2_297
timestamp 1682952543
transform 1 0 3184 0 -1 2570
box -9 -3 26 105
use AOI21X1  AOI21X1_14
timestamp 1682952543
transform -1 0 3232 0 -1 2570
box -7 -3 39 105
use M3_M2  M3_M2_4138
timestamp 1682952543
transform 1 0 3332 0 1 2475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_263
timestamp 1682952543
transform 1 0 3232 0 -1 2570
box -8 -3 104 105
use XOR2X1  XOR2X1_3
timestamp 1682952543
transform 1 0 3328 0 -1 2570
box -8 -3 64 105
use M3_M2  M3_M2_4139
timestamp 1682952543
transform 1 0 3412 0 1 2475
box -3 -3 3 3
use AND2X2  AND2X2_37
timestamp 1682952543
transform 1 0 3384 0 -1 2570
box -8 -3 40 105
use INVX2  INVX2_298
timestamp 1682952543
transform 1 0 3416 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_264
timestamp 1682952543
transform -1 0 3528 0 -1 2570
box -8 -3 104 105
use AOI21X1  AOI21X1_15
timestamp 1682952543
transform 1 0 3528 0 -1 2570
box -7 -3 39 105
use DFFNEGX1  DFFNEGX1_265
timestamp 1682952543
transform -1 0 3656 0 -1 2570
box -8 -3 104 105
use XOR2X1  XOR2X1_4
timestamp 1682952543
transform 1 0 3656 0 -1 2570
box -8 -3 64 105
use AND2X2  AND2X2_38
timestamp 1682952543
transform 1 0 3712 0 -1 2570
box -8 -3 40 105
use AOI22X1  AOI22X1_152
timestamp 1682952543
transform 1 0 3744 0 -1 2570
box -8 -3 46 105
use NAND2X1  NAND2X1_55
timestamp 1682952543
transform 1 0 3784 0 -1 2570
box -8 -3 32 105
use M3_M2  M3_M2_4140
timestamp 1682952543
transform 1 0 3820 0 1 2475
box -3 -3 3 3
use XOR2X1  XOR2X1_5
timestamp 1682952543
transform 1 0 3808 0 -1 2570
box -8 -3 64 105
use INVX2  INVX2_299
timestamp 1682952543
transform 1 0 3864 0 -1 2570
box -9 -3 26 105
use AND2X2  AND2X2_39
timestamp 1682952543
transform 1 0 3880 0 -1 2570
box -8 -3 40 105
use XOR2X1  XOR2X1_6
timestamp 1682952543
transform -1 0 3968 0 -1 2570
box -8 -3 64 105
use AOI22X1  AOI22X1_153
timestamp 1682952543
transform 1 0 3968 0 -1 2570
box -8 -3 46 105
use M3_M2  M3_M2_4141
timestamp 1682952543
transform 1 0 4028 0 1 2475
box -3 -3 3 3
use INVX2  INVX2_300
timestamp 1682952543
transform 1 0 4008 0 -1 2570
box -9 -3 26 105
use AOI21X1  AOI21X1_16
timestamp 1682952543
transform -1 0 4056 0 -1 2570
box -7 -3 39 105
use DFFNEGX1  DFFNEGX1_266
timestamp 1682952543
transform -1 0 4152 0 -1 2570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_33
timestamp 1682952543
transform 1 0 4201 0 1 2470
box -10 -3 10 3
use M3_M2  M3_M2_4206
timestamp 1682952543
transform 1 0 108 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4227
timestamp 1682952543
transform 1 0 100 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4149
timestamp 1682952543
transform 1 0 116 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4142
timestamp 1682952543
transform 1 0 124 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4183
timestamp 1682952543
transform 1 0 172 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4207
timestamp 1682952543
transform 1 0 164 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4228
timestamp 1682952543
transform 1 0 140 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4277
timestamp 1682952543
transform 1 0 124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4150
timestamp 1682952543
transform 1 0 140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4151
timestamp 1682952543
transform 1 0 148 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4270
timestamp 1682952543
transform 1 0 156 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4152
timestamp 1682952543
transform 1 0 164 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4271
timestamp 1682952543
transform 1 0 172 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4278
timestamp 1682952543
transform 1 0 140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1682952543
transform 1 0 156 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4329
timestamp 1682952543
transform 1 0 148 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1682952543
transform 1 0 172 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1682952543
transform 1 0 188 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4153
timestamp 1682952543
transform 1 0 188 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4272
timestamp 1682952543
transform 1 0 196 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4280
timestamp 1682952543
transform 1 0 196 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4229
timestamp 1682952543
transform 1 0 244 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4154
timestamp 1682952543
transform 1 0 228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4155
timestamp 1682952543
transform 1 0 244 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4273
timestamp 1682952543
transform 1 0 252 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4156
timestamp 1682952543
transform 1 0 260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1682952543
transform 1 0 276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4158
timestamp 1682952543
transform 1 0 284 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4281
timestamp 1682952543
transform 1 0 244 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1682952543
transform 1 0 252 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4331
timestamp 1682952543
transform 1 0 276 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4164
timestamp 1682952543
transform 1 0 324 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1682952543
transform 1 0 316 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4230
timestamp 1682952543
transform 1 0 340 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4159
timestamp 1682952543
transform 1 0 316 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4160
timestamp 1682952543
transform 1 0 332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4161
timestamp 1682952543
transform 1 0 340 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1682952543
transform 1 0 348 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1682952543
transform 1 0 324 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4231
timestamp 1682952543
transform 1 0 380 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4163
timestamp 1682952543
transform 1 0 380 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4295
timestamp 1682952543
transform 1 0 380 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4232
timestamp 1682952543
transform 1 0 420 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4164
timestamp 1682952543
transform 1 0 404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4165
timestamp 1682952543
transform 1 0 420 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4284
timestamp 1682952543
transform 1 0 388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4285
timestamp 1682952543
transform 1 0 396 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4332
timestamp 1682952543
transform 1 0 388 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1682952543
transform 1 0 404 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4286
timestamp 1682952543
transform 1 0 428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4166
timestamp 1682952543
transform 1 0 436 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4334
timestamp 1682952543
transform 1 0 428 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4144
timestamp 1682952543
transform 1 0 460 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1682952543
transform 1 0 452 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4167
timestamp 1682952543
transform 1 0 460 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4275
timestamp 1682952543
transform 1 0 468 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4168
timestamp 1682952543
transform 1 0 476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4169
timestamp 1682952543
transform 1 0 492 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4287
timestamp 1682952543
transform 1 0 452 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4288
timestamp 1682952543
transform 1 0 460 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1682952543
transform 1 0 484 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4335
timestamp 1682952543
transform 1 0 460 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4346
timestamp 1682952543
transform 1 0 460 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4296
timestamp 1682952543
transform 1 0 492 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4170
timestamp 1682952543
transform 1 0 508 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4276
timestamp 1682952543
transform 1 0 548 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4171
timestamp 1682952543
transform 1 0 556 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4290
timestamp 1682952543
transform 1 0 548 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4336
timestamp 1682952543
transform 1 0 556 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1682952543
transform 1 0 580 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4291
timestamp 1682952543
transform 1 0 580 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4185
timestamp 1682952543
transform 1 0 596 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4172
timestamp 1682952543
transform 1 0 596 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4186
timestamp 1682952543
transform 1 0 620 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4292
timestamp 1682952543
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4145
timestamp 1682952543
transform 1 0 660 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1682952543
transform 1 0 652 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4173
timestamp 1682952543
transform 1 0 636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4174
timestamp 1682952543
transform 1 0 652 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4297
timestamp 1682952543
transform 1 0 652 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1682952543
transform 1 0 644 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4146
timestamp 1682952543
transform 1 0 676 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4175
timestamp 1682952543
transform 1 0 668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1682952543
transform 1 0 676 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4348
timestamp 1682952543
transform 1 0 668 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1682952543
transform 1 0 684 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4176
timestamp 1682952543
transform 1 0 708 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4188
timestamp 1682952543
transform 1 0 732 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4177
timestamp 1682952543
transform 1 0 724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4294
timestamp 1682952543
transform 1 0 716 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4349
timestamp 1682952543
transform 1 0 724 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4350
timestamp 1682952543
transform 1 0 740 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1682952543
transform 1 0 756 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4178
timestamp 1682952543
transform 1 0 764 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4179
timestamp 1682952543
transform 1 0 772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1682952543
transform 1 0 756 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4299
timestamp 1682952543
transform 1 0 772 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4180
timestamp 1682952543
transform 1 0 828 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4181
timestamp 1682952543
transform 1 0 876 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1682952543
transform 1 0 796 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4300
timestamp 1682952543
transform 1 0 828 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1682952543
transform 1 0 828 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1682952543
transform 1 0 884 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1682952543
transform 1 0 884 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4365
timestamp 1682952543
transform 1 0 884 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4352
timestamp 1682952543
transform 1 0 884 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4278
timestamp 1682952543
transform 1 0 900 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4353
timestamp 1682952543
transform 1 0 900 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4182
timestamp 1682952543
transform 1 0 924 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4190
timestamp 1682952543
transform 1 0 948 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4183
timestamp 1682952543
transform 1 0 980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1682952543
transform 1 0 996 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4302
timestamp 1682952543
transform 1 0 964 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4297
timestamp 1682952543
transform 1 0 972 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4298
timestamp 1682952543
transform 1 0 1004 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4303
timestamp 1682952543
transform 1 0 1028 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4185
timestamp 1682952543
transform 1 0 1060 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4279
timestamp 1682952543
transform 1 0 1068 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4299
timestamp 1682952543
transform 1 0 1068 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4191
timestamp 1682952543
transform 1 0 1084 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1682952543
transform 1 0 1116 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4233
timestamp 1682952543
transform 1 0 1108 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4186
timestamp 1682952543
transform 1 0 1092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4187
timestamp 1682952543
transform 1 0 1108 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4234
timestamp 1682952543
transform 1 0 1132 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4188
timestamp 1682952543
transform 1 0 1124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1682952543
transform 1 0 1116 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4280
timestamp 1682952543
transform 1 0 1140 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4301
timestamp 1682952543
transform 1 0 1140 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4281
timestamp 1682952543
transform 1 0 1156 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4165
timestamp 1682952543
transform 1 0 1220 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1682952543
transform 1 0 1228 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4366
timestamp 1682952543
transform 1 0 1220 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4304
timestamp 1682952543
transform 1 0 1236 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4138
timestamp 1682952543
transform 1 0 1260 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4282
timestamp 1682952543
transform 1 0 1268 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4302
timestamp 1682952543
transform 1 0 1268 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4236
timestamp 1682952543
transform 1 0 1284 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4189
timestamp 1682952543
transform 1 0 1284 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4147
timestamp 1682952543
transform 1 0 1300 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4303
timestamp 1682952543
transform 1 0 1292 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1682952543
transform 1 0 1300 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4237
timestamp 1682952543
transform 1 0 1340 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4193
timestamp 1682952543
transform 1 0 1404 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4190
timestamp 1682952543
transform 1 0 1332 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4191
timestamp 1682952543
transform 1 0 1356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4192
timestamp 1682952543
transform 1 0 1364 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4305
timestamp 1682952543
transform 1 0 1332 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1682952543
transform 1 0 1356 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1682952543
transform 1 0 1380 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4193
timestamp 1682952543
transform 1 0 1388 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1682952543
transform 1 0 1412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1682952543
transform 1 0 1380 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1682952543
transform 1 0 1404 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4148
timestamp 1682952543
transform 1 0 1436 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4307
timestamp 1682952543
transform 1 0 1428 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1682952543
transform 1 0 1444 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4149
timestamp 1682952543
transform 1 0 1508 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4166
timestamp 1682952543
transform 1 0 1476 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1682952543
transform 1 0 1524 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4150
timestamp 1682952543
transform 1 0 1580 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1682952543
transform 1 0 1532 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4239
timestamp 1682952543
transform 1 0 1572 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4195
timestamp 1682952543
transform 1 0 1468 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4196
timestamp 1682952543
transform 1 0 1476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1682952543
transform 1 0 1532 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1682952543
transform 1 0 1572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1682952543
transform 1 0 1556 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4354
timestamp 1682952543
transform 1 0 1508 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1682952543
transform 1 0 1540 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1682952543
transform 1 0 1588 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4310
timestamp 1682952543
transform 1 0 1588 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4168
timestamp 1682952543
transform 1 0 1628 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4241
timestamp 1682952543
transform 1 0 1620 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4242
timestamp 1682952543
transform 1 0 1636 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4199
timestamp 1682952543
transform 1 0 1604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4200
timestamp 1682952543
transform 1 0 1620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1682952543
transform 1 0 1636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4311
timestamp 1682952543
transform 1 0 1596 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1682952543
transform 1 0 1628 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4356
timestamp 1682952543
transform 1 0 1644 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4202
timestamp 1682952543
transform 1 0 1668 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4307
timestamp 1682952543
transform 1 0 1660 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4151
timestamp 1682952543
transform 1 0 1684 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1682952543
transform 1 0 1684 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4203
timestamp 1682952543
transform 1 0 1684 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1682952543
transform 1 0 1692 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4152
timestamp 1682952543
transform 1 0 1740 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1682952543
transform 1 0 1716 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1682952543
transform 1 0 1716 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1682952543
transform 1 0 1732 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4204
timestamp 1682952543
transform 1 0 1716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4205
timestamp 1682952543
transform 1 0 1732 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1682952543
transform 1 0 1740 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4314
timestamp 1682952543
transform 1 0 1708 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4315
timestamp 1682952543
transform 1 0 1724 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4316
timestamp 1682952543
transform 1 0 1732 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4357
timestamp 1682952543
transform 1 0 1700 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1682952543
transform 1 0 1772 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1682952543
transform 1 0 1772 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4207
timestamp 1682952543
transform 1 0 1764 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4284
timestamp 1682952543
transform 1 0 1772 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4208
timestamp 1682952543
transform 1 0 1780 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1682952543
transform 1 0 1756 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1682952543
transform 1 0 1772 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4319
timestamp 1682952543
transform 1 0 1780 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4358
timestamp 1682952543
transform 1 0 1748 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4246
timestamp 1682952543
transform 1 0 1796 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4209
timestamp 1682952543
transform 1 0 1796 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4209
timestamp 1682952543
transform 1 0 1812 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4320
timestamp 1682952543
transform 1 0 1812 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4247
timestamp 1682952543
transform 1 0 1836 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4210
timestamp 1682952543
transform 1 0 1836 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1682952543
transform 1 0 1852 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4337
timestamp 1682952543
transform 1 0 1852 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4211
timestamp 1682952543
transform 1 0 1868 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4322
timestamp 1682952543
transform 1 0 1868 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4154
timestamp 1682952543
transform 1 0 1908 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1682952543
transform 1 0 1900 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4212
timestamp 1682952543
transform 1 0 1884 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4213
timestamp 1682952543
transform 1 0 1900 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1682952543
transform 1 0 1916 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4338
timestamp 1682952543
transform 1 0 1876 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4323
timestamp 1682952543
transform 1 0 1892 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4308
timestamp 1682952543
transform 1 0 1908 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4324
timestamp 1682952543
transform 1 0 1924 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4194
timestamp 1682952543
transform 1 0 1940 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4249
timestamp 1682952543
transform 1 0 1932 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4325
timestamp 1682952543
transform 1 0 1932 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4339
timestamp 1682952543
transform 1 0 1924 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4367
timestamp 1682952543
transform 1 0 1932 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4155
timestamp 1682952543
transform 1 0 1956 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4195
timestamp 1682952543
transform 1 0 1972 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4215
timestamp 1682952543
transform 1 0 1964 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4171
timestamp 1682952543
transform 1 0 2004 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1682952543
transform 1 0 2028 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1682952543
transform 1 0 2012 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4139
timestamp 1682952543
transform 1 0 2004 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1682952543
transform 1 0 2020 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4216
timestamp 1682952543
transform 1 0 2020 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4136
timestamp 1682952543
transform 1 0 2060 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4326
timestamp 1682952543
transform 1 0 2052 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4327
timestamp 1682952543
transform 1 0 2068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4141
timestamp 1682952543
transform 1 0 2092 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4142
timestamp 1682952543
transform 1 0 2108 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4340
timestamp 1682952543
transform 1 0 2100 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1682952543
transform 1 0 2148 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4197
timestamp 1682952543
transform 1 0 2140 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4198
timestamp 1682952543
transform 1 0 2164 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4217
timestamp 1682952543
transform 1 0 2140 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4218
timestamp 1682952543
transform 1 0 2156 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4328
timestamp 1682952543
transform 1 0 2116 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1682952543
transform 1 0 2124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1682952543
transform 1 0 2108 0 1 2385
box -2 -2 2 2
use M3_M2  M3_M2_4309
timestamp 1682952543
transform 1 0 2132 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4377
timestamp 1682952543
transform 1 0 2124 0 1 2385
box -2 -2 2 2
use M3_M2  M3_M2_4199
timestamp 1682952543
transform 1 0 2180 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4219
timestamp 1682952543
transform 1 0 2188 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4330
timestamp 1682952543
transform 1 0 2188 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4250
timestamp 1682952543
transform 1 0 2220 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4173
timestamp 1682952543
transform 1 0 2308 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1682952543
transform 1 0 2292 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4251
timestamp 1682952543
transform 1 0 2260 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4220
timestamp 1682952543
transform 1 0 2260 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4310
timestamp 1682952543
transform 1 0 2260 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4311
timestamp 1682952543
transform 1 0 2276 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4272
timestamp 1682952543
transform 1 0 2308 0 1 2407
box -2 -2 2 2
use M2_M1  M2_M1_4331
timestamp 1682952543
transform 1 0 2332 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4252
timestamp 1682952543
transform 1 0 2356 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4174
timestamp 1682952543
transform 1 0 2428 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4253
timestamp 1682952543
transform 1 0 2404 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4221
timestamp 1682952543
transform 1 0 2356 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1682952543
transform 1 0 2364 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1682952543
transform 1 0 2404 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4312
timestamp 1682952543
transform 1 0 2356 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1682952543
transform 1 0 2380 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4332
timestamp 1682952543
transform 1 0 2444 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4175
timestamp 1682952543
transform 1 0 2460 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4176
timestamp 1682952543
transform 1 0 2516 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1682952543
transform 1 0 2468 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1682952543
transform 1 0 2540 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4224
timestamp 1682952543
transform 1 0 2500 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1682952543
transform 1 0 2476 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4368
timestamp 1682952543
transform 1 0 2580 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4177
timestamp 1682952543
transform 1 0 2628 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1682952543
transform 1 0 2604 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1682952543
transform 1 0 2620 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4134
timestamp 1682952543
transform 1 0 2644 0 1 2445
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1682952543
transform 1 0 2604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4226
timestamp 1682952543
transform 1 0 2620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1682952543
transform 1 0 2628 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1682952543
transform 1 0 2636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4334
timestamp 1682952543
transform 1 0 2612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4255
timestamp 1682952543
transform 1 0 2668 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4135
timestamp 1682952543
transform 1 0 2684 0 1 2445
box -2 -2 2 2
use M3_M2  M3_M2_4211
timestamp 1682952543
transform 1 0 2684 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1682952543
transform 1 0 2724 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1682952543
transform 1 0 2708 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4229
timestamp 1682952543
transform 1 0 2708 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1682952543
transform 1 0 2724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1682952543
transform 1 0 2716 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4314
timestamp 1682952543
transform 1 0 2724 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4315
timestamp 1682952543
transform 1 0 2748 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1682952543
transform 1 0 2764 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4157
timestamp 1682952543
transform 1 0 2852 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4231
timestamp 1682952543
transform 1 0 2788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1682952543
transform 1 0 2836 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4213
timestamp 1682952543
transform 1 0 2916 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1682952543
transform 1 0 3004 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1682952543
transform 1 0 2964 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4233
timestamp 1682952543
transform 1 0 2900 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1682952543
transform 1 0 2908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1682952543
transform 1 0 2964 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4285
timestamp 1682952543
transform 1 0 2988 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4178
timestamp 1682952543
transform 1 0 3044 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4143
timestamp 1682952543
transform 1 0 3020 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4236
timestamp 1682952543
transform 1 0 3004 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4336
timestamp 1682952543
transform 1 0 2868 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1682952543
transform 1 0 2884 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4316
timestamp 1682952543
transform 1 0 2892 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4317
timestamp 1682952543
transform 1 0 2908 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4338
timestamp 1682952543
transform 1 0 2988 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4359
timestamp 1682952543
transform 1 0 2956 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1682952543
transform 1 0 3028 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1682952543
transform 1 0 3052 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4158
timestamp 1682952543
transform 1 0 3100 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1682952543
transform 1 0 3076 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4237
timestamp 1682952543
transform 1 0 3044 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1682952543
transform 1 0 3060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1682952543
transform 1 0 3028 0 1 2407
box -2 -2 2 2
use M3_M2  M3_M2_4318
timestamp 1682952543
transform 1 0 3036 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1682952543
transform 1 0 3068 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4179
timestamp 1682952543
transform 1 0 3124 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1682952543
transform 1 0 3116 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4239
timestamp 1682952543
transform 1 0 3076 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4287
timestamp 1682952543
transform 1 0 3092 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4240
timestamp 1682952543
transform 1 0 3108 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1682952543
transform 1 0 3124 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1682952543
transform 1 0 3052 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1682952543
transform 1 0 3068 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4319
timestamp 1682952543
transform 1 0 3076 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4341
timestamp 1682952543
transform 1 0 3100 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4369
timestamp 1682952543
transform 1 0 3076 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1682952543
transform 1 0 3084 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4360
timestamp 1682952543
transform 1 0 3068 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4320
timestamp 1682952543
transform 1 0 3108 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4342
timestamp 1682952543
transform 1 0 3116 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4361
timestamp 1682952543
transform 1 0 3100 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4159
timestamp 1682952543
transform 1 0 3220 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4216
timestamp 1682952543
transform 1 0 3204 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4144
timestamp 1682952543
transform 1 0 3164 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4261
timestamp 1682952543
transform 1 0 3196 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4262
timestamp 1682952543
transform 1 0 3228 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4217
timestamp 1682952543
transform 1 0 3284 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4218
timestamp 1682952543
transform 1 0 3308 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4263
timestamp 1682952543
transform 1 0 3372 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4242
timestamp 1682952543
transform 1 0 3196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4243
timestamp 1682952543
transform 1 0 3220 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4244
timestamp 1682952543
transform 1 0 3236 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4343
timestamp 1682952543
transform 1 0 3140 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4344
timestamp 1682952543
transform 1 0 3148 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1682952543
transform 1 0 3164 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4362
timestamp 1682952543
transform 1 0 3164 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4288
timestamp 1682952543
transform 1 0 3252 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4245
timestamp 1682952543
transform 1 0 3260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4246
timestamp 1682952543
transform 1 0 3268 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1682952543
transform 1 0 3276 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4289
timestamp 1682952543
transform 1 0 3308 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4160
timestamp 1682952543
transform 1 0 3540 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4204
timestamp 1682952543
transform 1 0 3420 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4205
timestamp 1682952543
transform 1 0 3540 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4219
timestamp 1682952543
transform 1 0 3444 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4220
timestamp 1682952543
transform 1 0 3476 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4180
timestamp 1682952543
transform 1 0 3580 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4137
timestamp 1682952543
transform 1 0 3540 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_4221
timestamp 1682952543
transform 1 0 3556 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4264
timestamp 1682952543
transform 1 0 3436 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1682952543
transform 1 0 3540 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4145
timestamp 1682952543
transform 1 0 3556 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1682952543
transform 1 0 3380 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1682952543
transform 1 0 3396 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4250
timestamp 1682952543
transform 1 0 3412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4251
timestamp 1682952543
transform 1 0 3420 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4252
timestamp 1682952543
transform 1 0 3428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1682952543
transform 1 0 3436 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4346
timestamp 1682952543
transform 1 0 3228 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4363
timestamp 1682952543
transform 1 0 3220 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4274
timestamp 1682952543
transform 1 0 3260 0 1 2407
box -2 -2 2 2
use M3_M2  M3_M2_4321
timestamp 1682952543
transform 1 0 3364 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4347
timestamp 1682952543
transform 1 0 3372 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4322
timestamp 1682952543
transform 1 0 3380 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4348
timestamp 1682952543
transform 1 0 3388 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4349
timestamp 1682952543
transform 1 0 3404 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1682952543
transform 1 0 3364 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4290
timestamp 1682952543
transform 1 0 3460 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4291
timestamp 1682952543
transform 1 0 3524 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1682952543
transform 1 0 3476 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4292
timestamp 1682952543
transform 1 0 3556 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4222
timestamp 1682952543
transform 1 0 3588 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4223
timestamp 1682952543
transform 1 0 3604 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4254
timestamp 1682952543
transform 1 0 3580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1682952543
transform 1 0 3532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1682952543
transform 1 0 3524 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4364
timestamp 1682952543
transform 1 0 3532 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4275
timestamp 1682952543
transform 1 0 3564 0 1 2407
box -2 -2 2 2
use M2_M1  M2_M1_4146
timestamp 1682952543
transform 1 0 3612 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4181
timestamp 1682952543
transform 1 0 3636 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1682952543
transform 1 0 3612 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4161
timestamp 1682952543
transform 1 0 3660 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1682952543
transform 1 0 3644 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4255
timestamp 1682952543
transform 1 0 3636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4256
timestamp 1682952543
transform 1 0 3652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4351
timestamp 1682952543
transform 1 0 3588 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4352
timestamp 1682952543
transform 1 0 3596 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4365
timestamp 1682952543
transform 1 0 3596 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4353
timestamp 1682952543
transform 1 0 3620 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4267
timestamp 1682952543
transform 1 0 3676 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4257
timestamp 1682952543
transform 1 0 3676 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1682952543
transform 1 0 3684 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1682952543
transform 1 0 3644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4355
timestamp 1682952543
transform 1 0 3660 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1682952543
transform 1 0 3676 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4182
timestamp 1682952543
transform 1 0 3812 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4224
timestamp 1682952543
transform 1 0 3708 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1682952543
transform 1 0 3788 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4147
timestamp 1682952543
transform 1 0 3796 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4259
timestamp 1682952543
transform 1 0 3692 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1682952543
transform 1 0 3756 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4261
timestamp 1682952543
transform 1 0 3788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4276
timestamp 1682952543
transform 1 0 3708 0 1 2407
box -2 -2 2 2
use M2_M1  M2_M1_4148
timestamp 1682952543
transform 1 0 3828 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1682952543
transform 1 0 3812 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1682952543
transform 1 0 3828 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4324
timestamp 1682952543
transform 1 0 3788 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4356
timestamp 1682952543
transform 1 0 3796 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4341
timestamp 1682952543
transform 1 0 3740 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1682952543
transform 1 0 3756 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4343
timestamp 1682952543
transform 1 0 3796 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4357
timestamp 1682952543
transform 1 0 3820 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4325
timestamp 1682952543
transform 1 0 3828 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4344
timestamp 1682952543
transform 1 0 3828 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4162
timestamp 1682952543
transform 1 0 3908 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4268
timestamp 1682952543
transform 1 0 3884 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4264
timestamp 1682952543
transform 1 0 3844 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1682952543
transform 1 0 3868 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4294
timestamp 1682952543
transform 1 0 3876 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4266
timestamp 1682952543
transform 1 0 3884 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4226
timestamp 1682952543
transform 1 0 3924 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4358
timestamp 1682952543
transform 1 0 3844 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4359
timestamp 1682952543
transform 1 0 3852 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4360
timestamp 1682952543
transform 1 0 3876 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1682952543
transform 1 0 3884 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4326
timestamp 1682952543
transform 1 0 3892 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4362
timestamp 1682952543
transform 1 0 3908 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4327
timestamp 1682952543
transform 1 0 3916 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4267
timestamp 1682952543
transform 1 0 3932 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4363
timestamp 1682952543
transform 1 0 3924 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4345
timestamp 1682952543
transform 1 0 3884 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4374
timestamp 1682952543
transform 1 0 3892 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4366
timestamp 1682952543
transform 1 0 3876 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4367
timestamp 1682952543
transform 1 0 3900 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4163
timestamp 1682952543
transform 1 0 4044 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1682952543
transform 1 0 4060 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4268
timestamp 1682952543
transform 1 0 3948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1682952543
transform 1 0 3956 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1682952543
transform 1 0 4060 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4271
timestamp 1682952543
transform 1 0 4100 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4328
timestamp 1682952543
transform 1 0 3996 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4375
timestamp 1682952543
transform 1 0 4044 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4364
timestamp 1682952543
transform 1 0 4140 0 1 2405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_34
timestamp 1682952543
transform 1 0 48 0 1 2370
box -10 -3 10 3
use FILL  FILL_1236
timestamp 1682952543
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1682952543
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_1238
timestamp 1682952543
transform 1 0 88 0 1 2370
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1682952543
transform 1 0 96 0 1 2370
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1682952543
transform 1 0 104 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_301
timestamp 1682952543
transform -1 0 128 0 1 2370
box -9 -3 26 105
use INVX2  INVX2_302
timestamp 1682952543
transform -1 0 144 0 1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_154
timestamp 1682952543
transform -1 0 184 0 1 2370
box -8 -3 46 105
use FILL  FILL_1241
timestamp 1682952543
transform 1 0 184 0 1 2370
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1682952543
transform 1 0 192 0 1 2370
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1682952543
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1682952543
transform 1 0 208 0 1 2370
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1682952543
transform 1 0 216 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_303
timestamp 1682952543
transform -1 0 240 0 1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_155
timestamp 1682952543
transform 1 0 240 0 1 2370
box -8 -3 46 105
use FILL  FILL_1248
timestamp 1682952543
transform 1 0 280 0 1 2370
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1682952543
transform 1 0 288 0 1 2370
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1682952543
transform 1 0 296 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4368
timestamp 1682952543
transform 1 0 340 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_197
timestamp 1682952543
transform -1 0 344 0 1 2370
box -8 -3 46 105
use FILL  FILL_1251
timestamp 1682952543
transform 1 0 344 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_305
timestamp 1682952543
transform -1 0 368 0 1 2370
box -9 -3 26 105
use FILL  FILL_1252
timestamp 1682952543
transform 1 0 368 0 1 2370
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1682952543
transform 1 0 376 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_158
timestamp 1682952543
transform -1 0 424 0 1 2370
box -8 -3 46 105
use FILL  FILL_1254
timestamp 1682952543
transform 1 0 424 0 1 2370
box -8 -3 16 105
use FILL  FILL_1255
timestamp 1682952543
transform 1 0 432 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_306
timestamp 1682952543
transform -1 0 456 0 1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_159
timestamp 1682952543
transform 1 0 456 0 1 2370
box -8 -3 46 105
use FILL  FILL_1256
timestamp 1682952543
transform 1 0 496 0 1 2370
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1682952543
transform 1 0 504 0 1 2370
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1682952543
transform 1 0 512 0 1 2370
box -8 -3 16 105
use FILL  FILL_1259
timestamp 1682952543
transform 1 0 520 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_198
timestamp 1682952543
transform 1 0 528 0 1 2370
box -8 -3 46 105
use FILL  FILL_1260
timestamp 1682952543
transform 1 0 568 0 1 2370
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1682952543
transform 1 0 576 0 1 2370
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1682952543
transform 1 0 584 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_43
timestamp 1682952543
transform 1 0 592 0 1 2370
box -5 -3 28 105
use FILL  FILL_1263
timestamp 1682952543
transform 1 0 616 0 1 2370
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1682952543
transform 1 0 624 0 1 2370
box -8 -3 16 105
use AND2X2  AND2X2_40
timestamp 1682952543
transform -1 0 664 0 1 2370
box -8 -3 40 105
use FILL  FILL_1265
timestamp 1682952543
transform 1 0 664 0 1 2370
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1682952543
transform 1 0 672 0 1 2370
box -8 -3 16 105
use FILL  FILL_1267
timestamp 1682952543
transform 1 0 680 0 1 2370
box -8 -3 16 105
use AND2X2  AND2X2_41
timestamp 1682952543
transform -1 0 720 0 1 2370
box -8 -3 40 105
use FILL  FILL_1268
timestamp 1682952543
transform 1 0 720 0 1 2370
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1682952543
transform 1 0 728 0 1 2370
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1682952543
transform 1 0 736 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4369
timestamp 1682952543
transform 1 0 756 0 1 2375
box -3 -3 3 3
use FILL  FILL_1271
timestamp 1682952543
transform 1 0 744 0 1 2370
box -8 -3 16 105
use FILL  FILL_1278
timestamp 1682952543
transform 1 0 752 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4370
timestamp 1682952543
transform 1 0 772 0 1 2375
box -3 -3 3 3
use INVX2  INVX2_310
timestamp 1682952543
transform 1 0 760 0 1 2370
box -9 -3 26 105
use FILL  FILL_1280
timestamp 1682952543
transform 1 0 776 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4371
timestamp 1682952543
transform 1 0 796 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4372
timestamp 1682952543
transform 1 0 812 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4373
timestamp 1682952543
transform 1 0 868 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_270
timestamp 1682952543
transform 1 0 784 0 1 2370
box -8 -3 104 105
use FILL  FILL_1284
timestamp 1682952543
transform 1 0 880 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_54
timestamp 1682952543
transform 1 0 888 0 1 2370
box -8 -3 32 105
use FILL  FILL_1293
timestamp 1682952543
transform 1 0 912 0 1 2370
box -8 -3 16 105
use FILL  FILL_1294
timestamp 1682952543
transform 1 0 920 0 1 2370
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1682952543
transform 1 0 928 0 1 2370
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1682952543
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1682952543
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1682952543
transform 1 0 952 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_164
timestamp 1682952543
transform 1 0 960 0 1 2370
box -8 -3 46 105
use FILL  FILL_1304
timestamp 1682952543
transform 1 0 1000 0 1 2370
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1682952543
transform 1 0 1008 0 1 2370
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1682952543
transform 1 0 1016 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4374
timestamp 1682952543
transform 1 0 1036 0 1 2375
box -3 -3 3 3
use FILL  FILL_1312
timestamp 1682952543
transform 1 0 1024 0 1 2370
box -8 -3 16 105
use FILL  FILL_1314
timestamp 1682952543
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use FILL  FILL_1316
timestamp 1682952543
transform 1 0 1040 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4375
timestamp 1682952543
transform 1 0 1068 0 1 2375
box -3 -3 3 3
use FILL  FILL_1318
timestamp 1682952543
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1682952543
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1682952543
transform 1 0 1064 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_165
timestamp 1682952543
transform -1 0 1112 0 1 2370
box -8 -3 46 105
use M3_M2  M3_M2_4376
timestamp 1682952543
transform 1 0 1124 0 1 2375
box -3 -3 3 3
use FILL  FILL_1323
timestamp 1682952543
transform 1 0 1112 0 1 2370
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1682952543
transform 1 0 1120 0 1 2370
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1682952543
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1682952543
transform 1 0 1136 0 1 2370
box -8 -3 16 105
use FILL  FILL_1333
timestamp 1682952543
transform 1 0 1144 0 1 2370
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1682952543
transform 1 0 1152 0 1 2370
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1682952543
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1682952543
transform 1 0 1168 0 1 2370
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1682952543
transform 1 0 1176 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_56
timestamp 1682952543
transform 1 0 1184 0 1 2370
box -8 -3 34 105
use FILL  FILL_1340
timestamp 1682952543
transform 1 0 1216 0 1 2370
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1682952543
transform 1 0 1224 0 1 2370
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1682952543
transform 1 0 1232 0 1 2370
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1682952543
transform 1 0 1240 0 1 2370
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1682952543
transform 1 0 1248 0 1 2370
box -8 -3 16 105
use FILL  FILL_1353
timestamp 1682952543
transform 1 0 1256 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_56
timestamp 1682952543
transform 1 0 1264 0 1 2370
box -8 -3 32 105
use FILL  FILL_1355
timestamp 1682952543
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1682952543
transform 1 0 1296 0 1 2370
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1682952543
transform 1 0 1304 0 1 2370
box -8 -3 16 105
use FILL  FILL_1358
timestamp 1682952543
transform 1 0 1312 0 1 2370
box -8 -3 16 105
use AND2X2  AND2X2_42
timestamp 1682952543
transform 1 0 1320 0 1 2370
box -8 -3 40 105
use FILL  FILL_1362
timestamp 1682952543
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_45
timestamp 1682952543
transform 1 0 1360 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_46
timestamp 1682952543
transform 1 0 1384 0 1 2370
box -5 -3 28 105
use M3_M2  M3_M2_4377
timestamp 1682952543
transform 1 0 1428 0 1 2375
box -3 -3 3 3
use BUFX2  BUFX2_47
timestamp 1682952543
transform 1 0 1408 0 1 2370
box -5 -3 28 105
use FILL  FILL_1372
timestamp 1682952543
transform 1 0 1432 0 1 2370
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1682952543
transform 1 0 1440 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_49
timestamp 1682952543
transform -1 0 1472 0 1 2370
box -5 -3 28 105
use M3_M2  M3_M2_4378
timestamp 1682952543
transform 1 0 1508 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_271
timestamp 1682952543
transform -1 0 1568 0 1 2370
box -8 -3 104 105
use INVX2  INVX2_312
timestamp 1682952543
transform -1 0 1584 0 1 2370
box -9 -3 26 105
use FILL  FILL_1374
timestamp 1682952543
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_1375
timestamp 1682952543
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_166
timestamp 1682952543
transform 1 0 1600 0 1 2370
box -8 -3 46 105
use FILL  FILL_1376
timestamp 1682952543
transform 1 0 1640 0 1 2370
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1682952543
transform 1 0 1648 0 1 2370
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1682952543
transform 1 0 1656 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_313
timestamp 1682952543
transform -1 0 1680 0 1 2370
box -9 -3 26 105
use FILL  FILL_1379
timestamp 1682952543
transform 1 0 1680 0 1 2370
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1682952543
transform 1 0 1688 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4379
timestamp 1682952543
transform 1 0 1724 0 1 2375
box -3 -3 3 3
use AOI22X1  AOI22X1_167
timestamp 1682952543
transform -1 0 1736 0 1 2370
box -8 -3 46 105
use FILL  FILL_1381
timestamp 1682952543
transform 1 0 1736 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4380
timestamp 1682952543
transform 1 0 1772 0 1 2375
box -3 -3 3 3
use AOI22X1  AOI22X1_168
timestamp 1682952543
transform -1 0 1784 0 1 2370
box -8 -3 46 105
use FILL  FILL_1382
timestamp 1682952543
transform 1 0 1784 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_50
timestamp 1682952543
transform 1 0 1792 0 1 2370
box -5 -3 28 105
use FILL  FILL_1383
timestamp 1682952543
transform 1 0 1816 0 1 2370
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1682952543
transform 1 0 1824 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_51
timestamp 1682952543
transform 1 0 1832 0 1 2370
box -5 -3 28 105
use M3_M2  M3_M2_4381
timestamp 1682952543
transform 1 0 1868 0 1 2375
box -3 -3 3 3
use FILL  FILL_1385
timestamp 1682952543
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_1401
timestamp 1682952543
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4382
timestamp 1682952543
transform 1 0 1884 0 1 2375
box -3 -3 3 3
use FILL  FILL_1403
timestamp 1682952543
transform 1 0 1872 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4383
timestamp 1682952543
transform 1 0 1916 0 1 2375
box -3 -3 3 3
use AOI22X1  AOI22X1_170
timestamp 1682952543
transform 1 0 1880 0 1 2370
box -8 -3 46 105
use FILL  FILL_1404
timestamp 1682952543
transform 1 0 1920 0 1 2370
box -8 -3 16 105
use FILL  FILL_1407
timestamp 1682952543
transform 1 0 1928 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_316
timestamp 1682952543
transform 1 0 1936 0 1 2370
box -9 -3 26 105
use FILL  FILL_1409
timestamp 1682952543
transform 1 0 1952 0 1 2370
box -8 -3 16 105
use FILL  FILL_1410
timestamp 1682952543
transform 1 0 1960 0 1 2370
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1682952543
transform 1 0 1968 0 1 2370
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1682952543
transform 1 0 1976 0 1 2370
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1682952543
transform 1 0 1984 0 1 2370
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1682952543
transform 1 0 1992 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4384
timestamp 1682952543
transform 1 0 2028 0 1 2375
box -3 -3 3 3
use NAND3X1  NAND3X1_25
timestamp 1682952543
transform -1 0 2032 0 1 2370
box -8 -3 40 105
use FILL  FILL_1415
timestamp 1682952543
transform 1 0 2032 0 1 2370
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1682952543
transform 1 0 2040 0 1 2370
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1682952543
transform 1 0 2048 0 1 2370
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1682952543
transform 1 0 2056 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_54
timestamp 1682952543
transform -1 0 2088 0 1 2370
box -5 -3 28 105
use FILL  FILL_1419
timestamp 1682952543
transform 1 0 2088 0 1 2370
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1682952543
transform 1 0 2096 0 1 2370
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1682952543
transform 1 0 2104 0 1 2370
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1682952543
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4385
timestamp 1682952543
transform 1 0 2132 0 1 2375
box -3 -3 3 3
use FILL  FILL_1423
timestamp 1682952543
transform 1 0 2120 0 1 2370
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1682952543
transform 1 0 2128 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_172
timestamp 1682952543
transform 1 0 2136 0 1 2370
box -8 -3 46 105
use FILL  FILL_1425
timestamp 1682952543
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1682952543
transform 1 0 2184 0 1 2370
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1682952543
transform 1 0 2192 0 1 2370
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1682952543
transform 1 0 2200 0 1 2370
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1682952543
transform 1 0 2208 0 1 2370
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1682952543
transform 1 0 2216 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_275
timestamp 1682952543
transform -1 0 2320 0 1 2370
box -8 -3 104 105
use M3_M2  M3_M2_4386
timestamp 1682952543
transform 1 0 2332 0 1 2375
box -3 -3 3 3
use FILL  FILL_1442
timestamp 1682952543
transform 1 0 2320 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_318
timestamp 1682952543
transform 1 0 2328 0 1 2370
box -9 -3 26 105
use FILL  FILL_1446
timestamp 1682952543
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1682952543
transform 1 0 2352 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4387
timestamp 1682952543
transform 1 0 2396 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4388
timestamp 1682952543
transform 1 0 2444 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_277
timestamp 1682952543
transform -1 0 2456 0 1 2370
box -8 -3 104 105
use FILL  FILL_1448
timestamp 1682952543
transform 1 0 2456 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4389
timestamp 1682952543
transform 1 0 2476 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_278
timestamp 1682952543
transform 1 0 2464 0 1 2370
box -8 -3 104 105
use FILL  FILL_1456
timestamp 1682952543
transform 1 0 2560 0 1 2370
box -8 -3 16 105
use FILL  FILL_1457
timestamp 1682952543
transform 1 0 2568 0 1 2370
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1682952543
transform 1 0 2576 0 1 2370
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1682952543
transform 1 0 2584 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_201
timestamp 1682952543
transform -1 0 2632 0 1 2370
box -8 -3 46 105
use FILL  FILL_1460
timestamp 1682952543
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_1476
timestamp 1682952543
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1682952543
transform 1 0 2648 0 1 2370
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1682952543
transform 1 0 2656 0 1 2370
box -8 -3 16 105
use FILL  FILL_1481
timestamp 1682952543
transform 1 0 2664 0 1 2370
box -8 -3 16 105
use FILL  FILL_1482
timestamp 1682952543
transform 1 0 2672 0 1 2370
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1682952543
transform 1 0 2680 0 1 2370
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1682952543
transform 1 0 2688 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_202
timestamp 1682952543
transform 1 0 2696 0 1 2370
box -8 -3 46 105
use FILL  FILL_1485
timestamp 1682952543
transform 1 0 2736 0 1 2370
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1682952543
transform 1 0 2744 0 1 2370
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1682952543
transform 1 0 2752 0 1 2370
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1682952543
transform 1 0 2760 0 1 2370
box -8 -3 16 105
use FILL  FILL_1497
timestamp 1682952543
transform 1 0 2768 0 1 2370
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1682952543
transform 1 0 2776 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4390
timestamp 1682952543
transform 1 0 2868 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_279
timestamp 1682952543
transform -1 0 2880 0 1 2370
box -8 -3 104 105
use BUFX2  BUFX2_58
timestamp 1682952543
transform -1 0 2904 0 1 2370
box -5 -3 28 105
use M3_M2  M3_M2_4391
timestamp 1682952543
transform 1 0 2940 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_280
timestamp 1682952543
transform -1 0 3000 0 1 2370
box -8 -3 104 105
use M3_M2  M3_M2_4392
timestamp 1682952543
transform 1 0 3012 0 1 2375
box -3 -3 3 3
use NAND2X1  NAND2X1_56
timestamp 1682952543
transform 1 0 3000 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_59
timestamp 1682952543
transform -1 0 3056 0 1 2370
box -8 -3 34 105
use M3_M2  M3_M2_4393
timestamp 1682952543
transform 1 0 3068 0 1 2375
box -3 -3 3 3
use NOR2X1  NOR2X1_57
timestamp 1682952543
transform -1 0 3080 0 1 2370
box -8 -3 32 105
use AOI21X1  AOI21X1_17
timestamp 1682952543
transform -1 0 3112 0 1 2370
box -7 -3 39 105
use OAI21X1  OAI21X1_60
timestamp 1682952543
transform 1 0 3112 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_57
timestamp 1682952543
transform 1 0 3144 0 1 2370
box -8 -3 32 105
use XOR2X1  XOR2X1_7
timestamp 1682952543
transform -1 0 3224 0 1 2370
box -8 -3 64 105
use AND2X2  AND2X2_43
timestamp 1682952543
transform 1 0 3224 0 1 2370
box -8 -3 40 105
use FAX1  FAX1_19
timestamp 1682952543
transform 1 0 3256 0 1 2370
box -5 -3 126 105
use AOI22X1  AOI22X1_175
timestamp 1682952543
transform 1 0 3376 0 1 2370
box -8 -3 46 105
use FAX1  FAX1_20
timestamp 1682952543
transform 1 0 3416 0 1 2370
box -5 -3 126 105
use NAND2X1  NAND2X1_58
timestamp 1682952543
transform 1 0 3536 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_61
timestamp 1682952543
transform -1 0 3592 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_59
timestamp 1682952543
transform 1 0 3592 0 1 2370
box -8 -3 32 105
use OAI21X1  OAI21X1_62
timestamp 1682952543
transform -1 0 3648 0 1 2370
box -8 -3 34 105
use AOI21X1  AOI21X1_18
timestamp 1682952543
transform 1 0 3648 0 1 2370
box -7 -3 39 105
use INVX2  INVX2_320
timestamp 1682952543
transform -1 0 3696 0 1 2370
box -9 -3 26 105
use M3_M2  M3_M2_4394
timestamp 1682952543
transform 1 0 3732 0 1 2375
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1682952543
transform 1 0 3764 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_281
timestamp 1682952543
transform 1 0 3696 0 1 2370
box -8 -3 104 105
use OAI21X1  OAI21X1_63
timestamp 1682952543
transform -1 0 3824 0 1 2370
box -8 -3 34 105
use NAND2X1  NAND2X1_60
timestamp 1682952543
transform -1 0 3848 0 1 2370
box -8 -3 32 105
use AOI22X1  AOI22X1_176
timestamp 1682952543
transform 1 0 3848 0 1 2370
box -8 -3 46 105
use AOI21X1  AOI21X1_19
timestamp 1682952543
transform -1 0 3920 0 1 2370
box -7 -3 39 105
use FILL  FILL_1499
timestamp 1682952543
transform 1 0 3920 0 1 2370
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1682952543
transform 1 0 3928 0 1 2370
box -8 -3 16 105
use FAX1  FAX1_21
timestamp 1682952543
transform 1 0 3936 0 1 2370
box -5 -3 126 105
use M3_M2  M3_M2_4396
timestamp 1682952543
transform 1 0 4092 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_282
timestamp 1682952543
transform -1 0 4152 0 1 2370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_35
timestamp 1682952543
transform 1 0 4177 0 1 2370
box -10 -3 10 3
use M3_M2  M3_M2_4397
timestamp 1682952543
transform 1 0 140 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4398
timestamp 1682952543
transform 1 0 188 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4424
timestamp 1682952543
transform 1 0 164 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4425
timestamp 1682952543
transform 1 0 180 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4384
timestamp 1682952543
transform 1 0 84 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4456
timestamp 1682952543
transform 1 0 156 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4385
timestamp 1682952543
transform 1 0 180 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1682952543
transform 1 0 196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1682952543
transform 1 0 204 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4457
timestamp 1682952543
transform 1 0 212 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4472
timestamp 1682952543
transform 1 0 108 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1682952543
transform 1 0 164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4474
timestamp 1682952543
transform 1 0 172 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1682952543
transform 1 0 188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4476
timestamp 1682952543
transform 1 0 212 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4481
timestamp 1682952543
transform 1 0 196 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4482
timestamp 1682952543
transform 1 0 220 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4426
timestamp 1682952543
transform 1 0 276 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4388
timestamp 1682952543
transform 1 0 244 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4389
timestamp 1682952543
transform 1 0 252 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4390
timestamp 1682952543
transform 1 0 268 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4391
timestamp 1682952543
transform 1 0 276 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1682952543
transform 1 0 244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4478
timestamp 1682952543
transform 1 0 260 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4483
timestamp 1682952543
transform 1 0 252 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4518
timestamp 1682952543
transform 1 0 244 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_4479
timestamp 1682952543
transform 1 0 284 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4399
timestamp 1682952543
transform 1 0 308 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4427
timestamp 1682952543
transform 1 0 324 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4428
timestamp 1682952543
transform 1 0 372 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4392
timestamp 1682952543
transform 1 0 308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4393
timestamp 1682952543
transform 1 0 324 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4458
timestamp 1682952543
transform 1 0 340 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4394
timestamp 1682952543
transform 1 0 348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4395
timestamp 1682952543
transform 1 0 356 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1682952543
transform 1 0 372 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4397
timestamp 1682952543
transform 1 0 380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4480
timestamp 1682952543
transform 1 0 300 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1682952543
transform 1 0 316 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1682952543
transform 1 0 324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4483
timestamp 1682952543
transform 1 0 340 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1682952543
transform 1 0 364 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4484
timestamp 1682952543
transform 1 0 356 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4485
timestamp 1682952543
transform 1 0 380 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4398
timestamp 1682952543
transform 1 0 412 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4459
timestamp 1682952543
transform 1 0 500 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4485
timestamp 1682952543
transform 1 0 396 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1682952543
transform 1 0 436 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1682952543
transform 1 0 492 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1682952543
transform 1 0 500 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4519
timestamp 1682952543
transform 1 0 388 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1682952543
transform 1 0 460 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4429
timestamp 1682952543
transform 1 0 612 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4399
timestamp 1682952543
transform 1 0 516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4400
timestamp 1682952543
transform 1 0 532 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4546
timestamp 1682952543
transform 1 0 508 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4489
timestamp 1682952543
transform 1 0 580 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1682952543
transform 1 0 612 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1682952543
transform 1 0 628 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4487
timestamp 1682952543
transform 1 0 580 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4547
timestamp 1682952543
transform 1 0 540 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4488
timestamp 1682952543
transform 1 0 628 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4405
timestamp 1682952543
transform 1 0 644 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4406
timestamp 1682952543
transform 1 0 668 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4430
timestamp 1682952543
transform 1 0 692 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4401
timestamp 1682952543
transform 1 0 668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1682952543
transform 1 0 676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4403
timestamp 1682952543
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4492
timestamp 1682952543
transform 1 0 660 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4489
timestamp 1682952543
transform 1 0 652 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4431
timestamp 1682952543
transform 1 0 716 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4404
timestamp 1682952543
transform 1 0 716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4493
timestamp 1682952543
transform 1 0 684 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1682952543
transform 1 0 700 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1682952543
transform 1 0 708 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1682952543
transform 1 0 724 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4497
timestamp 1682952543
transform 1 0 740 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4490
timestamp 1682952543
transform 1 0 684 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1682952543
transform 1 0 700 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4520
timestamp 1682952543
transform 1 0 676 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1682952543
transform 1 0 740 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1682952543
transform 1 0 716 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4526
timestamp 1682952543
transform 1 0 708 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4498
timestamp 1682952543
transform 1 0 756 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4527
timestamp 1682952543
transform 1 0 748 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4405
timestamp 1682952543
transform 1 0 772 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4493
timestamp 1682952543
transform 1 0 772 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4432
timestamp 1682952543
transform 1 0 788 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4406
timestamp 1682952543
transform 1 0 788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4407
timestamp 1682952543
transform 1 0 812 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4408
timestamp 1682952543
transform 1 0 820 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4499
timestamp 1682952543
transform 1 0 804 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1682952543
transform 1 0 820 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1682952543
transform 1 0 828 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4494
timestamp 1682952543
transform 1 0 828 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4522
timestamp 1682952543
transform 1 0 820 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4528
timestamp 1682952543
transform 1 0 796 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4529
timestamp 1682952543
transform 1 0 820 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4588
timestamp 1682952543
transform 1 0 836 0 1 2295
box -2 -2 2 2
use M2_M1  M2_M1_4409
timestamp 1682952543
transform 1 0 852 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4530
timestamp 1682952543
transform 1 0 852 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4589
timestamp 1682952543
transform 1 0 852 0 1 2285
box -2 -2 2 2
use M3_M2  M3_M2_4407
timestamp 1682952543
transform 1 0 868 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4410
timestamp 1682952543
transform 1 0 868 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1682952543
transform 1 0 868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1682952543
transform 1 0 876 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4531
timestamp 1682952543
transform 1 0 868 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4408
timestamp 1682952543
transform 1 0 900 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1682952543
transform 1 0 900 0 1 2335
box -3 -3 3 3
use M3_M2  M3_M2_4400
timestamp 1682952543
transform 1 0 924 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4378
timestamp 1682952543
transform 1 0 924 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4461
timestamp 1682952543
transform 1 0 924 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4411
timestamp 1682952543
transform 1 0 932 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4433
timestamp 1682952543
transform 1 0 948 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1682952543
transform 1 0 964 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4412
timestamp 1682952543
transform 1 0 956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4580
timestamp 1682952543
transform 1 0 972 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4495
timestamp 1682952543
transform 1 0 980 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4523
timestamp 1682952543
transform 1 0 972 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4532
timestamp 1682952543
transform 1 0 980 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4524
timestamp 1682952543
transform 1 0 1004 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_4413
timestamp 1682952543
transform 1 0 1036 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4402
timestamp 1682952543
transform 1 0 1060 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4434
timestamp 1682952543
transform 1 0 1060 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4403
timestamp 1682952543
transform 1 0 1076 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4504
timestamp 1682952543
transform 1 0 1060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1682952543
transform 1 0 1068 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4435
timestamp 1682952543
transform 1 0 1092 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4414
timestamp 1682952543
transform 1 0 1092 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1682952543
transform 1 0 1092 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4415
timestamp 1682952543
transform 1 0 1108 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4496
timestamp 1682952543
transform 1 0 1108 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4507
timestamp 1682952543
transform 1 0 1164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1682952543
transform 1 0 1156 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4462
timestamp 1682952543
transform 1 0 1188 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4582
timestamp 1682952543
transform 1 0 1172 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4548
timestamp 1682952543
transform 1 0 1172 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4508
timestamp 1682952543
transform 1 0 1220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1682952543
transform 1 0 1212 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4497
timestamp 1682952543
transform 1 0 1220 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4549
timestamp 1682952543
transform 1 0 1212 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4379
timestamp 1682952543
transform 1 0 1260 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_4416
timestamp 1682952543
transform 1 0 1268 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4550
timestamp 1682952543
transform 1 0 1268 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4436
timestamp 1682952543
transform 1 0 1292 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4509
timestamp 1682952543
transform 1 0 1300 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4498
timestamp 1682952543
transform 1 0 1300 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4551
timestamp 1682952543
transform 1 0 1284 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4552
timestamp 1682952543
transform 1 0 1356 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4409
timestamp 1682952543
transform 1 0 1372 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4437
timestamp 1682952543
transform 1 0 1364 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4417
timestamp 1682952543
transform 1 0 1364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4510
timestamp 1682952543
transform 1 0 1372 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4467
timestamp 1682952543
transform 1 0 1380 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4511
timestamp 1682952543
transform 1 0 1388 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4410
timestamp 1682952543
transform 1 0 1436 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4438
timestamp 1682952543
transform 1 0 1428 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4463
timestamp 1682952543
transform 1 0 1420 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4418
timestamp 1682952543
transform 1 0 1428 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4419
timestamp 1682952543
transform 1 0 1436 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4533
timestamp 1682952543
transform 1 0 1444 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4439
timestamp 1682952543
transform 1 0 1460 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4512
timestamp 1682952543
transform 1 0 1460 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4513
timestamp 1682952543
transform 1 0 1468 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1682952543
transform 1 0 1484 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4411
timestamp 1682952543
transform 1 0 1524 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4440
timestamp 1682952543
transform 1 0 1516 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4515
timestamp 1682952543
transform 1 0 1516 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4420
timestamp 1682952543
transform 1 0 1524 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4516
timestamp 1682952543
transform 1 0 1540 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4441
timestamp 1682952543
transform 1 0 1556 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4421
timestamp 1682952543
transform 1 0 1564 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4422
timestamp 1682952543
transform 1 0 1572 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4423
timestamp 1682952543
transform 1 0 1588 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1682952543
transform 1 0 1580 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4468
timestamp 1682952543
transform 1 0 1604 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4518
timestamp 1682952543
transform 1 0 1620 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4442
timestamp 1682952543
transform 1 0 1636 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1682952543
transform 1 0 1652 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4424
timestamp 1682952543
transform 1 0 1636 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4469
timestamp 1682952543
transform 1 0 1636 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4519
timestamp 1682952543
transform 1 0 1668 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4470
timestamp 1682952543
transform 1 0 1700 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4520
timestamp 1682952543
transform 1 0 1716 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4444
timestamp 1682952543
transform 1 0 1740 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4425
timestamp 1682952543
transform 1 0 1740 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4471
timestamp 1682952543
transform 1 0 1740 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4521
timestamp 1682952543
transform 1 0 1780 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1682952543
transform 1 0 1820 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1682952543
transform 1 0 1828 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4499
timestamp 1682952543
transform 1 0 1780 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4500
timestamp 1682952543
transform 1 0 1828 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1682952543
transform 1 0 1820 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4445
timestamp 1682952543
transform 1 0 1844 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1682952543
transform 1 0 1852 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4426
timestamp 1682952543
transform 1 0 1876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4427
timestamp 1682952543
transform 1 0 1884 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4428
timestamp 1682952543
transform 1 0 1900 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1682952543
transform 1 0 1908 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1682952543
transform 1 0 1868 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4535
timestamp 1682952543
transform 1 0 1860 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4524
timestamp 1682952543
transform 1 0 1892 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4536
timestamp 1682952543
transform 1 0 1900 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1682952543
transform 1 0 1932 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1682952543
transform 1 0 1932 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4525
timestamp 1682952543
transform 1 0 1940 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4537
timestamp 1682952543
transform 1 0 1932 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1682952543
transform 1 0 1964 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4430
timestamp 1682952543
transform 1 0 1964 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4431
timestamp 1682952543
transform 1 0 2052 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1682952543
transform 1 0 1964 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4527
timestamp 1682952543
transform 1 0 2028 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4474
timestamp 1682952543
transform 1 0 2052 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4448
timestamp 1682952543
transform 1 0 2068 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4528
timestamp 1682952543
transform 1 0 2068 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4585
timestamp 1682952543
transform 1 0 2068 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4586
timestamp 1682952543
transform 1 0 2084 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1682952543
transform 1 0 2108 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1682952543
transform 1 0 2132 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4529
timestamp 1682952543
transform 1 0 2116 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4434
timestamp 1682952543
transform 1 0 2196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4435
timestamp 1682952543
transform 1 0 2292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4530
timestamp 1682952543
transform 1 0 2204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1682952543
transform 1 0 2212 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1682952543
transform 1 0 2252 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4475
timestamp 1682952543
transform 1 0 2292 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1682952543
transform 1 0 2204 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4502
timestamp 1682952543
transform 1 0 2252 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4436
timestamp 1682952543
transform 1 0 2324 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1682952543
transform 1 0 2364 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1682952543
transform 1 0 2332 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1682952543
transform 1 0 2348 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4535
timestamp 1682952543
transform 1 0 2364 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4503
timestamp 1682952543
transform 1 0 2396 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4438
timestamp 1682952543
transform 1 0 2436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1682952543
transform 1 0 2428 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4476
timestamp 1682952543
transform 1 0 2444 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4439
timestamp 1682952543
transform 1 0 2460 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4504
timestamp 1682952543
transform 1 0 2452 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4538
timestamp 1682952543
transform 1 0 2428 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4537
timestamp 1682952543
transform 1 0 2476 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4553
timestamp 1682952543
transform 1 0 2476 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4440
timestamp 1682952543
transform 1 0 2492 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4538
timestamp 1682952543
transform 1 0 2500 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4539
timestamp 1682952543
transform 1 0 2508 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4505
timestamp 1682952543
transform 1 0 2492 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4540
timestamp 1682952543
transform 1 0 2516 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4539
timestamp 1682952543
transform 1 0 2540 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4441
timestamp 1682952543
transform 1 0 2564 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4442
timestamp 1682952543
transform 1 0 2580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4443
timestamp 1682952543
transform 1 0 2588 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4477
timestamp 1682952543
transform 1 0 2556 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4541
timestamp 1682952543
transform 1 0 2572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1682952543
transform 1 0 2588 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4506
timestamp 1682952543
transform 1 0 2572 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1682952543
transform 1 0 2580 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4380
timestamp 1682952543
transform 1 0 2612 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1682952543
transform 1 0 2612 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1682952543
transform 1 0 2636 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1682952543
transform 1 0 2652 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4412
timestamp 1682952543
transform 1 0 2668 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4446
timestamp 1682952543
transform 1 0 2676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4543
timestamp 1682952543
transform 1 0 2668 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4544
timestamp 1682952543
transform 1 0 2684 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4554
timestamp 1682952543
transform 1 0 2660 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4545
timestamp 1682952543
transform 1 0 2700 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4555
timestamp 1682952543
transform 1 0 2716 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4447
timestamp 1682952543
transform 1 0 2748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1682952543
transform 1 0 2756 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4541
timestamp 1682952543
transform 1 0 2748 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4449
timestamp 1682952543
transform 1 0 2788 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1682952543
transform 1 0 2780 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4547
timestamp 1682952543
transform 1 0 2796 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4507
timestamp 1682952543
transform 1 0 2780 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4450
timestamp 1682952543
transform 1 0 2820 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4508
timestamp 1682952543
transform 1 0 2820 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4413
timestamp 1682952543
transform 1 0 2844 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4548
timestamp 1682952543
transform 1 0 2836 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1682952543
transform 1 0 2844 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4414
timestamp 1682952543
transform 1 0 2876 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1682952543
transform 1 0 2940 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4449
timestamp 1682952543
transform 1 0 2972 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4451
timestamp 1682952543
transform 1 0 2940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1682952543
transform 1 0 2956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1682952543
transform 1 0 2852 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1682952543
transform 1 0 2860 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4552
timestamp 1682952543
transform 1 0 2892 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4509
timestamp 1682952543
transform 1 0 2852 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1682952543
transform 1 0 2892 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4542
timestamp 1682952543
transform 1 0 2860 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_4553
timestamp 1682952543
transform 1 0 2964 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4554
timestamp 1682952543
transform 1 0 2972 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4511
timestamp 1682952543
transform 1 0 2972 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1682952543
transform 1 0 2988 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4453
timestamp 1682952543
transform 1 0 2996 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4454
timestamp 1682952543
transform 1 0 3020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4555
timestamp 1682952543
transform 1 0 3004 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1682952543
transform 1 0 3028 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4416
timestamp 1682952543
transform 1 0 3052 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4455
timestamp 1682952543
transform 1 0 3052 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4557
timestamp 1682952543
transform 1 0 3060 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4478
timestamp 1682952543
transform 1 0 3068 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4512
timestamp 1682952543
transform 1 0 3060 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4456
timestamp 1682952543
transform 1 0 3084 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1682952543
transform 1 0 3100 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4464
timestamp 1682952543
transform 1 0 3108 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4558
timestamp 1682952543
transform 1 0 3124 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4451
timestamp 1682952543
transform 1 0 3140 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4458
timestamp 1682952543
transform 1 0 3140 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4417
timestamp 1682952543
transform 1 0 3308 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1682952543
transform 1 0 3268 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4459
timestamp 1682952543
transform 1 0 3308 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1682952543
transform 1 0 3164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4560
timestamp 1682952543
transform 1 0 3220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4561
timestamp 1682952543
transform 1 0 3228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4562
timestamp 1682952543
transform 1 0 3260 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4543
timestamp 1682952543
transform 1 0 3172 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1682952543
transform 1 0 3324 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4563
timestamp 1682952543
transform 1 0 3324 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4418
timestamp 1682952543
transform 1 0 3412 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4460
timestamp 1682952543
transform 1 0 3412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1682952543
transform 1 0 3364 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4565
timestamp 1682952543
transform 1 0 3380 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4479
timestamp 1682952543
transform 1 0 3388 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4404
timestamp 1682952543
transform 1 0 3484 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1682952543
transform 1 0 3508 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4461
timestamp 1682952543
transform 1 0 3508 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4420
timestamp 1682952543
transform 1 0 3604 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1682952543
transform 1 0 3660 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1682952543
transform 1 0 3740 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4382
timestamp 1682952543
transform 1 0 3636 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_4462
timestamp 1682952543
transform 1 0 3532 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4566
timestamp 1682952543
transform 1 0 3428 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1682952543
transform 1 0 3460 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4568
timestamp 1682952543
transform 1 0 3524 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4556
timestamp 1682952543
transform 1 0 3452 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4557
timestamp 1682952543
transform 1 0 3476 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4558
timestamp 1682952543
transform 1 0 3508 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1682952543
transform 1 0 3644 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4463
timestamp 1682952543
transform 1 0 3644 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1682952543
transform 1 0 3660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4569
timestamp 1682952543
transform 1 0 3548 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4480
timestamp 1682952543
transform 1 0 3572 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4513
timestamp 1682952543
transform 1 0 3548 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4544
timestamp 1682952543
transform 1 0 3604 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4559
timestamp 1682952543
transform 1 0 3588 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4570
timestamp 1682952543
transform 1 0 3708 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4571
timestamp 1682952543
transform 1 0 3740 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4572
timestamp 1682952543
transform 1 0 3748 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4514
timestamp 1682952543
transform 1 0 3708 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4465
timestamp 1682952543
transform 1 0 3764 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4466
timestamp 1682952543
transform 1 0 3772 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4525
timestamp 1682952543
transform 1 0 3756 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4515
timestamp 1682952543
transform 1 0 3772 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4587
timestamp 1682952543
transform 1 0 3788 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1682952543
transform 1 0 3812 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4423
timestamp 1682952543
transform 1 0 3836 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1682952543
transform 1 0 3852 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4383
timestamp 1682952543
transform 1 0 3940 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_4467
timestamp 1682952543
transform 1 0 3828 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4468
timestamp 1682952543
transform 1 0 3836 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4574
timestamp 1682952543
transform 1 0 3844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4575
timestamp 1682952543
transform 1 0 3852 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4516
timestamp 1682952543
transform 1 0 3844 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4469
timestamp 1682952543
transform 1 0 3956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4576
timestamp 1682952543
transform 1 0 3956 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4454
timestamp 1682952543
transform 1 0 4044 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4470
timestamp 1682952543
transform 1 0 4044 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4455
timestamp 1682952543
transform 1 0 4140 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4471
timestamp 1682952543
transform 1 0 4140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4577
timestamp 1682952543
transform 1 0 3996 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1682952543
transform 1 0 4060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1682952543
transform 1 0 4092 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4517
timestamp 1682952543
transform 1 0 4060 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4545
timestamp 1682952543
transform 1 0 3996 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4560
timestamp 1682952543
transform 1 0 4044 0 1 2285
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_36
timestamp 1682952543
transform 1 0 24 0 1 2270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_267
timestamp 1682952543
transform 1 0 72 0 -1 2370
box -8 -3 104 105
use AOI22X1  AOI22X1_156
timestamp 1682952543
transform -1 0 208 0 -1 2370
box -8 -3 46 105
use INVX2  INVX2_304
timestamp 1682952543
transform -1 0 224 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1246
timestamp 1682952543
transform 1 0 224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1682952543
transform 1 0 232 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_157
timestamp 1682952543
transform 1 0 240 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1272
timestamp 1682952543
transform 1 0 280 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4561
timestamp 1682952543
transform 1 0 316 0 1 2275
box -3 -3 3 3
use OAI22X1  OAI22X1_199
timestamp 1682952543
transform -1 0 328 0 -1 2370
box -8 -3 46 105
use INVX2  INVX2_307
timestamp 1682952543
transform -1 0 344 0 -1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_160
timestamp 1682952543
transform 1 0 344 0 -1 2370
box -8 -3 46 105
use INVX2  INVX2_308
timestamp 1682952543
transform 1 0 384 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_268
timestamp 1682952543
transform 1 0 400 0 -1 2370
box -8 -3 104 105
use BUFX2  BUFX2_44
timestamp 1682952543
transform 1 0 496 0 -1 2370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_269
timestamp 1682952543
transform 1 0 520 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_309
timestamp 1682952543
transform -1 0 632 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1273
timestamp 1682952543
transform 1 0 632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1682952543
transform 1 0 640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1682952543
transform 1 0 648 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1276
timestamp 1682952543
transform 1 0 656 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_161
timestamp 1682952543
transform 1 0 664 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_162
timestamp 1682952543
transform 1 0 704 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1277
timestamp 1682952543
transform 1 0 744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1279
timestamp 1682952543
transform 1 0 752 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1281
timestamp 1682952543
transform 1 0 760 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1682952543
transform 1 0 768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1283
timestamp 1682952543
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_163
timestamp 1682952543
transform 1 0 784 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1285
timestamp 1682952543
transform 1 0 824 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1286
timestamp 1682952543
transform 1 0 832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1682952543
transform 1 0 840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1682952543
transform 1 0 848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1682952543
transform 1 0 856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1290
timestamp 1682952543
transform 1 0 864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1682952543
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1682952543
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_54
timestamp 1682952543
transform 1 0 888 0 -1 2370
box -8 -3 34 105
use FILL  FILL_1295
timestamp 1682952543
transform 1 0 920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1297
timestamp 1682952543
transform 1 0 928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1682952543
transform 1 0 936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1682952543
transform 1 0 944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1682952543
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1682952543
transform 1 0 960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1306
timestamp 1682952543
transform 1 0 968 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_55
timestamp 1682952543
transform 1 0 976 0 -1 2370
box -8 -3 32 105
use FILL  FILL_1307
timestamp 1682952543
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1309
timestamp 1682952543
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1682952543
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1313
timestamp 1682952543
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1682952543
transform 1 0 1032 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1682952543
transform 1 0 1040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1319
timestamp 1682952543
transform 1 0 1048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1682952543
transform 1 0 1056 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_55
timestamp 1682952543
transform 1 0 1064 0 -1 2370
box -8 -3 34 105
use FILL  FILL_1324
timestamp 1682952543
transform 1 0 1096 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1682952543
transform 1 0 1104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1682952543
transform 1 0 1112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1682952543
transform 1 0 1120 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1682952543
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1682952543
transform 1 0 1136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1334
timestamp 1682952543
transform 1 0 1144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1682952543
transform 1 0 1152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1682952543
transform 1 0 1160 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_57
timestamp 1682952543
transform -1 0 1200 0 -1 2370
box -8 -3 34 105
use FILL  FILL_1342
timestamp 1682952543
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1343
timestamp 1682952543
transform 1 0 1208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1682952543
transform 1 0 1216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1346
timestamp 1682952543
transform 1 0 1224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1682952543
transform 1 0 1232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1682952543
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1682952543
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1682952543
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1682952543
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1360
timestamp 1682952543
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_58
timestamp 1682952543
transform -1 0 1312 0 -1 2370
box -8 -3 34 105
use FILL  FILL_1361
timestamp 1682952543
transform 1 0 1312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1682952543
transform 1 0 1320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1364
timestamp 1682952543
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1682952543
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1682952543
transform 1 0 1344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1367
timestamp 1682952543
transform 1 0 1352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1682952543
transform 1 0 1360 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_311
timestamp 1682952543
transform 1 0 1368 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1369
timestamp 1682952543
transform 1 0 1384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1682952543
transform 1 0 1392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1682952543
transform 1 0 1400 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_48
timestamp 1682952543
transform 1 0 1408 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1386
timestamp 1682952543
transform 1 0 1432 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_52
timestamp 1682952543
transform -1 0 1464 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1387
timestamp 1682952543
transform 1 0 1464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1682952543
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_53
timestamp 1682952543
transform 1 0 1480 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1389
timestamp 1682952543
transform 1 0 1504 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4562
timestamp 1682952543
transform 1 0 1524 0 1 2275
box -3 -3 3 3
use FILL  FILL_1390
timestamp 1682952543
transform 1 0 1512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1682952543
transform 1 0 1520 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_314
timestamp 1682952543
transform -1 0 1544 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1392
timestamp 1682952543
transform 1 0 1544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1682952543
transform 1 0 1552 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_169
timestamp 1682952543
transform 1 0 1560 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1394
timestamp 1682952543
transform 1 0 1600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1682952543
transform 1 0 1608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1682952543
transform 1 0 1616 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_272
timestamp 1682952543
transform 1 0 1624 0 -1 2370
box -8 -3 104 105
use FILL  FILL_1397
timestamp 1682952543
transform 1 0 1720 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4563
timestamp 1682952543
transform 1 0 1812 0 1 2275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_273
timestamp 1682952543
transform 1 0 1728 0 -1 2370
box -8 -3 104 105
use M3_M2  M3_M2_4564
timestamp 1682952543
transform 1 0 1844 0 1 2275
box -3 -3 3 3
use INVX2  INVX2_315
timestamp 1682952543
transform -1 0 1840 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1398
timestamp 1682952543
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1682952543
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1682952543
transform 1 0 1856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1402
timestamp 1682952543
transform 1 0 1864 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_171
timestamp 1682952543
transform 1 0 1872 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1405
timestamp 1682952543
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1406
timestamp 1682952543
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1682952543
transform 1 0 1928 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_55
timestamp 1682952543
transform 1 0 1936 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1426
timestamp 1682952543
transform 1 0 1960 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_274
timestamp 1682952543
transform -1 0 2064 0 -1 2370
box -8 -3 104 105
use FILL  FILL_1427
timestamp 1682952543
transform 1 0 2064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1682952543
transform 1 0 2072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1682952543
transform 1 0 2080 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_56
timestamp 1682952543
transform 1 0 2088 0 -1 2370
box -5 -3 28 105
use BUFX2  BUFX2_57
timestamp 1682952543
transform 1 0 2112 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1430
timestamp 1682952543
transform 1 0 2136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1682952543
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1432
timestamp 1682952543
transform 1 0 2152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1682952543
transform 1 0 2160 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1682952543
transform 1 0 2168 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1435
timestamp 1682952543
transform 1 0 2176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1437
timestamp 1682952543
transform 1 0 2184 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_317
timestamp 1682952543
transform 1 0 2192 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_276
timestamp 1682952543
transform -1 0 2304 0 -1 2370
box -8 -3 104 105
use FILL  FILL_1443
timestamp 1682952543
transform 1 0 2304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1682952543
transform 1 0 2312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1445
timestamp 1682952543
transform 1 0 2320 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_173
timestamp 1682952543
transform 1 0 2328 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1449
timestamp 1682952543
transform 1 0 2368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1682952543
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1682952543
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1452
timestamp 1682952543
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4565
timestamp 1682952543
transform 1 0 2412 0 1 2275
box -3 -3 3 3
use FILL  FILL_1453
timestamp 1682952543
transform 1 0 2400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1682952543
transform 1 0 2408 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_200
timestamp 1682952543
transform -1 0 2456 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1455
timestamp 1682952543
transform 1 0 2456 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1461
timestamp 1682952543
transform 1 0 2464 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1682952543
transform 1 0 2472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1682952543
transform 1 0 2480 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_319
timestamp 1682952543
transform 1 0 2488 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1464
timestamp 1682952543
transform 1 0 2504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1465
timestamp 1682952543
transform 1 0 2512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1682952543
transform 1 0 2520 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1467
timestamp 1682952543
transform 1 0 2528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1682952543
transform 1 0 2536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1469
timestamp 1682952543
transform 1 0 2544 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_174
timestamp 1682952543
transform 1 0 2552 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1470
timestamp 1682952543
transform 1 0 2592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1471
timestamp 1682952543
transform 1 0 2600 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4566
timestamp 1682952543
transform 1 0 2620 0 1 2275
box -3 -3 3 3
use FILL  FILL_1472
timestamp 1682952543
transform 1 0 2608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1473
timestamp 1682952543
transform 1 0 2616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1682952543
transform 1 0 2624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1475
timestamp 1682952543
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1682952543
transform 1 0 2640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1682952543
transform 1 0 2648 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_203
timestamp 1682952543
transform 1 0 2656 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1486
timestamp 1682952543
transform 1 0 2696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1487
timestamp 1682952543
transform 1 0 2704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1682952543
transform 1 0 2712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1682952543
transform 1 0 2720 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4567
timestamp 1682952543
transform 1 0 2740 0 1 2275
box -3 -3 3 3
use FILL  FILL_1490
timestamp 1682952543
transform 1 0 2728 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1682952543
transform 1 0 2736 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1682952543
transform 1 0 2744 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1682952543
transform 1 0 2752 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_177
timestamp 1682952543
transform 1 0 2760 0 -1 2370
box -8 -3 46 105
use FILL  FILL_1501
timestamp 1682952543
transform 1 0 2800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1502
timestamp 1682952543
transform 1 0 2808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1682952543
transform 1 0 2816 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4568
timestamp 1682952543
transform 1 0 2844 0 1 2275
box -3 -3 3 3
use INVX2  INVX2_321
timestamp 1682952543
transform 1 0 2824 0 -1 2370
box -9 -3 26 105
use INVX2  INVX2_322
timestamp 1682952543
transform 1 0 2840 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_283
timestamp 1682952543
transform -1 0 2952 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_323
timestamp 1682952543
transform 1 0 2952 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1504
timestamp 1682952543
transform 1 0 2968 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_59
timestamp 1682952543
transform 1 0 2976 0 -1 2370
box -5 -3 28 105
use M3_M2  M3_M2_4569
timestamp 1682952543
transform 1 0 3028 0 1 2275
box -3 -3 3 3
use BUFX2  BUFX2_60
timestamp 1682952543
transform 1 0 3000 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1505
timestamp 1682952543
transform 1 0 3024 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_61
timestamp 1682952543
transform 1 0 3032 0 -1 2370
box -5 -3 28 105
use M3_M2  M3_M2_4570
timestamp 1682952543
transform 1 0 3068 0 1 2275
box -3 -3 3 3
use FILL  FILL_1506
timestamp 1682952543
transform 1 0 3056 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_62
timestamp 1682952543
transform 1 0 3064 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1507
timestamp 1682952543
transform 1 0 3088 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_324
timestamp 1682952543
transform 1 0 3096 0 -1 2370
box -9 -3 26 105
use FILL  FILL_1508
timestamp 1682952543
transform 1 0 3112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1682952543
transform 1 0 3120 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_284
timestamp 1682952543
transform 1 0 3128 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_285
timestamp 1682952543
transform -1 0 3320 0 -1 2370
box -8 -3 104 105
use FILL  FILL_1510
timestamp 1682952543
transform 1 0 3320 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_286
timestamp 1682952543
transform -1 0 3424 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_287
timestamp 1682952543
transform -1 0 3520 0 -1 2370
box -8 -3 104 105
use FILL  FILL_1511
timestamp 1682952543
transform 1 0 3520 0 -1 2370
box -8 -3 16 105
use FAX1  FAX1_22
timestamp 1682952543
transform 1 0 3528 0 -1 2370
box -5 -3 126 105
use DFFNEGX1  DFFNEGX1_288
timestamp 1682952543
transform 1 0 3648 0 -1 2370
box -8 -3 104 105
use BUFX2  BUFX2_63
timestamp 1682952543
transform 1 0 3744 0 -1 2370
box -5 -3 28 105
use FILL  FILL_1512
timestamp 1682952543
transform 1 0 3768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1682952543
transform 1 0 3776 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_64
timestamp 1682952543
transform -1 0 3816 0 -1 2370
box -8 -3 34 105
use FILL  FILL_1514
timestamp 1682952543
transform 1 0 3816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1682952543
transform 1 0 3824 0 -1 2370
box -8 -3 16 105
use FAX1  FAX1_23
timestamp 1682952543
transform 1 0 3832 0 -1 2370
box -5 -3 126 105
use FILL  FILL_1516
timestamp 1682952543
transform 1 0 3952 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_289
timestamp 1682952543
transform -1 0 4056 0 -1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_290
timestamp 1682952543
transform -1 0 4152 0 -1 2370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_37
timestamp 1682952543
transform 1 0 4201 0 1 2270
box -10 -3 10 3
use M3_M2  M3_M2_4578
timestamp 1682952543
transform 1 0 228 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4608
timestamp 1682952543
transform 1 0 172 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1682952543
transform 1 0 204 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_4606
timestamp 1682952543
transform 1 0 116 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4607
timestamp 1682952543
transform 1 0 164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1682952543
transform 1 0 212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1682952543
transform 1 0 84 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4672
timestamp 1682952543
transform 1 0 84 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4711
timestamp 1682952543
transform 1 0 180 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4673
timestamp 1682952543
transform 1 0 180 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1682952543
transform 1 0 196 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4675
timestamp 1682952543
transform 1 0 220 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4609
timestamp 1682952543
transform 1 0 268 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4664
timestamp 1682952543
transform 1 0 268 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1682952543
transform 1 0 300 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_4610
timestamp 1682952543
transform 1 0 324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1682952543
transform 1 0 372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4712
timestamp 1682952543
transform 1 0 292 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4676
timestamp 1682952543
transform 1 0 292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1682952543
transform 1 0 324 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1682952543
transform 1 0 396 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1682952543
transform 1 0 428 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4610
timestamp 1682952543
transform 1 0 412 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4624
timestamp 1682952543
transform 1 0 412 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4612
timestamp 1682952543
transform 1 0 388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1682952543
transform 1 0 404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4614
timestamp 1682952543
transform 1 0 428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1682952543
transform 1 0 380 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1682952543
transform 1 0 412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1682952543
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4611
timestamp 1682952543
transform 1 0 444 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_4615
timestamp 1682952543
transform 1 0 436 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4716
timestamp 1682952543
transform 1 0 444 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4612
timestamp 1682952543
transform 1 0 476 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1682952543
transform 1 0 492 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4616
timestamp 1682952543
transform 1 0 492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4717
timestamp 1682952543
transform 1 0 484 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4678
timestamp 1682952543
transform 1 0 484 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1682952543
transform 1 0 508 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4613
timestamp 1682952543
transform 1 0 556 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1682952543
transform 1 0 524 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4617
timestamp 1682952543
transform 1 0 516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1682952543
transform 1 0 540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1682952543
transform 1 0 556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1682952543
transform 1 0 524 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1682952543
transform 1 0 548 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4665
timestamp 1682952543
transform 1 0 556 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_4720
timestamp 1682952543
transform 1 0 564 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4679
timestamp 1682952543
transform 1 0 548 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4620
timestamp 1682952543
transform 1 0 580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1682952543
transform 1 0 612 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4593
timestamp 1682952543
transform 1 0 644 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4627
timestamp 1682952543
transform 1 0 644 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1682952543
transform 1 0 676 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4622
timestamp 1682952543
transform 1 0 652 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1682952543
transform 1 0 676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1682952543
transform 1 0 636 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1682952543
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1682952543
transform 1 0 660 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4724
timestamp 1682952543
transform 1 0 668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4725
timestamp 1682952543
transform 1 0 676 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4716
timestamp 1682952543
transform 1 0 668 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4594
timestamp 1682952543
transform 1 0 708 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_4624
timestamp 1682952543
transform 1 0 700 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4717
timestamp 1682952543
transform 1 0 700 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4596
timestamp 1682952543
transform 1 0 724 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4680
timestamp 1682952543
transform 1 0 740 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4788
timestamp 1682952543
transform 1 0 748 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4573
timestamp 1682952543
transform 1 0 764 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_4625
timestamp 1682952543
transform 1 0 756 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4580
timestamp 1682952543
transform 1 0 772 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4574
timestamp 1682952543
transform 1 0 804 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_4626
timestamp 1682952543
transform 1 0 836 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4681
timestamp 1682952543
transform 1 0 836 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4718
timestamp 1682952543
transform 1 0 836 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4595
timestamp 1682952543
transform 1 0 860 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4614
timestamp 1682952543
transform 1 0 868 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_4627
timestamp 1682952543
transform 1 0 860 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1682952543
transform 1 0 852 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4682
timestamp 1682952543
transform 1 0 868 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4590
timestamp 1682952543
transform 1 0 884 0 1 2255
box -2 -2 2 2
use M3_M2  M3_M2_4596
timestamp 1682952543
transform 1 0 884 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4719
timestamp 1682952543
transform 1 0 876 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4628
timestamp 1682952543
transform 1 0 900 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4597
timestamp 1682952543
transform 1 0 964 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_4629
timestamp 1682952543
transform 1 0 956 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4630
timestamp 1682952543
transform 1 0 972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1682952543
transform 1 0 940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1682952543
transform 1 0 948 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1682952543
transform 1 0 964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1682952543
transform 1 0 972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1682952543
transform 1 0 980 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4666
timestamp 1682952543
transform 1 0 996 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_4790
timestamp 1682952543
transform 1 0 996 0 1 2195
box -2 -2 2 2
use M3_M2  M3_M2_4629
timestamp 1682952543
transform 1 0 1036 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4631
timestamp 1682952543
transform 1 0 1036 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4683
timestamp 1682952543
transform 1 0 1036 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4575
timestamp 1682952543
transform 1 0 1132 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4576
timestamp 1682952543
transform 1 0 1148 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4581
timestamp 1682952543
transform 1 0 1052 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4598
timestamp 1682952543
transform 1 0 1052 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4630
timestamp 1682952543
transform 1 0 1084 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4631
timestamp 1682952543
transform 1 0 1148 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4632
timestamp 1682952543
transform 1 0 1052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1682952543
transform 1 0 1084 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4634
timestamp 1682952543
transform 1 0 1148 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4667
timestamp 1682952543
transform 1 0 1108 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_4731
timestamp 1682952543
transform 1 0 1132 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4684
timestamp 1682952543
transform 1 0 1100 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4720
timestamp 1682952543
transform 1 0 1140 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4732
timestamp 1682952543
transform 1 0 1164 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4685
timestamp 1682952543
transform 1 0 1164 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4721
timestamp 1682952543
transform 1 0 1228 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4647
timestamp 1682952543
transform 1 0 1252 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4635
timestamp 1682952543
transform 1 0 1276 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4733
timestamp 1682952543
transform 1 0 1252 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4686
timestamp 1682952543
transform 1 0 1252 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4722
timestamp 1682952543
transform 1 0 1252 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4668
timestamp 1682952543
transform 1 0 1340 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_4636
timestamp 1682952543
transform 1 0 1356 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4637
timestamp 1682952543
transform 1 0 1364 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4638
timestamp 1682952543
transform 1 0 1404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1682952543
transform 1 0 1444 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4687
timestamp 1682952543
transform 1 0 1364 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1682952543
transform 1 0 1404 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4723
timestamp 1682952543
transform 1 0 1412 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4639
timestamp 1682952543
transform 1 0 1516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1682952543
transform 1 0 1468 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4582
timestamp 1682952543
transform 1 0 1596 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1682952543
transform 1 0 1620 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4640
timestamp 1682952543
transform 1 0 1580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1682952543
transform 1 0 1588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1682952543
transform 1 0 1604 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1682952543
transform 1 0 1620 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4736
timestamp 1682952543
transform 1 0 1572 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1682952543
transform 1 0 1596 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1682952543
transform 1 0 1612 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4689
timestamp 1682952543
transform 1 0 1596 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1682952543
transform 1 0 1612 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4739
timestamp 1682952543
transform 1 0 1628 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4690
timestamp 1682952543
transform 1 0 1628 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4583
timestamp 1682952543
transform 1 0 1660 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4599
timestamp 1682952543
transform 1 0 1660 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_4644
timestamp 1682952543
transform 1 0 1644 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4648
timestamp 1682952543
transform 1 0 1652 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1682952543
transform 1 0 1692 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4645
timestamp 1682952543
transform 1 0 1660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1682952543
transform 1 0 1676 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4649
timestamp 1682952543
transform 1 0 1684 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4647
timestamp 1682952543
transform 1 0 1692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1682952543
transform 1 0 1668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1682952543
transform 1 0 1684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1682952543
transform 1 0 1692 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4691
timestamp 1682952543
transform 1 0 1668 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4725
timestamp 1682952543
transform 1 0 1668 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4648
timestamp 1682952543
transform 1 0 1708 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4650
timestamp 1682952543
transform 1 0 1716 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4743
timestamp 1682952543
transform 1 0 1716 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4692
timestamp 1682952543
transform 1 0 1716 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4649
timestamp 1682952543
transform 1 0 1740 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4600
timestamp 1682952543
transform 1 0 1772 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4634
timestamp 1682952543
transform 1 0 1780 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4651
timestamp 1682952543
transform 1 0 1756 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4650
timestamp 1682952543
transform 1 0 1764 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4652
timestamp 1682952543
transform 1 0 1772 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4651
timestamp 1682952543
transform 1 0 1780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4744
timestamp 1682952543
transform 1 0 1772 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1682952543
transform 1 0 1780 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4726
timestamp 1682952543
transform 1 0 1780 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4652
timestamp 1682952543
transform 1 0 1820 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4653
timestamp 1682952543
transform 1 0 1844 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4746
timestamp 1682952543
transform 1 0 1852 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4693
timestamp 1682952543
transform 1 0 1852 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4727
timestamp 1682952543
transform 1 0 1844 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1682952543
transform 1 0 1900 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4653
timestamp 1682952543
transform 1 0 1868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1682952543
transform 1 0 1884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1682952543
transform 1 0 1900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1682952543
transform 1 0 1916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4747
timestamp 1682952543
transform 1 0 1916 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4654
timestamp 1682952543
transform 1 0 1932 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4748
timestamp 1682952543
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4694
timestamp 1682952543
transform 1 0 1940 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4636
timestamp 1682952543
transform 1 0 1980 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4657
timestamp 1682952543
transform 1 0 1964 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4655
timestamp 1682952543
transform 1 0 1972 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4658
timestamp 1682952543
transform 1 0 1980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1682952543
transform 1 0 1972 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1682952543
transform 1 0 1980 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4584
timestamp 1682952543
transform 1 0 1996 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_4659
timestamp 1682952543
transform 1 0 2028 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4585
timestamp 1682952543
transform 1 0 2052 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4601
timestamp 1682952543
transform 1 0 2060 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_4660
timestamp 1682952543
transform 1 0 2044 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4656
timestamp 1682952543
transform 1 0 2052 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4586
timestamp 1682952543
transform 1 0 2084 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4657
timestamp 1682952543
transform 1 0 2076 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4587
timestamp 1682952543
transform 1 0 2116 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4602
timestamp 1682952543
transform 1 0 2116 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4658
timestamp 1682952543
transform 1 0 2108 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4661
timestamp 1682952543
transform 1 0 2116 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4659
timestamp 1682952543
transform 1 0 2124 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4662
timestamp 1682952543
transform 1 0 2132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1682952543
transform 1 0 2116 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1682952543
transform 1 0 2124 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1682952543
transform 1 0 2140 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4695
timestamp 1682952543
transform 1 0 2108 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1682952543
transform 1 0 2156 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4663
timestamp 1682952543
transform 1 0 2156 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4603
timestamp 1682952543
transform 1 0 2204 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_4664
timestamp 1682952543
transform 1 0 2204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1682952543
transform 1 0 2220 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4660
timestamp 1682952543
transform 1 0 2228 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4666
timestamp 1682952543
transform 1 0 2236 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1682952543
transform 1 0 2212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1682952543
transform 1 0 2228 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4756
timestamp 1682952543
transform 1 0 2252 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4757
timestamp 1682952543
transform 1 0 2260 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4667
timestamp 1682952543
transform 1 0 2284 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4661
timestamp 1682952543
transform 1 0 2292 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4668
timestamp 1682952543
transform 1 0 2300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1682952543
transform 1 0 2324 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4604
timestamp 1682952543
transform 1 0 2364 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1682952543
transform 1 0 2388 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4638
timestamp 1682952543
transform 1 0 2372 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4670
timestamp 1682952543
transform 1 0 2356 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4662
timestamp 1682952543
transform 1 0 2364 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4671
timestamp 1682952543
transform 1 0 2372 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1682952543
transform 1 0 2388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4758
timestamp 1682952543
transform 1 0 2364 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4728
timestamp 1682952543
transform 1 0 2356 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4759
timestamp 1682952543
transform 1 0 2396 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4696
timestamp 1682952543
transform 1 0 2396 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1682952543
transform 1 0 2412 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4639
timestamp 1682952543
transform 1 0 2420 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4760
timestamp 1682952543
transform 1 0 2420 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4730
timestamp 1682952543
transform 1 0 2428 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4640
timestamp 1682952543
transform 1 0 2460 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1682952543
transform 1 0 2500 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4673
timestamp 1682952543
transform 1 0 2460 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1682952543
transform 1 0 2468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4675
timestamp 1682952543
transform 1 0 2500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4761
timestamp 1682952543
transform 1 0 2548 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4697
timestamp 1682952543
transform 1 0 2468 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1682952543
transform 1 0 2508 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1682952543
transform 1 0 2500 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1682952543
transform 1 0 2564 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_4762
timestamp 1682952543
transform 1 0 2564 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4588
timestamp 1682952543
transform 1 0 2588 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1682952543
transform 1 0 2588 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_4676
timestamp 1682952543
transform 1 0 2588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4763
timestamp 1682952543
transform 1 0 2588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4699
timestamp 1682952543
transform 1 0 2588 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4764
timestamp 1682952543
transform 1 0 2604 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4700
timestamp 1682952543
transform 1 0 2604 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4615
timestamp 1682952543
transform 1 0 2668 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_4677
timestamp 1682952543
transform 1 0 2644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1682952543
transform 1 0 2660 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4589
timestamp 1682952543
transform 1 0 2684 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_4597
timestamp 1682952543
transform 1 0 2684 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4765
timestamp 1682952543
transform 1 0 2668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1682952543
transform 1 0 2676 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4701
timestamp 1682952543
transform 1 0 2676 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4732
timestamp 1682952543
transform 1 0 2668 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4679
timestamp 1682952543
transform 1 0 2700 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4702
timestamp 1682952543
transform 1 0 2700 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4591
timestamp 1682952543
transform 1 0 2716 0 1 2235
box -2 -2 2 2
use M3_M2  M3_M2_4590
timestamp 1682952543
transform 1 0 2788 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4616
timestamp 1682952543
transform 1 0 2764 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4617
timestamp 1682952543
transform 1 0 2788 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4618
timestamp 1682952543
transform 1 0 2812 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1682952543
transform 1 0 2732 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4643
timestamp 1682952543
transform 1 0 2756 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_4680
timestamp 1682952543
transform 1 0 2724 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1682952543
transform 1 0 2740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4682
timestamp 1682952543
transform 1 0 2764 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4767
timestamp 1682952543
transform 1 0 2732 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4768
timestamp 1682952543
transform 1 0 2748 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4769
timestamp 1682952543
transform 1 0 2756 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4703
timestamp 1682952543
transform 1 0 2756 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4644
timestamp 1682952543
transform 1 0 2772 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4645
timestamp 1682952543
transform 1 0 2812 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1682952543
transform 1 0 2900 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4592
timestamp 1682952543
transform 1 0 3052 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4619
timestamp 1682952543
transform 1 0 2964 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1682952543
transform 1 0 3028 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_4683
timestamp 1682952543
transform 1 0 2772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4684
timestamp 1682952543
transform 1 0 2780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4685
timestamp 1682952543
transform 1 0 2812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1682952543
transform 1 0 2876 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1682952543
transform 1 0 2932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4770
timestamp 1682952543
transform 1 0 2860 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4704
timestamp 1682952543
transform 1 0 2860 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4733
timestamp 1682952543
transform 1 0 2780 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4771
timestamp 1682952543
transform 1 0 2956 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4705
timestamp 1682952543
transform 1 0 2956 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4688
timestamp 1682952543
transform 1 0 3004 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4689
timestamp 1682952543
transform 1 0 3060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1682952543
transform 1 0 3068 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4772
timestamp 1682952543
transform 1 0 2980 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4734
timestamp 1682952543
transform 1 0 2980 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4706
timestamp 1682952543
transform 1 0 3068 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4691
timestamp 1682952543
transform 1 0 3148 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1682952543
transform 1 0 3100 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1682952543
transform 1 0 3116 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4707
timestamp 1682952543
transform 1 0 3116 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4735
timestamp 1682952543
transform 1 0 3100 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4692
timestamp 1682952543
transform 1 0 3212 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4693
timestamp 1682952543
transform 1 0 3252 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1682952543
transform 1 0 3228 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4708
timestamp 1682952543
transform 1 0 3228 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4694
timestamp 1682952543
transform 1 0 3332 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4607
timestamp 1682952543
transform 1 0 3356 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_4592
timestamp 1682952543
transform 1 0 3356 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1682952543
transform 1 0 3348 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4599
timestamp 1682952543
transform 1 0 3372 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1682952543
transform 1 0 3364 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1682952543
transform 1 0 3484 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4600
timestamp 1682952543
transform 1 0 3476 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4695
timestamp 1682952543
transform 1 0 3436 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1682952543
transform 1 0 3468 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4777
timestamp 1682952543
transform 1 0 3388 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4709
timestamp 1682952543
transform 1 0 3436 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4736
timestamp 1682952543
transform 1 0 3388 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4737
timestamp 1682952543
transform 1 0 3436 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1682952543
transform 1 0 3548 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1682952543
transform 1 0 3564 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_4601
timestamp 1682952543
transform 1 0 3500 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4577
timestamp 1682952543
transform 1 0 3612 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_4594
timestamp 1682952543
transform 1 0 3612 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4602
timestamp 1682952543
transform 1 0 3604 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1682952543
transform 1 0 3508 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1682952543
transform 1 0 3564 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1682952543
transform 1 0 3492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1682952543
transform 1 0 3588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4710
timestamp 1682952543
transform 1 0 3508 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1682952543
transform 1 0 3636 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_4595
timestamp 1682952543
transform 1 0 3644 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_4603
timestamp 1682952543
transform 1 0 3628 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1682952543
transform 1 0 3636 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4780
timestamp 1682952543
transform 1 0 3620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4605
timestamp 1682952543
transform 1 0 3660 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1682952543
transform 1 0 3652 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4669
timestamp 1682952543
transform 1 0 3644 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4738
timestamp 1682952543
transform 1 0 3652 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4700
timestamp 1682952543
transform 1 0 3700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4781
timestamp 1682952543
transform 1 0 3676 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4711
timestamp 1682952543
transform 1 0 3676 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1682952543
transform 1 0 3692 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4740
timestamp 1682952543
transform 1 0 3716 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4701
timestamp 1682952543
transform 1 0 3772 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4702
timestamp 1682952543
transform 1 0 3836 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1682952543
transform 1 0 3884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1682952543
transform 1 0 3932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4705
timestamp 1682952543
transform 1 0 3980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1682952543
transform 1 0 3996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1682952543
transform 1 0 4012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4782
timestamp 1682952543
transform 1 0 3788 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4670
timestamp 1682952543
transform 1 0 3836 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4671
timestamp 1682952543
transform 1 0 3868 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4712
timestamp 1682952543
transform 1 0 3788 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_4708
timestamp 1682952543
transform 1 0 4060 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1682952543
transform 1 0 3900 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4784
timestamp 1682952543
transform 1 0 3988 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1682952543
transform 1 0 4004 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4786
timestamp 1682952543
transform 1 0 4020 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1682952543
transform 1 0 4036 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4713
timestamp 1682952543
transform 1 0 3988 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4714
timestamp 1682952543
transform 1 0 4004 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4741
timestamp 1682952543
transform 1 0 3900 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4715
timestamp 1682952543
transform 1 0 4060 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4742
timestamp 1682952543
transform 1 0 4036 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4743
timestamp 1682952543
transform 1 0 4068 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_4709
timestamp 1682952543
transform 1 0 4132 0 1 2215
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_38
timestamp 1682952543
transform 1 0 48 0 1 2170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_291
timestamp 1682952543
transform 1 0 72 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_292
timestamp 1682952543
transform 1 0 168 0 1 2170
box -8 -3 104 105
use FILL  FILL_1517
timestamp 1682952543
transform 1 0 264 0 1 2170
box -8 -3 16 105
use FILL  FILL_1518
timestamp 1682952543
transform 1 0 272 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_293
timestamp 1682952543
transform 1 0 280 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4744
timestamp 1682952543
transform 1 0 388 0 1 2175
box -3 -3 3 3
use FILL  FILL_1519
timestamp 1682952543
transform 1 0 376 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_180
timestamp 1682952543
transform 1 0 384 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_329
timestamp 1682952543
transform 1 0 424 0 1 2170
box -9 -3 26 105
use FILL  FILL_1536
timestamp 1682952543
transform 1 0 440 0 1 2170
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1682952543
transform 1 0 448 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_64
timestamp 1682952543
transform -1 0 480 0 1 2170
box -5 -3 28 105
use FILL  FILL_1538
timestamp 1682952543
transform 1 0 480 0 1 2170
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1682952543
transform 1 0 488 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_65
timestamp 1682952543
transform -1 0 520 0 1 2170
box -5 -3 28 105
use FILL  FILL_1540
timestamp 1682952543
transform 1 0 520 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_205
timestamp 1682952543
transform 1 0 528 0 1 2170
box -8 -3 46 105
use FILL  FILL_1541
timestamp 1682952543
transform 1 0 568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1542
timestamp 1682952543
transform 1 0 576 0 1 2170
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1682952543
transform 1 0 584 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4745
timestamp 1682952543
transform 1 0 612 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_330
timestamp 1682952543
transform -1 0 608 0 1 2170
box -9 -3 26 105
use FILL  FILL_1544
timestamp 1682952543
transform 1 0 608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1682952543
transform 1 0 616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1682952543
transform 1 0 624 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_182
timestamp 1682952543
transform 1 0 632 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_331
timestamp 1682952543
transform 1 0 672 0 1 2170
box -9 -3 26 105
use FILL  FILL_1549
timestamp 1682952543
transform 1 0 688 0 1 2170
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1682952543
transform 1 0 696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1682952543
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1682952543
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1682952543
transform 1 0 720 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_332
timestamp 1682952543
transform 1 0 728 0 1 2170
box -9 -3 26 105
use FILL  FILL_1560
timestamp 1682952543
transform 1 0 744 0 1 2170
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1682952543
transform 1 0 752 0 1 2170
box -8 -3 16 105
use FILL  FILL_1562
timestamp 1682952543
transform 1 0 760 0 1 2170
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1682952543
transform 1 0 768 0 1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_58
timestamp 1682952543
transform 1 0 776 0 1 2170
box -8 -3 32 105
use FILL  FILL_1564
timestamp 1682952543
transform 1 0 800 0 1 2170
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1682952543
transform 1 0 808 0 1 2170
box -8 -3 16 105
use FILL  FILL_1566
timestamp 1682952543
transform 1 0 816 0 1 2170
box -8 -3 16 105
use FILL  FILL_1568
timestamp 1682952543
transform 1 0 824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1682952543
transform 1 0 832 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_184
timestamp 1682952543
transform 1 0 840 0 1 2170
box -8 -3 46 105
use FILL  FILL_1571
timestamp 1682952543
transform 1 0 880 0 1 2170
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1682952543
transform 1 0 888 0 1 2170
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1682952543
transform 1 0 896 0 1 2170
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1682952543
transform 1 0 904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1682952543
transform 1 0 912 0 1 2170
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1682952543
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_1583
timestamp 1682952543
transform 1 0 928 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4746
timestamp 1682952543
transform 1 0 964 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_185
timestamp 1682952543
transform 1 0 936 0 1 2170
box -8 -3 46 105
use FILL  FILL_1584
timestamp 1682952543
transform 1 0 976 0 1 2170
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1682952543
transform 1 0 984 0 1 2170
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1682952543
transform 1 0 992 0 1 2170
box -8 -3 16 105
use FILL  FILL_1593
timestamp 1682952543
transform 1 0 1000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1682952543
transform 1 0 1008 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_333
timestamp 1682952543
transform 1 0 1016 0 1 2170
box -9 -3 26 105
use FILL  FILL_1595
timestamp 1682952543
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1682952543
transform 1 0 1040 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4747
timestamp 1682952543
transform 1 0 1092 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_297
timestamp 1682952543
transform -1 0 1144 0 1 2170
box -8 -3 104 105
use BUFX2  BUFX2_66
timestamp 1682952543
transform 1 0 1144 0 1 2170
box -5 -3 28 105
use FILL  FILL_1599
timestamp 1682952543
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1600
timestamp 1682952543
transform 1 0 1176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1682952543
transform 1 0 1184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1682952543
transform 1 0 1192 0 1 2170
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1682952543
transform 1 0 1200 0 1 2170
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1682952543
transform 1 0 1208 0 1 2170
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1682952543
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_1621
timestamp 1682952543
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1682952543
transform 1 0 1232 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_298
timestamp 1682952543
transform 1 0 1240 0 1 2170
box -8 -3 104 105
use FILL  FILL_1625
timestamp 1682952543
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_334
timestamp 1682952543
transform 1 0 1344 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_299
timestamp 1682952543
transform -1 0 1456 0 1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_300
timestamp 1682952543
transform 1 0 1456 0 1 2170
box -8 -3 104 105
use FILL  FILL_1626
timestamp 1682952543
transform 1 0 1552 0 1 2170
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1682952543
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1682952543
transform 1 0 1568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1682952543
transform 1 0 1576 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_187
timestamp 1682952543
transform 1 0 1584 0 1 2170
box -8 -3 46 105
use FILL  FILL_1647
timestamp 1682952543
transform 1 0 1624 0 1 2170
box -8 -3 16 105
use FILL  FILL_1648
timestamp 1682952543
transform 1 0 1632 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4748
timestamp 1682952543
transform 1 0 1652 0 1 2175
box -3 -3 3 3
use FILL  FILL_1649
timestamp 1682952543
transform 1 0 1640 0 1 2170
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1682952543
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4749
timestamp 1682952543
transform 1 0 1700 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_189
timestamp 1682952543
transform 1 0 1656 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_337
timestamp 1682952543
transform 1 0 1696 0 1 2170
box -9 -3 26 105
use FILL  FILL_1654
timestamp 1682952543
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1682952543
transform 1 0 1720 0 1 2170
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1682952543
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use FILL  FILL_1657
timestamp 1682952543
transform 1 0 1736 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4750
timestamp 1682952543
transform 1 0 1772 0 1 2175
box -3 -3 3 3
use M3_M2  M3_M2_4751
timestamp 1682952543
transform 1 0 1788 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_190
timestamp 1682952543
transform 1 0 1744 0 1 2170
box -8 -3 46 105
use FILL  FILL_1658
timestamp 1682952543
transform 1 0 1784 0 1 2170
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1682952543
transform 1 0 1792 0 1 2170
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1682952543
transform 1 0 1800 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_338
timestamp 1682952543
transform 1 0 1808 0 1 2170
box -9 -3 26 105
use FILL  FILL_1661
timestamp 1682952543
transform 1 0 1824 0 1 2170
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1682952543
transform 1 0 1832 0 1 2170
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1682952543
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_1664
timestamp 1682952543
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4752
timestamp 1682952543
transform 1 0 1868 0 1 2175
box -3 -3 3 3
use FILL  FILL_1665
timestamp 1682952543
transform 1 0 1856 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_191
timestamp 1682952543
transform 1 0 1864 0 1 2170
box -8 -3 46 105
use FILL  FILL_1666
timestamp 1682952543
transform 1 0 1904 0 1 2170
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1682952543
transform 1 0 1912 0 1 2170
box -8 -3 16 105
use FILL  FILL_1668
timestamp 1682952543
transform 1 0 1920 0 1 2170
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1682952543
transform 1 0 1928 0 1 2170
box -8 -3 16 105
use FILL  FILL_1670
timestamp 1682952543
transform 1 0 1936 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_192
timestamp 1682952543
transform 1 0 1944 0 1 2170
box -8 -3 46 105
use FILL  FILL_1671
timestamp 1682952543
transform 1 0 1984 0 1 2170
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1682952543
transform 1 0 1992 0 1 2170
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1682952543
transform 1 0 2000 0 1 2170
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1682952543
transform 1 0 2008 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_339
timestamp 1682952543
transform 1 0 2016 0 1 2170
box -9 -3 26 105
use FILL  FILL_1675
timestamp 1682952543
transform 1 0 2032 0 1 2170
box -8 -3 16 105
use FILL  FILL_1676
timestamp 1682952543
transform 1 0 2040 0 1 2170
box -8 -3 16 105
use FILL  FILL_1677
timestamp 1682952543
transform 1 0 2048 0 1 2170
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1682952543
transform 1 0 2056 0 1 2170
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1682952543
transform 1 0 2064 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_340
timestamp 1682952543
transform -1 0 2088 0 1 2170
box -9 -3 26 105
use FILL  FILL_1680
timestamp 1682952543
transform 1 0 2088 0 1 2170
box -8 -3 16 105
use FILL  FILL_1681
timestamp 1682952543
transform 1 0 2096 0 1 2170
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1682952543
transform 1 0 2104 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4753
timestamp 1682952543
transform 1 0 2124 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_193
timestamp 1682952543
transform 1 0 2112 0 1 2170
box -8 -3 46 105
use M3_M2  M3_M2_4754
timestamp 1682952543
transform 1 0 2164 0 1 2175
box -3 -3 3 3
use FILL  FILL_1686
timestamp 1682952543
transform 1 0 2152 0 1 2170
box -8 -3 16 105
use FILL  FILL_1688
timestamp 1682952543
transform 1 0 2160 0 1 2170
box -8 -3 16 105
use FILL  FILL_1690
timestamp 1682952543
transform 1 0 2168 0 1 2170
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1682952543
transform 1 0 2176 0 1 2170
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1682952543
transform 1 0 2184 0 1 2170
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1682952543
transform 1 0 2192 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_195
timestamp 1682952543
transform -1 0 2240 0 1 2170
box -8 -3 46 105
use FILL  FILL_1694
timestamp 1682952543
transform 1 0 2240 0 1 2170
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1682952543
transform 1 0 2248 0 1 2170
box -8 -3 16 105
use FILL  FILL_1696
timestamp 1682952543
transform 1 0 2256 0 1 2170
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1682952543
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use AND2X2  AND2X2_44
timestamp 1682952543
transform 1 0 2272 0 1 2170
box -8 -3 40 105
use M3_M2  M3_M2_4755
timestamp 1682952543
transform 1 0 2316 0 1 2175
box -3 -3 3 3
use FILL  FILL_1698
timestamp 1682952543
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1682952543
transform 1 0 2312 0 1 2170
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1682952543
transform 1 0 2320 0 1 2170
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1682952543
transform 1 0 2328 0 1 2170
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1682952543
transform 1 0 2336 0 1 2170
box -8 -3 16 105
use FILL  FILL_1703
timestamp 1682952543
transform 1 0 2344 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_196
timestamp 1682952543
transform 1 0 2352 0 1 2170
box -8 -3 46 105
use FILL  FILL_1704
timestamp 1682952543
transform 1 0 2392 0 1 2170
box -8 -3 16 105
use FILL  FILL_1705
timestamp 1682952543
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_1706
timestamp 1682952543
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use FILL  FILL_1707
timestamp 1682952543
transform 1 0 2416 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_342
timestamp 1682952543
transform 1 0 2424 0 1 2170
box -9 -3 26 105
use FILL  FILL_1708
timestamp 1682952543
transform 1 0 2440 0 1 2170
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1682952543
transform 1 0 2448 0 1 2170
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1682952543
transform 1 0 2456 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_307
timestamp 1682952543
transform -1 0 2560 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4756
timestamp 1682952543
transform 1 0 2572 0 1 2175
box -3 -3 3 3
use FILL  FILL_1719
timestamp 1682952543
transform 1 0 2560 0 1 2170
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1682952543
transform 1 0 2568 0 1 2170
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1682952543
transform 1 0 2576 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4757
timestamp 1682952543
transform 1 0 2612 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_346
timestamp 1682952543
transform 1 0 2584 0 1 2170
box -9 -3 26 105
use FILL  FILL_1731
timestamp 1682952543
transform 1 0 2600 0 1 2170
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1682952543
transform 1 0 2608 0 1 2170
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1682952543
transform 1 0 2616 0 1 2170
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1682952543
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1682952543
transform 1 0 2632 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4758
timestamp 1682952543
transform 1 0 2676 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_200
timestamp 1682952543
transform 1 0 2640 0 1 2170
box -8 -3 46 105
use FILL  FILL_1738
timestamp 1682952543
transform 1 0 2680 0 1 2170
box -8 -3 16 105
use FILL  FILL_1743
timestamp 1682952543
transform 1 0 2688 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4759
timestamp 1682952543
transform 1 0 2716 0 1 2175
box -3 -3 3 3
use FILL  FILL_1745
timestamp 1682952543
transform 1 0 2696 0 1 2170
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1682952543
transform 1 0 2704 0 1 2170
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1682952543
transform 1 0 2712 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4760
timestamp 1682952543
transform 1 0 2732 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_201
timestamp 1682952543
transform 1 0 2720 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_348
timestamp 1682952543
transform 1 0 2760 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_308
timestamp 1682952543
transform -1 0 2872 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4761
timestamp 1682952543
transform 1 0 2916 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_309
timestamp 1682952543
transform -1 0 2968 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4762
timestamp 1682952543
transform 1 0 2996 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_310
timestamp 1682952543
transform 1 0 2968 0 1 2170
box -8 -3 104 105
use FILL  FILL_1749
timestamp 1682952543
transform 1 0 3064 0 1 2170
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1682952543
transform 1 0 3072 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_67
timestamp 1682952543
transform 1 0 3080 0 1 2170
box -5 -3 28 105
use M3_M2  M3_M2_4763
timestamp 1682952543
transform 1 0 3140 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_311
timestamp 1682952543
transform 1 0 3104 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_351
timestamp 1682952543
transform 1 0 3200 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_312
timestamp 1682952543
transform 1 0 3216 0 1 2170
box -8 -3 104 105
use FILL  FILL_1772
timestamp 1682952543
transform 1 0 3312 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_352
timestamp 1682952543
transform 1 0 3320 0 1 2170
box -9 -3 26 105
use FILL  FILL_1773
timestamp 1682952543
transform 1 0 3336 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_27
timestamp 1682952543
transform -1 0 3376 0 1 2170
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_313
timestamp 1682952543
transform 1 0 3376 0 1 2170
box -8 -3 104 105
use NAND3X1  NAND3X1_28
timestamp 1682952543
transform -1 0 3504 0 1 2170
box -8 -3 40 105
use M3_M2  M3_M2_4764
timestamp 1682952543
transform 1 0 3532 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_314
timestamp 1682952543
transform -1 0 3600 0 1 2170
box -8 -3 104 105
use NAND3X1  NAND3X1_29
timestamp 1682952543
transform -1 0 3632 0 1 2170
box -8 -3 40 105
use NAND3X1  NAND3X1_30
timestamp 1682952543
transform -1 0 3664 0 1 2170
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_315
timestamp 1682952543
transform 1 0 3664 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4765
timestamp 1682952543
transform 1 0 3772 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_353
timestamp 1682952543
transform 1 0 3760 0 1 2170
box -9 -3 26 105
use M3_M2  M3_M2_4766
timestamp 1682952543
transform 1 0 3812 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_316
timestamp 1682952543
transform 1 0 3776 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_354
timestamp 1682952543
transform 1 0 3872 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_317
timestamp 1682952543
transform 1 0 3888 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4767
timestamp 1682952543
transform 1 0 4012 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_211
timestamp 1682952543
transform 1 0 3984 0 1 2170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_318
timestamp 1682952543
transform 1 0 4024 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4768
timestamp 1682952543
transform 1 0 4132 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_355
timestamp 1682952543
transform 1 0 4120 0 1 2170
box -9 -3 26 105
use FILL  FILL_1774
timestamp 1682952543
transform 1 0 4136 0 1 2170
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1682952543
transform 1 0 4144 0 1 2170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_39
timestamp 1682952543
transform 1 0 4177 0 1 2170
box -10 -3 10 3
use M3_M2  M3_M2_4868
timestamp 1682952543
transform 1 0 108 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4899
timestamp 1682952543
transform 1 0 116 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4843
timestamp 1682952543
transform 1 0 140 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4900
timestamp 1682952543
transform 1 0 140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4795
timestamp 1682952543
transform 1 0 148 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4898
timestamp 1682952543
transform 1 0 148 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4807
timestamp 1682952543
transform 1 0 164 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4796
timestamp 1682952543
transform 1 0 164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1682952543
transform 1 0 180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1682952543
transform 1 0 172 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4899
timestamp 1682952543
transform 1 0 172 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4798
timestamp 1682952543
transform 1 0 196 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4844
timestamp 1682952543
transform 1 0 204 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4902
timestamp 1682952543
transform 1 0 196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4903
timestamp 1682952543
transform 1 0 204 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4900
timestamp 1682952543
transform 1 0 196 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4950
timestamp 1682952543
transform 1 0 204 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4808
timestamp 1682952543
transform 1 0 220 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4769
timestamp 1682952543
transform 1 0 260 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_4799
timestamp 1682952543
transform 1 0 220 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4800
timestamp 1682952543
transform 1 0 236 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4845
timestamp 1682952543
transform 1 0 244 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4809
timestamp 1682952543
transform 1 0 268 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4801
timestamp 1682952543
transform 1 0 252 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4802
timestamp 1682952543
transform 1 0 268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4803
timestamp 1682952543
transform 1 0 284 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1682952543
transform 1 0 292 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4869
timestamp 1682952543
transform 1 0 220 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4904
timestamp 1682952543
transform 1 0 228 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1682952543
transform 1 0 244 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4870
timestamp 1682952543
transform 1 0 252 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4906
timestamp 1682952543
transform 1 0 260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1682952543
transform 1 0 276 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4871
timestamp 1682952543
transform 1 0 284 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4908
timestamp 1682952543
transform 1 0 292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4909
timestamp 1682952543
transform 1 0 300 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4901
timestamp 1682952543
transform 1 0 260 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4951
timestamp 1682952543
transform 1 0 228 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4952
timestamp 1682952543
transform 1 0 244 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4980
timestamp 1682952543
transform 1 0 292 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4953
timestamp 1682952543
transform 1 0 316 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_4805
timestamp 1682952543
transform 1 0 348 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4902
timestamp 1682952543
transform 1 0 348 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4810
timestamp 1682952543
transform 1 0 364 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4806
timestamp 1682952543
transform 1 0 364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4807
timestamp 1682952543
transform 1 0 380 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4811
timestamp 1682952543
transform 1 0 412 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4808
timestamp 1682952543
transform 1 0 396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4809
timestamp 1682952543
transform 1 0 412 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4793
timestamp 1682952543
transform 1 0 532 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4812
timestamp 1682952543
transform 1 0 516 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4813
timestamp 1682952543
transform 1 0 564 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4814
timestamp 1682952543
transform 1 0 604 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4810
timestamp 1682952543
transform 1 0 436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1682952543
transform 1 0 380 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1682952543
transform 1 0 388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4912
timestamp 1682952543
transform 1 0 404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1682952543
transform 1 0 420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1682952543
transform 1 0 460 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4954
timestamp 1682952543
transform 1 0 380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1682952543
transform 1 0 404 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1682952543
transform 1 0 484 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4811
timestamp 1682952543
transform 1 0 532 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4915
timestamp 1682952543
transform 1 0 516 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4916
timestamp 1682952543
transform 1 0 580 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4955
timestamp 1682952543
transform 1 0 460 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4981
timestamp 1682952543
transform 1 0 420 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1682952543
transform 1 0 444 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1682952543
transform 1 0 484 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4873
timestamp 1682952543
transform 1 0 604 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4904
timestamp 1682952543
transform 1 0 596 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4984
timestamp 1682952543
transform 1 0 540 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1682952543
transform 1 0 636 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4812
timestamp 1682952543
transform 1 0 628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1682952543
transform 1 0 636 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1682952543
transform 1 0 644 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4905
timestamp 1682952543
transform 1 0 636 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1682952543
transform 1 0 660 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4813
timestamp 1682952543
transform 1 0 684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4919
timestamp 1682952543
transform 1 0 668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1682952543
transform 1 0 684 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4956
timestamp 1682952543
transform 1 0 668 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1682952543
transform 1 0 700 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4960
timestamp 1682952543
transform 1 0 708 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4794
timestamp 1682952543
transform 1 0 732 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4795
timestamp 1682952543
transform 1 0 764 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_4814
timestamp 1682952543
transform 1 0 732 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1682952543
transform 1 0 756 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4874
timestamp 1682952543
transform 1 0 812 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4961
timestamp 1682952543
transform 1 0 748 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_4815
timestamp 1682952543
transform 1 0 828 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1682952543
transform 1 0 836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4791
timestamp 1682952543
transform 1 0 876 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4816
timestamp 1682952543
transform 1 0 868 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4846
timestamp 1682952543
transform 1 0 876 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4923
timestamp 1682952543
transform 1 0 868 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4875
timestamp 1682952543
transform 1 0 900 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4924
timestamp 1682952543
transform 1 0 908 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4906
timestamp 1682952543
transform 1 0 892 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5029
timestamp 1682952543
transform 1 0 900 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4907
timestamp 1682952543
transform 1 0 908 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4770
timestamp 1682952543
transform 1 0 940 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4847
timestamp 1682952543
transform 1 0 940 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1682952543
transform 1 0 956 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4818
timestamp 1682952543
transform 1 0 980 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4925
timestamp 1682952543
transform 1 0 980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4817
timestamp 1682952543
transform 1 0 996 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4848
timestamp 1682952543
transform 1 0 1020 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4926
timestamp 1682952543
transform 1 0 1004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4818
timestamp 1682952543
transform 1 0 1036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4819
timestamp 1682952543
transform 1 0 1052 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1682952543
transform 1 0 1052 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1682952543
transform 1 0 1068 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4819
timestamp 1682952543
transform 1 0 1100 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4820
timestamp 1682952543
transform 1 0 1100 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1682952543
transform 1 0 1124 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4821
timestamp 1682952543
transform 1 0 1156 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4877
timestamp 1682952543
transform 1 0 1180 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5031
timestamp 1682952543
transform 1 0 1164 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4962
timestamp 1682952543
transform 1 0 1172 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_4929
timestamp 1682952543
transform 1 0 1212 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4963
timestamp 1682952543
transform 1 0 1204 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_4930
timestamp 1682952543
transform 1 0 1228 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4964
timestamp 1682952543
transform 1 0 1220 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_4822
timestamp 1682952543
transform 1 0 1244 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4878
timestamp 1682952543
transform 1 0 1244 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4823
timestamp 1682952543
transform 1 0 1268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1682952543
transform 1 0 1260 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1682952543
transform 1 0 1276 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4908
timestamp 1682952543
transform 1 0 1260 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4965
timestamp 1682952543
transform 1 0 1292 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4909
timestamp 1682952543
transform 1 0 1308 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4985
timestamp 1682952543
transform 1 0 1316 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_4824
timestamp 1682952543
transform 1 0 1332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1682952543
transform 1 0 1364 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1682952543
transform 1 0 1356 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4879
timestamp 1682952543
transform 1 0 1364 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4934
timestamp 1682952543
transform 1 0 1372 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4910
timestamp 1682952543
transform 1 0 1372 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4826
timestamp 1682952543
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4771
timestamp 1682952543
transform 1 0 1428 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4772
timestamp 1682952543
transform 1 0 1508 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4820
timestamp 1682952543
transform 1 0 1492 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4827
timestamp 1682952543
transform 1 0 1492 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1682952543
transform 1 0 1412 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4936
timestamp 1682952543
transform 1 0 1468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1682952543
transform 1 0 1508 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4911
timestamp 1682952543
transform 1 0 1468 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1682952543
transform 1 0 1508 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1682952543
transform 1 0 1556 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_4828
timestamp 1682952543
transform 1 0 1556 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4880
timestamp 1682952543
transform 1 0 1556 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4938
timestamp 1682952543
transform 1 0 1564 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4913
timestamp 1682952543
transform 1 0 1580 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1682952543
transform 1 0 1588 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4774
timestamp 1682952543
transform 1 0 1604 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_4829
timestamp 1682952543
transform 1 0 1604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4830
timestamp 1682952543
transform 1 0 1612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1682952543
transform 1 0 1628 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4832
timestamp 1682952543
transform 1 0 1636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4939
timestamp 1682952543
transform 1 0 1596 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4986
timestamp 1682952543
transform 1 0 1596 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_4940
timestamp 1682952543
transform 1 0 1620 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4914
timestamp 1682952543
transform 1 0 1620 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4987
timestamp 1682952543
transform 1 0 1636 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4775
timestamp 1682952543
transform 1 0 1700 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1682952543
transform 1 0 1740 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4821
timestamp 1682952543
transform 1 0 1740 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4833
timestamp 1682952543
transform 1 0 1740 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1682952543
transform 1 0 1660 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1682952543
transform 1 0 1708 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4915
timestamp 1682952543
transform 1 0 1740 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4966
timestamp 1682952543
transform 1 0 1724 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4988
timestamp 1682952543
transform 1 0 1700 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1682952543
transform 1 0 1732 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1682952543
transform 1 0 1796 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4778
timestamp 1682952543
transform 1 0 1836 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1682952543
transform 1 0 1844 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1682952543
transform 1 0 1892 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4834
timestamp 1682952543
transform 1 0 1844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4835
timestamp 1682952543
transform 1 0 1860 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4836
timestamp 1682952543
transform 1 0 1876 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1682952543
transform 1 0 1892 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4838
timestamp 1682952543
transform 1 0 1900 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1682952543
transform 1 0 1764 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1682952543
transform 1 0 1820 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4882
timestamp 1682952543
transform 1 0 1860 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4945
timestamp 1682952543
transform 1 0 1868 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4946
timestamp 1682952543
transform 1 0 1884 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4916
timestamp 1682952543
transform 1 0 1772 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4917
timestamp 1682952543
transform 1 0 1844 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4967
timestamp 1682952543
transform 1 0 1796 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4779
timestamp 1682952543
transform 1 0 1964 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4780
timestamp 1682952543
transform 1 0 2004 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4824
timestamp 1682952543
transform 1 0 1916 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4849
timestamp 1682952543
transform 1 0 1908 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4839
timestamp 1682952543
transform 1 0 1996 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4947
timestamp 1682952543
transform 1 0 1908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1682952543
transform 1 0 1916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1682952543
transform 1 0 1948 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4918
timestamp 1682952543
transform 1 0 1908 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4919
timestamp 1682952543
transform 1 0 1948 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4968
timestamp 1682952543
transform 1 0 1996 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_4840
timestamp 1682952543
transform 1 0 2020 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4883
timestamp 1682952543
transform 1 0 2020 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4950
timestamp 1682952543
transform 1 0 2044 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4781
timestamp 1682952543
transform 1 0 2108 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4782
timestamp 1682952543
transform 1 0 2140 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1682952543
transform 1 0 2140 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4841
timestamp 1682952543
transform 1 0 2116 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4842
timestamp 1682952543
transform 1 0 2140 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4951
timestamp 1682952543
transform 1 0 2108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1682952543
transform 1 0 2116 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1682952543
transform 1 0 2132 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4920
timestamp 1682952543
transform 1 0 2044 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1682952543
transform 1 0 2100 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4969
timestamp 1682952543
transform 1 0 2068 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1682952543
transform 1 0 2132 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4970
timestamp 1682952543
transform 1 0 2116 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_4843
timestamp 1682952543
transform 1 0 2156 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4826
timestamp 1682952543
transform 1 0 2172 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4954
timestamp 1682952543
transform 1 0 2164 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4923
timestamp 1682952543
transform 1 0 2156 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4971
timestamp 1682952543
transform 1 0 2164 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4783
timestamp 1682952543
transform 1 0 2252 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4827
timestamp 1682952543
transform 1 0 2196 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4850
timestamp 1682952543
transform 1 0 2236 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4844
timestamp 1682952543
transform 1 0 2276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4955
timestamp 1682952543
transform 1 0 2188 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4956
timestamp 1682952543
transform 1 0 2196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1682952543
transform 1 0 2228 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4924
timestamp 1682952543
transform 1 0 2188 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4884
timestamp 1682952543
transform 1 0 2276 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4925
timestamp 1682952543
transform 1 0 2228 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4851
timestamp 1682952543
transform 1 0 2292 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4828
timestamp 1682952543
transform 1 0 2308 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4845
timestamp 1682952543
transform 1 0 2308 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1682952543
transform 1 0 2324 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4847
timestamp 1682952543
transform 1 0 2332 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4958
timestamp 1682952543
transform 1 0 2292 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4959
timestamp 1682952543
transform 1 0 2300 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4960
timestamp 1682952543
transform 1 0 2316 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1682952543
transform 1 0 2332 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1682952543
transform 1 0 2340 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4926
timestamp 1682952543
transform 1 0 2332 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4990
timestamp 1682952543
transform 1 0 2316 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4972
timestamp 1682952543
transform 1 0 2348 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1682952543
transform 1 0 2388 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1682952543
transform 1 0 2420 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4848
timestamp 1682952543
transform 1 0 2388 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4852
timestamp 1682952543
transform 1 0 2396 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4849
timestamp 1682952543
transform 1 0 2404 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4792
timestamp 1682952543
transform 1 0 2444 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1682952543
transform 1 0 2396 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4964
timestamp 1682952543
transform 1 0 2404 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4965
timestamp 1682952543
transform 1 0 2420 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4966
timestamp 1682952543
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4991
timestamp 1682952543
transform 1 0 2404 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4927
timestamp 1682952543
transform 1 0 2436 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1682952543
transform 1 0 2460 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_4967
timestamp 1682952543
transform 1 0 2468 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4784
timestamp 1682952543
transform 1 0 2492 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1682952543
transform 1 0 2484 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4850
timestamp 1682952543
transform 1 0 2484 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1682952543
transform 1 0 2492 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4885
timestamp 1682952543
transform 1 0 2484 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4968
timestamp 1682952543
transform 1 0 2492 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4797
timestamp 1682952543
transform 1 0 2516 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4853
timestamp 1682952543
transform 1 0 2548 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4969
timestamp 1682952543
transform 1 0 2532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4970
timestamp 1682952543
transform 1 0 2548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4971
timestamp 1682952543
transform 1 0 2556 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4928
timestamp 1682952543
transform 1 0 2556 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4992
timestamp 1682952543
transform 1 0 2548 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4929
timestamp 1682952543
transform 1 0 2572 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1682952543
transform 1 0 2612 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4799
timestamp 1682952543
transform 1 0 2628 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_4852
timestamp 1682952543
transform 1 0 2596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4853
timestamp 1682952543
transform 1 0 2604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1682952543
transform 1 0 2620 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1682952543
transform 1 0 2628 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4886
timestamp 1682952543
transform 1 0 2596 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4972
timestamp 1682952543
transform 1 0 2612 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4973
timestamp 1682952543
transform 1 0 2628 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4930
timestamp 1682952543
transform 1 0 2628 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4974
timestamp 1682952543
transform 1 0 2644 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4800
timestamp 1682952543
transform 1 0 2660 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_4793
timestamp 1682952543
transform 1 0 2684 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1682952543
transform 1 0 2692 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4785
timestamp 1682952543
transform 1 0 2708 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4801
timestamp 1682952543
transform 1 0 2724 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_4976
timestamp 1682952543
transform 1 0 2724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1682952543
transform 1 0 2732 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1682952543
transform 1 0 2748 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4973
timestamp 1682952543
transform 1 0 2740 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4993
timestamp 1682952543
transform 1 0 2748 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4786
timestamp 1682952543
transform 1 0 2780 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_4977
timestamp 1682952543
transform 1 0 2772 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1682952543
transform 1 0 2764 0 1 2105
box -2 -2 2 2
use M2_M1  M2_M1_4978
timestamp 1682952543
transform 1 0 2788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5033
timestamp 1682952543
transform 1 0 2788 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4832
timestamp 1682952543
transform 1 0 2828 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4857
timestamp 1682952543
transform 1 0 2828 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4833
timestamp 1682952543
transform 1 0 2860 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4979
timestamp 1682952543
transform 1 0 2820 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4980
timestamp 1682952543
transform 1 0 2836 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1682952543
transform 1 0 2852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4982
timestamp 1682952543
transform 1 0 2860 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4931
timestamp 1682952543
transform 1 0 2820 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4932
timestamp 1682952543
transform 1 0 2844 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4858
timestamp 1682952543
transform 1 0 2868 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4933
timestamp 1682952543
transform 1 0 2868 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4859
timestamp 1682952543
transform 1 0 2884 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4887
timestamp 1682952543
transform 1 0 2892 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1682952543
transform 1 0 2948 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_4860
timestamp 1682952543
transform 1 0 2924 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4983
timestamp 1682952543
transform 1 0 2916 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4854
timestamp 1682952543
transform 1 0 2932 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4861
timestamp 1682952543
transform 1 0 2940 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4855
timestamp 1682952543
transform 1 0 2948 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4984
timestamp 1682952543
transform 1 0 2932 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4974
timestamp 1682952543
transform 1 0 2932 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1682952543
transform 1 0 2972 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1682952543
transform 1 0 3020 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4862
timestamp 1682952543
transform 1 0 2988 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4863
timestamp 1682952543
transform 1 0 3004 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1682952543
transform 1 0 3020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1682952543
transform 1 0 2972 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4986
timestamp 1682952543
transform 1 0 2980 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4888
timestamp 1682952543
transform 1 0 3004 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4987
timestamp 1682952543
transform 1 0 3012 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4934
timestamp 1682952543
transform 1 0 3012 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4988
timestamp 1682952543
transform 1 0 3028 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4889
timestamp 1682952543
transform 1 0 3036 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4935
timestamp 1682952543
transform 1 0 3028 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1682952543
transform 1 0 3020 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_4865
timestamp 1682952543
transform 1 0 3060 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4890
timestamp 1682952543
transform 1 0 3060 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4866
timestamp 1682952543
transform 1 0 3092 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4788
timestamp 1682952543
transform 1 0 3132 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_4867
timestamp 1682952543
transform 1 0 3124 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1682952543
transform 1 0 3132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1682952543
transform 1 0 3148 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4857
timestamp 1682952543
transform 1 0 3156 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4870
timestamp 1682952543
transform 1 0 3164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1682952543
transform 1 0 3084 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1682952543
transform 1 0 3100 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1682952543
transform 1 0 3116 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4976
timestamp 1682952543
transform 1 0 3076 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4891
timestamp 1682952543
transform 1 0 3124 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4992
timestamp 1682952543
transform 1 0 3140 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1682952543
transform 1 0 3156 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4936
timestamp 1682952543
transform 1 0 3092 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4937
timestamp 1682952543
transform 1 0 3140 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4994
timestamp 1682952543
transform 1 0 3180 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1682952543
transform 1 0 3180 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_4794
timestamp 1682952543
transform 1 0 3204 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_4858
timestamp 1682952543
transform 1 0 3204 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4835
timestamp 1682952543
transform 1 0 3252 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4871
timestamp 1682952543
transform 1 0 3236 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4872
timestamp 1682952543
transform 1 0 3252 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1682952543
transform 1 0 3220 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5035
timestamp 1682952543
transform 1 0 3204 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1682952543
transform 1 0 3188 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4957
timestamp 1682952543
transform 1 0 3196 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4977
timestamp 1682952543
transform 1 0 3188 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1682952543
transform 1 0 3212 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4892
timestamp 1682952543
transform 1 0 3236 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_4996
timestamp 1682952543
transform 1 0 3244 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4939
timestamp 1682952543
transform 1 0 3228 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4859
timestamp 1682952543
transform 1 0 3260 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4873
timestamp 1682952543
transform 1 0 3268 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1682952543
transform 1 0 3260 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4940
timestamp 1682952543
transform 1 0 3260 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1682952543
transform 1 0 3300 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4874
timestamp 1682952543
transform 1 0 3300 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4860
timestamp 1682952543
transform 1 0 3308 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4875
timestamp 1682952543
transform 1 0 3316 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4998
timestamp 1682952543
transform 1 0 3308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4999
timestamp 1682952543
transform 1 0 3324 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4893
timestamp 1682952543
transform 1 0 3332 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1682952543
transform 1 0 3388 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4876
timestamp 1682952543
transform 1 0 3436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5000
timestamp 1682952543
transform 1 0 3388 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1682952543
transform 1 0 3468 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4861
timestamp 1682952543
transform 1 0 3484 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4878
timestamp 1682952543
transform 1 0 3492 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4862
timestamp 1682952543
transform 1 0 3500 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4879
timestamp 1682952543
transform 1 0 3508 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5001
timestamp 1682952543
transform 1 0 3484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1682952543
transform 1 0 3500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1682952543
transform 1 0 3516 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4941
timestamp 1682952543
transform 1 0 3492 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4942
timestamp 1682952543
transform 1 0 3516 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5004
timestamp 1682952543
transform 1 0 3540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5005
timestamp 1682952543
transform 1 0 3548 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4978
timestamp 1682952543
transform 1 0 3548 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4863
timestamp 1682952543
transform 1 0 3564 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5036
timestamp 1682952543
transform 1 0 3564 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4789
timestamp 1682952543
transform 1 0 3572 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5006
timestamp 1682952543
transform 1 0 3572 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4802
timestamp 1682952543
transform 1 0 3604 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1682952543
transform 1 0 3612 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5007
timestamp 1682952543
transform 1 0 3612 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4894
timestamp 1682952543
transform 1 0 3620 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5037
timestamp 1682952543
transform 1 0 3620 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1682952543
transform 1 0 3604 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4895
timestamp 1682952543
transform 1 0 3636 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4803
timestamp 1682952543
transform 1 0 3684 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4804
timestamp 1682952543
transform 1 0 3716 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4838
timestamp 1682952543
transform 1 0 3716 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4880
timestamp 1682952543
transform 1 0 3684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1682952543
transform 1 0 3700 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1682952543
transform 1 0 3716 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1682952543
transform 1 0 3668 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5009
timestamp 1682952543
transform 1 0 3684 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5010
timestamp 1682952543
transform 1 0 3708 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1682952543
transform 1 0 3652 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4896
timestamp 1682952543
transform 1 0 3716 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5011
timestamp 1682952543
transform 1 0 3724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5039
timestamp 1682952543
transform 1 0 3676 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4943
timestamp 1682952543
transform 1 0 3684 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1682952543
transform 1 0 3708 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5045
timestamp 1682952543
transform 1 0 3660 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4958
timestamp 1682952543
transform 1 0 3668 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4994
timestamp 1682952543
transform 1 0 3660 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4995
timestamp 1682952543
transform 1 0 3684 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4805
timestamp 1682952543
transform 1 0 3788 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_4883
timestamp 1682952543
transform 1 0 3772 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1682952543
transform 1 0 3780 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4865
timestamp 1682952543
transform 1 0 3788 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4839
timestamp 1682952543
transform 1 0 3820 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4885
timestamp 1682952543
transform 1 0 3812 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4886
timestamp 1682952543
transform 1 0 3820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1682952543
transform 1 0 3836 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1682952543
transform 1 0 3852 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4866
timestamp 1682952543
transform 1 0 3860 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4889
timestamp 1682952543
transform 1 0 3868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1682952543
transform 1 0 3884 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5012
timestamp 1682952543
transform 1 0 3756 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1682952543
transform 1 0 3772 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5014
timestamp 1682952543
transform 1 0 3788 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5015
timestamp 1682952543
transform 1 0 3812 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5016
timestamp 1682952543
transform 1 0 3828 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5017
timestamp 1682952543
transform 1 0 3844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5018
timestamp 1682952543
transform 1 0 3852 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5019
timestamp 1682952543
transform 1 0 3876 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1682952543
transform 1 0 3740 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5041
timestamp 1682952543
transform 1 0 3756 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4996
timestamp 1682952543
transform 1 0 3724 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5046
timestamp 1682952543
transform 1 0 3748 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4945
timestamp 1682952543
transform 1 0 3780 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4997
timestamp 1682952543
transform 1 0 3772 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1682952543
transform 1 0 3836 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1682952543
transform 1 0 3828 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4897
timestamp 1682952543
transform 1 0 3884 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5020
timestamp 1682952543
transform 1 0 3892 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4947
timestamp 1682952543
transform 1 0 3876 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4998
timestamp 1682952543
transform 1 0 3844 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4806
timestamp 1682952543
transform 1 0 3900 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4979
timestamp 1682952543
transform 1 0 3892 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4790
timestamp 1682952543
transform 1 0 3948 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4840
timestamp 1682952543
transform 1 0 3940 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4891
timestamp 1682952543
transform 1 0 3916 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4867
timestamp 1682952543
transform 1 0 3924 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_4892
timestamp 1682952543
transform 1 0 3932 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1682952543
transform 1 0 3948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1682952543
transform 1 0 3916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5022
timestamp 1682952543
transform 1 0 3940 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4948
timestamp 1682952543
transform 1 0 3916 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5023
timestamp 1682952543
transform 1 0 3956 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1682952543
transform 1 0 3980 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1682952543
transform 1 0 3980 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4949
timestamp 1682952543
transform 1 0 3980 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_4895
timestamp 1682952543
transform 1 0 4004 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5025
timestamp 1682952543
transform 1 0 3996 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4791
timestamp 1682952543
transform 1 0 4020 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4792
timestamp 1682952543
transform 1 0 4044 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4841
timestamp 1682952543
transform 1 0 4028 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4896
timestamp 1682952543
transform 1 0 4028 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1682952543
transform 1 0 4044 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5026
timestamp 1682952543
transform 1 0 4036 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4842
timestamp 1682952543
transform 1 0 4092 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_4898
timestamp 1682952543
transform 1 0 4068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5027
timestamp 1682952543
transform 1 0 4092 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5028
timestamp 1682952543
transform 1 0 4148 0 1 2125
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_40
timestamp 1682952543
transform 1 0 24 0 1 2070
box -10 -3 10 3
use FILL  FILL_1520
timestamp 1682952543
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1682952543
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1682952543
transform 1 0 88 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1682952543
transform 1 0 96 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1682952543
transform 1 0 104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1682952543
transform 1 0 112 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_325
timestamp 1682952543
transform -1 0 136 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1526
timestamp 1682952543
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1527
timestamp 1682952543
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_178
timestamp 1682952543
transform -1 0 192 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1528
timestamp 1682952543
transform 1 0 192 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_326
timestamp 1682952543
transform 1 0 200 0 -1 2170
box -9 -3 26 105
use OAI22X1  OAI22X1_204
timestamp 1682952543
transform -1 0 256 0 -1 2170
box -8 -3 46 105
use AOI22X1  AOI22X1_179
timestamp 1682952543
transform 1 0 256 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_327
timestamp 1682952543
transform 1 0 296 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1529
timestamp 1682952543
transform 1 0 312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1682952543
transform 1 0 320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1682952543
transform 1 0 328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1682952543
transform 1 0 336 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_328
timestamp 1682952543
transform 1 0 344 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1533
timestamp 1682952543
transform 1 0 360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1534
timestamp 1682952543
transform 1 0 368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1682952543
transform 1 0 376 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_181
timestamp 1682952543
transform 1 0 384 0 -1 2170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_294
timestamp 1682952543
transform 1 0 424 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_295
timestamp 1682952543
transform 1 0 520 0 -1 2170
box -8 -3 104 105
use FILL  FILL_1546
timestamp 1682952543
transform 1 0 616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1682952543
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1682952543
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1551
timestamp 1682952543
transform 1 0 640 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_183
timestamp 1682952543
transform 1 0 648 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1552
timestamp 1682952543
transform 1 0 688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1682952543
transform 1 0 696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1682952543
transform 1 0 704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1558
timestamp 1682952543
transform 1 0 712 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_296
timestamp 1682952543
transform 1 0 720 0 -1 2170
box -8 -3 104 105
use FILL  FILL_1567
timestamp 1682952543
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1682952543
transform 1 0 824 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_65
timestamp 1682952543
transform 1 0 832 0 -1 2170
box -8 -3 34 105
use FILL  FILL_1572
timestamp 1682952543
transform 1 0 864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1682952543
transform 1 0 872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1574
timestamp 1682952543
transform 1 0 880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1682952543
transform 1 0 888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1682952543
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1682952543
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_59
timestamp 1682952543
transform 1 0 912 0 -1 2170
box -8 -3 32 105
use FILL  FILL_1585
timestamp 1682952543
transform 1 0 936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1682952543
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1587
timestamp 1682952543
transform 1 0 952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1588
timestamp 1682952543
transform 1 0 960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1589
timestamp 1682952543
transform 1 0 968 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4999
timestamp 1682952543
transform 1 0 988 0 1 2075
box -3 -3 3 3
use FILL  FILL_1590
timestamp 1682952543
transform 1 0 976 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_186
timestamp 1682952543
transform 1 0 984 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1596
timestamp 1682952543
transform 1 0 1024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1682952543
transform 1 0 1032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1682952543
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1604
timestamp 1682952543
transform 1 0 1048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1682952543
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1682952543
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_66
timestamp 1682952543
transform 1 0 1072 0 -1 2170
box -8 -3 34 105
use FILL  FILL_1607
timestamp 1682952543
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1608
timestamp 1682952543
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1682952543
transform 1 0 1120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1682952543
transform 1 0 1128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1682952543
transform 1 0 1136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1682952543
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1613
timestamp 1682952543
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_67
timestamp 1682952543
transform -1 0 1192 0 -1 2170
box -8 -3 34 105
use FILL  FILL_1614
timestamp 1682952543
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1682952543
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1682952543
transform 1 0 1208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1682952543
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1682952543
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1624
timestamp 1682952543
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1682952543
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_206
timestamp 1682952543
transform 1 0 1248 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1631
timestamp 1682952543
transform 1 0 1288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1682952543
transform 1 0 1296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1682952543
transform 1 0 1304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1682952543
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1682952543
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1682952543
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1682952543
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_207
timestamp 1682952543
transform -1 0 1384 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1638
timestamp 1682952543
transform 1 0 1384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1682952543
transform 1 0 1392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1682952543
transform 1 0 1400 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_301
timestamp 1682952543
transform -1 0 1504 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_335
timestamp 1682952543
transform -1 0 1520 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1641
timestamp 1682952543
transform 1 0 1520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1682952543
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1643
timestamp 1682952543
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1682952543
transform 1 0 1544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1682952543
transform 1 0 1552 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_336
timestamp 1682952543
transform -1 0 1576 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1646
timestamp 1682952543
transform 1 0 1576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1682952543
transform 1 0 1584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1651
timestamp 1682952543
transform 1 0 1592 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_188
timestamp 1682952543
transform -1 0 1640 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1652
timestamp 1682952543
transform 1 0 1640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1682952543
transform 1 0 1648 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_302
timestamp 1682952543
transform -1 0 1752 0 -1 2170
box -8 -3 104 105
use FILL  FILL_1684
timestamp 1682952543
transform 1 0 1752 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_303
timestamp 1682952543
transform -1 0 1856 0 -1 2170
box -8 -3 104 105
use OAI22X1  OAI22X1_208
timestamp 1682952543
transform 1 0 1856 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_341
timestamp 1682952543
transform 1 0 1896 0 -1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_304
timestamp 1682952543
transform -1 0 2008 0 -1 2170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_305
timestamp 1682952543
transform 1 0 2008 0 -1 2170
box -8 -3 104 105
use FILL  FILL_1685
timestamp 1682952543
transform 1 0 2104 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_194
timestamp 1682952543
transform 1 0 2112 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1687
timestamp 1682952543
transform 1 0 2152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1682952543
transform 1 0 2160 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_343
timestamp 1682952543
transform 1 0 2168 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1709
timestamp 1682952543
transform 1 0 2184 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_306
timestamp 1682952543
transform -1 0 2288 0 -1 2170
box -8 -3 104 105
use FILL  FILL_1710
timestamp 1682952543
transform 1 0 2288 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_197
timestamp 1682952543
transform 1 0 2296 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_344
timestamp 1682952543
transform 1 0 2336 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1711
timestamp 1682952543
transform 1 0 2352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1682952543
transform 1 0 2360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1682952543
transform 1 0 2368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1714
timestamp 1682952543
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_345
timestamp 1682952543
transform 1 0 2384 0 -1 2170
box -9 -3 26 105
use AOI22X1  AOI22X1_198
timestamp 1682952543
transform 1 0 2400 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1715
timestamp 1682952543
transform 1 0 2440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1717
timestamp 1682952543
transform 1 0 2448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1682952543
transform 1 0 2456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1682952543
transform 1 0 2464 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_60
timestamp 1682952543
transform 1 0 2472 0 -1 2170
box -8 -3 32 105
use FILL  FILL_1722
timestamp 1682952543
transform 1 0 2496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1682952543
transform 1 0 2504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1682952543
transform 1 0 2512 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_45
timestamp 1682952543
transform 1 0 2520 0 -1 2170
box -8 -3 40 105
use FILL  FILL_1725
timestamp 1682952543
transform 1 0 2552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1682952543
transform 1 0 2560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1682952543
transform 1 0 2568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1730
timestamp 1682952543
transform 1 0 2576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1736
timestamp 1682952543
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_199
timestamp 1682952543
transform -1 0 2632 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1737
timestamp 1682952543
transform 1 0 2632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1739
timestamp 1682952543
transform 1 0 2640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1740
timestamp 1682952543
transform 1 0 2648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1682952543
transform 1 0 2656 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_347
timestamp 1682952543
transform 1 0 2664 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1742
timestamp 1682952543
transform 1 0 2680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1682952543
transform 1 0 2688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1746
timestamp 1682952543
transform 1 0 2696 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_61
timestamp 1682952543
transform 1 0 2704 0 -1 2170
box -8 -3 32 105
use FILL  FILL_1750
timestamp 1682952543
transform 1 0 2728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1682952543
transform 1 0 2736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1682952543
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_26
timestamp 1682952543
transform -1 0 2784 0 -1 2170
box -8 -3 40 105
use FILL  FILL_1753
timestamp 1682952543
transform 1 0 2784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1754
timestamp 1682952543
transform 1 0 2792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1755
timestamp 1682952543
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1682952543
transform 1 0 2808 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_202
timestamp 1682952543
transform 1 0 2816 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1757
timestamp 1682952543
transform 1 0 2856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1682952543
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1682952543
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1682952543
transform 1 0 2880 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_349
timestamp 1682952543
transform 1 0 2888 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1761
timestamp 1682952543
transform 1 0 2904 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1682952543
transform 1 0 2912 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5000
timestamp 1682952543
transform 1 0 2932 0 1 2075
box -3 -3 3 3
use OAI22X1  OAI22X1_209
timestamp 1682952543
transform -1 0 2960 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1763
timestamp 1682952543
transform 1 0 2960 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5001
timestamp 1682952543
transform 1 0 2980 0 1 2075
box -3 -3 3 3
use FILL  FILL_1764
timestamp 1682952543
transform 1 0 2968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1765
timestamp 1682952543
transform 1 0 2976 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_210
timestamp 1682952543
transform 1 0 2984 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1766
timestamp 1682952543
transform 1 0 3024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1682952543
transform 1 0 3032 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_350
timestamp 1682952543
transform -1 0 3056 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1768
timestamp 1682952543
transform 1 0 3056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1682952543
transform 1 0 3064 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1771
timestamp 1682952543
transform 1 0 3072 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_203
timestamp 1682952543
transform 1 0 3080 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1776
timestamp 1682952543
transform 1 0 3120 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_212
timestamp 1682952543
transform -1 0 3168 0 -1 2170
box -8 -3 46 105
use NAND3X1  NAND3X1_31
timestamp 1682952543
transform 1 0 3168 0 -1 2170
box -8 -3 40 105
use FILL  FILL_1777
timestamp 1682952543
transform 1 0 3200 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_5002
timestamp 1682952543
transform 1 0 3220 0 1 2075
box -3 -3 3 3
use FILL  FILL_1778
timestamp 1682952543
transform 1 0 3208 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_213
timestamp 1682952543
transform 1 0 3216 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1779
timestamp 1682952543
transform 1 0 3256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1682952543
transform 1 0 3264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1682952543
transform 1 0 3272 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_214
timestamp 1682952543
transform 1 0 3280 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_356
timestamp 1682952543
transform -1 0 3336 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1782
timestamp 1682952543
transform 1 0 3336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1682952543
transform 1 0 3344 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_319
timestamp 1682952543
transform -1 0 3448 0 -1 2170
box -8 -3 104 105
use FILL  FILL_1784
timestamp 1682952543
transform 1 0 3448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1682952543
transform 1 0 3456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1786
timestamp 1682952543
transform 1 0 3464 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_357
timestamp 1682952543
transform 1 0 3472 0 -1 2170
box -9 -3 26 105
use OAI22X1  OAI22X1_215
timestamp 1682952543
transform -1 0 3528 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1787
timestamp 1682952543
transform 1 0 3528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1682952543
transform 1 0 3536 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_358
timestamp 1682952543
transform -1 0 3560 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1789
timestamp 1682952543
transform 1 0 3560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1682952543
transform 1 0 3568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1791
timestamp 1682952543
transform 1 0 3576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1792
timestamp 1682952543
transform 1 0 3584 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_32
timestamp 1682952543
transform -1 0 3624 0 -1 2170
box -8 -3 40 105
use FILL  FILL_1793
timestamp 1682952543
transform 1 0 3624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1682952543
transform 1 0 3632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1682952543
transform 1 0 3640 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_33
timestamp 1682952543
transform -1 0 3680 0 -1 2170
box -8 -3 40 105
use OAI22X1  OAI22X1_216
timestamp 1682952543
transform 1 0 3680 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_359
timestamp 1682952543
transform 1 0 3720 0 -1 2170
box -9 -3 26 105
use NAND3X1  NAND3X1_34
timestamp 1682952543
transform -1 0 3768 0 -1 2170
box -8 -3 40 105
use AOI22X1  AOI22X1_204
timestamp 1682952543
transform -1 0 3808 0 -1 2170
box -8 -3 46 105
use M3_M2  M3_M2_5003
timestamp 1682952543
transform 1 0 3852 0 1 2075
box -3 -3 3 3
use AOI22X1  AOI22X1_205
timestamp 1682952543
transform 1 0 3808 0 -1 2170
box -8 -3 46 105
use OAI22X1  OAI22X1_217
timestamp 1682952543
transform 1 0 3848 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1796
timestamp 1682952543
transform 1 0 3888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1682952543
transform 1 0 3896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1682952543
transform 1 0 3904 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_218
timestamp 1682952543
transform 1 0 3912 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1799
timestamp 1682952543
transform 1 0 3952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1682952543
transform 1 0 3960 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_360
timestamp 1682952543
transform -1 0 3984 0 -1 2170
box -9 -3 26 105
use FILL  FILL_1801
timestamp 1682952543
transform 1 0 3984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1682952543
transform 1 0 3992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_1803
timestamp 1682952543
transform 1 0 4000 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_219
timestamp 1682952543
transform 1 0 4008 0 -1 2170
box -8 -3 46 105
use FILL  FILL_1804
timestamp 1682952543
transform 1 0 4048 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_320
timestamp 1682952543
transform 1 0 4056 0 -1 2170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_41
timestamp 1682952543
transform 1 0 4201 0 1 2070
box -10 -3 10 3
use M3_M2  M3_M2_5057
timestamp 1682952543
transform 1 0 116 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1682952543
transform 1 0 172 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5066
timestamp 1682952543
transform 1 0 116 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5067
timestamp 1682952543
transform 1 0 164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1682952543
transform 1 0 172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5174
timestamp 1682952543
transform 1 0 84 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5138
timestamp 1682952543
transform 1 0 164 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5034
timestamp 1682952543
transform 1 0 196 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5059
timestamp 1682952543
transform 1 0 188 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5060
timestamp 1682952543
transform 1 0 212 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5069
timestamp 1682952543
transform 1 0 196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5070
timestamp 1682952543
transform 1 0 212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5071
timestamp 1682952543
transform 1 0 228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5175
timestamp 1682952543
transform 1 0 188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5176
timestamp 1682952543
transform 1 0 196 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1682952543
transform 1 0 220 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5170
timestamp 1682952543
transform 1 0 180 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1682952543
transform 1 0 220 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1682952543
transform 1 0 284 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5072
timestamp 1682952543
transform 1 0 244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1682952543
transform 1 0 300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1682952543
transform 1 0 324 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5171
timestamp 1682952543
transform 1 0 236 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5179
timestamp 1682952543
transform 1 0 340 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5140
timestamp 1682952543
transform 1 0 340 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1682952543
transform 1 0 388 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5074
timestamp 1682952543
transform 1 0 364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1682952543
transform 1 0 380 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5180
timestamp 1682952543
transform 1 0 372 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5172
timestamp 1682952543
transform 1 0 372 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5076
timestamp 1682952543
transform 1 0 396 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1682952543
transform 1 0 412 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1682952543
transform 1 0 428 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5037
timestamp 1682952543
transform 1 0 460 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5078
timestamp 1682952543
transform 1 0 452 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5114
timestamp 1682952543
transform 1 0 436 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5182
timestamp 1682952543
transform 1 0 460 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5183
timestamp 1682952543
transform 1 0 468 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5079
timestamp 1682952543
transform 1 0 484 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5038
timestamp 1682952543
transform 1 0 524 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5061
timestamp 1682952543
transform 1 0 516 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5062
timestamp 1682952543
transform 1 0 556 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5080
timestamp 1682952543
transform 1 0 516 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5081
timestamp 1682952543
transform 1 0 524 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1682952543
transform 1 0 556 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1682952543
transform 1 0 604 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5275
timestamp 1682952543
transform 1 0 628 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5173
timestamp 1682952543
transform 1 0 628 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5185
timestamp 1682952543
transform 1 0 644 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5174
timestamp 1682952543
transform 1 0 652 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5083
timestamp 1682952543
transform 1 0 692 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5063
timestamp 1682952543
transform 1 0 716 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5084
timestamp 1682952543
transform 1 0 708 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5186
timestamp 1682952543
transform 1 0 700 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5141
timestamp 1682952543
transform 1 0 692 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5175
timestamp 1682952543
transform 1 0 684 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5187
timestamp 1682952543
transform 1 0 724 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5142
timestamp 1682952543
transform 1 0 724 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5085
timestamp 1682952543
transform 1 0 740 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1682952543
transform 1 0 756 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1682952543
transform 1 0 748 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5143
timestamp 1682952543
transform 1 0 756 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1682952543
transform 1 0 788 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5064
timestamp 1682952543
transform 1 0 804 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5086
timestamp 1682952543
transform 1 0 788 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5087
timestamp 1682952543
transform 1 0 804 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5115
timestamp 1682952543
transform 1 0 772 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5189
timestamp 1682952543
transform 1 0 796 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5190
timestamp 1682952543
transform 1 0 804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1682952543
transform 1 0 876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1682952543
transform 1 0 892 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5191
timestamp 1682952543
transform 1 0 868 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5176
timestamp 1682952543
transform 1 0 876 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1682952543
transform 1 0 900 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5192
timestamp 1682952543
transform 1 0 924 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1682952543
transform 1 0 988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5193
timestamp 1682952543
transform 1 0 972 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1682952543
transform 1 0 980 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5195
timestamp 1682952543
transform 1 0 1012 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5100
timestamp 1682952543
transform 1 0 1020 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5196
timestamp 1682952543
transform 1 0 1020 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5004
timestamp 1682952543
transform 1 0 1068 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5091
timestamp 1682952543
transform 1 0 1076 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5144
timestamp 1682952543
transform 1 0 1068 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1682952543
transform 1 0 1084 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5054
timestamp 1682952543
transform 1 0 1084 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5092
timestamp 1682952543
transform 1 0 1100 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5101
timestamp 1682952543
transform 1 0 1132 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5197
timestamp 1682952543
transform 1 0 1116 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5198
timestamp 1682952543
transform 1 0 1124 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5145
timestamp 1682952543
transform 1 0 1124 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1682952543
transform 1 0 1164 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5055
timestamp 1682952543
transform 1 0 1164 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5093
timestamp 1682952543
transform 1 0 1204 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5094
timestamp 1682952543
transform 1 0 1212 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5146
timestamp 1682952543
transform 1 0 1204 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1682952543
transform 1 0 1228 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1682952543
transform 1 0 1268 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5065
timestamp 1682952543
transform 1 0 1292 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5066
timestamp 1682952543
transform 1 0 1316 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5095
timestamp 1682952543
transform 1 0 1292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1682952543
transform 1 0 1308 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1682952543
transform 1 0 1316 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5199
timestamp 1682952543
transform 1 0 1276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5200
timestamp 1682952543
transform 1 0 1284 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5201
timestamp 1682952543
transform 1 0 1300 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5117
timestamp 1682952543
transform 1 0 1308 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1682952543
transform 1 0 1284 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5102
timestamp 1682952543
transform 1 0 1324 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5179
timestamp 1682952543
transform 1 0 1332 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5202
timestamp 1682952543
transform 1 0 1356 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5017
timestamp 1682952543
transform 1 0 1484 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5098
timestamp 1682952543
transform 1 0 1412 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5103
timestamp 1682952543
transform 1 0 1476 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5118
timestamp 1682952543
transform 1 0 1412 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5203
timestamp 1682952543
transform 1 0 1460 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1682952543
transform 1 0 1476 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5099
timestamp 1682952543
transform 1 0 1500 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5180
timestamp 1682952543
transform 1 0 1492 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5018
timestamp 1682952543
transform 1 0 1540 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5041
timestamp 1682952543
transform 1 0 1532 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5042
timestamp 1682952543
transform 1 0 1580 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1682952543
transform 1 0 1644 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5067
timestamp 1682952543
transform 1 0 1628 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5100
timestamp 1682952543
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5101
timestamp 1682952543
transform 1 0 1612 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5102
timestamp 1682952543
transform 1 0 1628 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1682952543
transform 1 0 1644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1682952543
transform 1 0 1516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5206
timestamp 1682952543
transform 1 0 1532 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5119
timestamp 1682952543
transform 1 0 1564 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5120
timestamp 1682952543
transform 1 0 1580 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5207
timestamp 1682952543
transform 1 0 1620 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5208
timestamp 1682952543
transform 1 0 1636 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5121
timestamp 1682952543
transform 1 0 1644 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5209
timestamp 1682952543
transform 1 0 1652 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5210
timestamp 1682952543
transform 1 0 1660 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5181
timestamp 1682952543
transform 1 0 1532 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1682952543
transform 1 0 1580 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1682952543
transform 1 0 1612 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5276
timestamp 1682952543
transform 1 0 1660 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5044
timestamp 1682952543
transform 1 0 1676 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5277
timestamp 1682952543
transform 1 0 1676 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5068
timestamp 1682952543
transform 1 0 1692 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5104
timestamp 1682952543
transform 1 0 1692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1682952543
transform 1 0 1708 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5211
timestamp 1682952543
transform 1 0 1700 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5122
timestamp 1682952543
transform 1 0 1708 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5106
timestamp 1682952543
transform 1 0 1724 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5212
timestamp 1682952543
transform 1 0 1716 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5123
timestamp 1682952543
transform 1 0 1756 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5213
timestamp 1682952543
transform 1 0 1764 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5214
timestamp 1682952543
transform 1 0 1772 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5045
timestamp 1682952543
transform 1 0 1796 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5107
timestamp 1682952543
transform 1 0 1796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1682952543
transform 1 0 1812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5215
timestamp 1682952543
transform 1 0 1804 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1682952543
transform 1 0 1820 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1682952543
transform 1 0 1828 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5124
timestamp 1682952543
transform 1 0 1844 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5005
timestamp 1682952543
transform 1 0 1908 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5046
timestamp 1682952543
transform 1 0 1884 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5047
timestamp 1682952543
transform 1 0 1900 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5069
timestamp 1682952543
transform 1 0 1876 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5109
timestamp 1682952543
transform 1 0 1868 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1682952543
transform 1 0 1900 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1682952543
transform 1 0 1892 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1682952543
transform 1 0 1916 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5147
timestamp 1682952543
transform 1 0 1916 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5184
timestamp 1682952543
transform 1 0 1916 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5219
timestamp 1682952543
transform 1 0 1932 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5104
timestamp 1682952543
transform 1 0 1948 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5047
timestamp 1682952543
transform 1 0 1996 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1682952543
transform 1 0 1988 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1682952543
transform 1 0 1980 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5185
timestamp 1682952543
transform 1 0 1964 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5070
timestamp 1682952543
transform 1 0 2036 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5220
timestamp 1682952543
transform 1 0 2044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1682952543
transform 1 0 2060 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5148
timestamp 1682952543
transform 1 0 2060 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5112
timestamp 1682952543
transform 1 0 2084 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5222
timestamp 1682952543
transform 1 0 2092 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5048
timestamp 1682952543
transform 1 0 2124 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5071
timestamp 1682952543
transform 1 0 2108 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5072
timestamp 1682952543
transform 1 0 2140 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5113
timestamp 1682952543
transform 1 0 2116 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5105
timestamp 1682952543
transform 1 0 2124 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5114
timestamp 1682952543
transform 1 0 2132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5223
timestamp 1682952543
transform 1 0 2124 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5125
timestamp 1682952543
transform 1 0 2132 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5224
timestamp 1682952543
transform 1 0 2140 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5073
timestamp 1682952543
transform 1 0 2156 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5186
timestamp 1682952543
transform 1 0 2156 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5049
timestamp 1682952543
transform 1 0 2196 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5074
timestamp 1682952543
transform 1 0 2180 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5115
timestamp 1682952543
transform 1 0 2180 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1682952543
transform 1 0 2196 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5225
timestamp 1682952543
transform 1 0 2172 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5126
timestamp 1682952543
transform 1 0 2180 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5226
timestamp 1682952543
transform 1 0 2188 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1682952543
transform 1 0 2204 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1682952543
transform 1 0 2212 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5187
timestamp 1682952543
transform 1 0 2180 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5050
timestamp 1682952543
transform 1 0 2236 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5075
timestamp 1682952543
transform 1 0 2244 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5076
timestamp 1682952543
transform 1 0 2260 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5117
timestamp 1682952543
transform 1 0 2228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1682952543
transform 1 0 2244 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5127
timestamp 1682952543
transform 1 0 2228 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5229
timestamp 1682952543
transform 1 0 2236 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5128
timestamp 1682952543
transform 1 0 2244 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5006
timestamp 1682952543
transform 1 0 2380 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5007
timestamp 1682952543
transform 1 0 2420 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5077
timestamp 1682952543
transform 1 0 2284 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5078
timestamp 1682952543
transform 1 0 2324 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1682952543
transform 1 0 2268 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5119
timestamp 1682952543
transform 1 0 2284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1682952543
transform 1 0 2340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5230
timestamp 1682952543
transform 1 0 2260 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1682952543
transform 1 0 2268 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5232
timestamp 1682952543
transform 1 0 2276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5233
timestamp 1682952543
transform 1 0 2364 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5278
timestamp 1682952543
transform 1 0 2260 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5188
timestamp 1682952543
transform 1 0 2236 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1682952543
transform 1 0 2260 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5149
timestamp 1682952543
transform 1 0 2364 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5019
timestamp 1682952543
transform 1 0 2476 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5020
timestamp 1682952543
transform 1 0 2492 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1682952543
transform 1 0 2500 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5121
timestamp 1682952543
transform 1 0 2412 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5122
timestamp 1682952543
transform 1 0 2468 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1682952543
transform 1 0 2484 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5124
timestamp 1682952543
transform 1 0 2500 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1682952543
transform 1 0 2388 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5129
timestamp 1682952543
transform 1 0 2412 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5190
timestamp 1682952543
transform 1 0 2372 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1682952543
transform 1 0 2388 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1682952543
transform 1 0 2452 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5235
timestamp 1682952543
transform 1 0 2492 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5236
timestamp 1682952543
transform 1 0 2508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1682952543
transform 1 0 2516 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5193
timestamp 1682952543
transform 1 0 2508 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5125
timestamp 1682952543
transform 1 0 2532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1682952543
transform 1 0 2540 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5008
timestamp 1682952543
transform 1 0 2572 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5021
timestamp 1682952543
transform 1 0 2580 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5051
timestamp 1682952543
transform 1 0 2564 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5237
timestamp 1682952543
transform 1 0 2548 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5194
timestamp 1682952543
transform 1 0 2548 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5022
timestamp 1682952543
transform 1 0 2612 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5080
timestamp 1682952543
transform 1 0 2580 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5081
timestamp 1682952543
transform 1 0 2604 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5127
timestamp 1682952543
transform 1 0 2580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1682952543
transform 1 0 2596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1682952543
transform 1 0 2604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5238
timestamp 1682952543
transform 1 0 2564 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1682952543
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1682952543
transform 1 0 2588 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1682952543
transform 1 0 2564 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5023
timestamp 1682952543
transform 1 0 2628 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5009
timestamp 1682952543
transform 1 0 2668 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5082
timestamp 1682952543
transform 1 0 2644 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1682952543
transform 1 0 2700 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1682952543
transform 1 0 2724 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5130
timestamp 1682952543
transform 1 0 2636 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5131
timestamp 1682952543
transform 1 0 2644 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1682952543
transform 1 0 2692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5241
timestamp 1682952543
transform 1 0 2628 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5281
timestamp 1682952543
transform 1 0 2620 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5026
timestamp 1682952543
transform 1 0 2764 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5133
timestamp 1682952543
transform 1 0 2748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1682952543
transform 1 0 2724 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1682952543
transform 1 0 2740 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5150
timestamp 1682952543
transform 1 0 2724 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5130
timestamp 1682952543
transform 1 0 2748 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5085
timestamp 1682952543
transform 1 0 2908 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5134
timestamp 1682952543
transform 1 0 2820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5135
timestamp 1682952543
transform 1 0 2828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5136
timestamp 1682952543
transform 1 0 2884 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5131
timestamp 1682952543
transform 1 0 2820 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5244
timestamp 1682952543
transform 1 0 2908 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5151
timestamp 1682952543
transform 1 0 2884 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5245
timestamp 1682952543
transform 1 0 2932 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5132
timestamp 1682952543
transform 1 0 2940 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5086
timestamp 1682952543
transform 1 0 2956 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5137
timestamp 1682952543
transform 1 0 2956 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1682952543
transform 1 0 2980 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5246
timestamp 1682952543
transform 1 0 2964 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1682952543
transform 1 0 2980 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5152
timestamp 1682952543
transform 1 0 2964 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5058
timestamp 1682952543
transform 1 0 2996 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1682952543
transform 1 0 2996 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5010
timestamp 1682952543
transform 1 0 3036 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5048
timestamp 1682952543
transform 1 0 3036 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5248
timestamp 1682952543
transform 1 0 3044 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5049
timestamp 1682952543
transform 1 0 3092 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5140
timestamp 1682952543
transform 1 0 3100 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5133
timestamp 1682952543
transform 1 0 3084 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5050
timestamp 1682952543
transform 1 0 3116 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_5107
timestamp 1682952543
transform 1 0 3116 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1682952543
transform 1 0 3108 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5195
timestamp 1682952543
transform 1 0 3092 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5011
timestamp 1682952543
transform 1 0 3132 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1682952543
transform 1 0 3156 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5059
timestamp 1682952543
transform 1 0 3132 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1682952543
transform 1 0 3140 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5087
timestamp 1682952543
transform 1 0 3148 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5141
timestamp 1682952543
transform 1 0 3148 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5134
timestamp 1682952543
transform 1 0 3140 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5154
timestamp 1682952543
transform 1 0 3140 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5061
timestamp 1682952543
transform 1 0 3180 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5142
timestamp 1682952543
transform 1 0 3188 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5088
timestamp 1682952543
transform 1 0 3228 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5143
timestamp 1682952543
transform 1 0 3212 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5108
timestamp 1682952543
transform 1 0 3220 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5144
timestamp 1682952543
transform 1 0 3228 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1682952543
transform 1 0 3212 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5250
timestamp 1682952543
transform 1 0 3220 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5028
timestamp 1682952543
transform 1 0 3268 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5089
timestamp 1682952543
transform 1 0 3260 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5145
timestamp 1682952543
transform 1 0 3252 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5155
timestamp 1682952543
transform 1 0 3244 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1682952543
transform 1 0 3212 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5012
timestamp 1682952543
transform 1 0 3300 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5090
timestamp 1682952543
transform 1 0 3292 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5146
timestamp 1682952543
transform 1 0 3268 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1682952543
transform 1 0 3276 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5148
timestamp 1682952543
transform 1 0 3292 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1682952543
transform 1 0 3260 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1682952543
transform 1 0 3268 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5253
timestamp 1682952543
transform 1 0 3284 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5135
timestamp 1682952543
transform 1 0 3292 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5109
timestamp 1682952543
transform 1 0 3308 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5254
timestamp 1682952543
transform 1 0 3300 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5156
timestamp 1682952543
transform 1 0 3268 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1682952543
transform 1 0 3300 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5197
timestamp 1682952543
transform 1 0 3284 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5029
timestamp 1682952543
transform 1 0 3372 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5149
timestamp 1682952543
transform 1 0 3356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1682952543
transform 1 0 3332 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5136
timestamp 1682952543
transform 1 0 3356 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1682952543
transform 1 0 3380 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5198
timestamp 1682952543
transform 1 0 3332 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1682952543
transform 1 0 3348 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5013
timestamp 1682952543
transform 1 0 3444 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5030
timestamp 1682952543
transform 1 0 3436 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5091
timestamp 1682952543
transform 1 0 3428 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5062
timestamp 1682952543
transform 1 0 3436 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1682952543
transform 1 0 3428 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5031
timestamp 1682952543
transform 1 0 3460 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5051
timestamp 1682952543
transform 1 0 3460 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_5092
timestamp 1682952543
transform 1 0 3468 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5063
timestamp 1682952543
transform 1 0 3476 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5151
timestamp 1682952543
transform 1 0 3468 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5137
timestamp 1682952543
transform 1 0 3468 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5200
timestamp 1682952543
transform 1 0 3452 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5014
timestamp 1682952543
transform 1 0 3532 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5093
timestamp 1682952543
transform 1 0 3516 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1682952543
transform 1 0 3508 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5152
timestamp 1682952543
transform 1 0 3516 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1682952543
transform 1 0 3532 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5154
timestamp 1682952543
transform 1 0 3540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1682952543
transform 1 0 3548 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5111
timestamp 1682952543
transform 1 0 3556 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5156
timestamp 1682952543
transform 1 0 3564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1682952543
transform 1 0 3612 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1682952543
transform 1 0 3500 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5257
timestamp 1682952543
transform 1 0 3508 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5258
timestamp 1682952543
transform 1 0 3524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1682952543
transform 1 0 3540 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5260
timestamp 1682952543
transform 1 0 3556 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1682952543
transform 1 0 3572 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5262
timestamp 1682952543
transform 1 0 3588 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5201
timestamp 1682952543
transform 1 0 3500 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1682952543
transform 1 0 3556 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1682952543
transform 1 0 3612 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5032
timestamp 1682952543
transform 1 0 3708 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5094
timestamp 1682952543
transform 1 0 3700 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5158
timestamp 1682952543
transform 1 0 3700 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5159
timestamp 1682952543
transform 1 0 3724 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5015
timestamp 1682952543
transform 1 0 3748 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5016
timestamp 1682952543
transform 1 0 3764 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5263
timestamp 1682952543
transform 1 0 3740 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5161
timestamp 1682952543
transform 1 0 3740 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5024
timestamp 1682952543
transform 1 0 3764 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5052
timestamp 1682952543
transform 1 0 3764 0 1 2035
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1682952543
transform 1 0 3756 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5095
timestamp 1682952543
transform 1 0 3772 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5160
timestamp 1682952543
transform 1 0 3772 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5033
timestamp 1682952543
transform 1 0 3804 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5065
timestamp 1682952543
transform 1 0 3796 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5161
timestamp 1682952543
transform 1 0 3788 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5162
timestamp 1682952543
transform 1 0 3788 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5112
timestamp 1682952543
transform 1 0 3804 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5052
timestamp 1682952543
transform 1 0 3836 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5096
timestamp 1682952543
transform 1 0 3828 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5162
timestamp 1682952543
transform 1 0 3812 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5163
timestamp 1682952543
transform 1 0 3828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5164
timestamp 1682952543
transform 1 0 3844 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1682952543
transform 1 0 3852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5166
timestamp 1682952543
transform 1 0 3876 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1682952543
transform 1 0 3804 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5053
timestamp 1682952543
transform 1 0 3964 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5054
timestamp 1682952543
transform 1 0 4004 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5097
timestamp 1682952543
transform 1 0 3980 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5098
timestamp 1682952543
transform 1 0 4004 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5167
timestamp 1682952543
transform 1 0 3924 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1682952543
transform 1 0 3844 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1682952543
transform 1 0 3852 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1682952543
transform 1 0 3868 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5268
timestamp 1682952543
transform 1 0 3884 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1682952543
transform 1 0 3900 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5163
timestamp 1682952543
transform 1 0 3820 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5164
timestamp 1682952543
transform 1 0 3836 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1682952543
transform 1 0 3852 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1682952543
transform 1 0 3868 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1682952543
transform 1 0 3844 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5203
timestamp 1682952543
transform 1 0 3876 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5167
timestamp 1682952543
transform 1 0 3924 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5055
timestamp 1682952543
transform 1 0 4036 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5168
timestamp 1682952543
transform 1 0 3996 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1682952543
transform 1 0 4004 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5170
timestamp 1682952543
transform 1 0 4028 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5113
timestamp 1682952543
transform 1 0 4036 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5056
timestamp 1682952543
transform 1 0 4140 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5171
timestamp 1682952543
transform 1 0 4076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5172
timestamp 1682952543
transform 1 0 4132 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1682952543
transform 1 0 4140 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5270
timestamp 1682952543
transform 1 0 4004 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1682952543
transform 1 0 4020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1682952543
transform 1 0 4036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1682952543
transform 1 0 4052 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5168
timestamp 1682952543
transform 1 0 4020 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1682952543
transform 1 0 4076 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5204
timestamp 1682952543
transform 1 0 3996 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5205
timestamp 1682952543
transform 1 0 4012 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5206
timestamp 1682952543
transform 1 0 4036 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5274
timestamp 1682952543
transform 1 0 4148 0 1 2005
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_42
timestamp 1682952543
transform 1 0 48 0 1 1970
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_321
timestamp 1682952543
transform 1 0 72 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_361
timestamp 1682952543
transform -1 0 184 0 1 1970
box -9 -3 26 105
use FILL  FILL_1805
timestamp 1682952543
transform 1 0 184 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_206
timestamp 1682952543
transform 1 0 192 0 1 1970
box -8 -3 46 105
use FILL  FILL_1806
timestamp 1682952543
transform 1 0 232 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_323
timestamp 1682952543
transform -1 0 336 0 1 1970
box -8 -3 104 105
use FILL  FILL_1807
timestamp 1682952543
transform 1 0 336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1682952543
transform 1 0 344 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5207
timestamp 1682952543
transform 1 0 388 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_220
timestamp 1682952543
transform -1 0 392 0 1 1970
box -8 -3 46 105
use FILL  FILL_1809
timestamp 1682952543
transform 1 0 392 0 1 1970
box -8 -3 16 105
use FILL  FILL_1810
timestamp 1682952543
transform 1 0 400 0 1 1970
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1682952543
transform 1 0 408 0 1 1970
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1682952543
transform 1 0 416 0 1 1970
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1682952543
transform 1 0 424 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_207
timestamp 1682952543
transform 1 0 432 0 1 1970
box -8 -3 46 105
use FILL  FILL_1814
timestamp 1682952543
transform 1 0 472 0 1 1970
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1682952543
transform 1 0 480 0 1 1970
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1682952543
transform 1 0 488 0 1 1970
box -8 -3 16 105
use FILL  FILL_1817
timestamp 1682952543
transform 1 0 496 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_362
timestamp 1682952543
transform 1 0 504 0 1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_324
timestamp 1682952543
transform -1 0 616 0 1 1970
box -8 -3 104 105
use FILL  FILL_1818
timestamp 1682952543
transform 1 0 616 0 1 1970
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1682952543
transform 1 0 624 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_62
timestamp 1682952543
transform 1 0 632 0 1 1970
box -8 -3 32 105
use FILL  FILL_1825
timestamp 1682952543
transform 1 0 656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1682952543
transform 1 0 664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1830
timestamp 1682952543
transform 1 0 672 0 1 1970
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1682952543
transform 1 0 680 0 1 1970
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1682952543
transform 1 0 688 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_68
timestamp 1682952543
transform 1 0 696 0 1 1970
box -8 -3 34 105
use FILL  FILL_1833
timestamp 1682952543
transform 1 0 728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1837
timestamp 1682952543
transform 1 0 736 0 1 1970
box -8 -3 16 105
use FILL  FILL_1839
timestamp 1682952543
transform 1 0 744 0 1 1970
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1682952543
transform 1 0 752 0 1 1970
box -8 -3 16 105
use FILL  FILL_1842
timestamp 1682952543
transform 1 0 760 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_210
timestamp 1682952543
transform 1 0 768 0 1 1970
box -8 -3 46 105
use FILL  FILL_1843
timestamp 1682952543
transform 1 0 808 0 1 1970
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1682952543
transform 1 0 816 0 1 1970
box -8 -3 16 105
use FILL  FILL_1848
timestamp 1682952543
transform 1 0 824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1682952543
transform 1 0 832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1682952543
transform 1 0 840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1854
timestamp 1682952543
transform 1 0 848 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_211
timestamp 1682952543
transform 1 0 856 0 1 1970
box -8 -3 46 105
use FILL  FILL_1855
timestamp 1682952543
transform 1 0 896 0 1 1970
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1682952543
transform 1 0 904 0 1 1970
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1682952543
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1682952543
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1682952543
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1682952543
transform 1 0 936 0 1 1970
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1682952543
transform 1 0 944 0 1 1970
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1682952543
transform 1 0 952 0 1 1970
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1682952543
transform 1 0 960 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_213
timestamp 1682952543
transform 1 0 968 0 1 1970
box -8 -3 46 105
use FILL  FILL_1868
timestamp 1682952543
transform 1 0 1008 0 1 1970
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1682952543
transform 1 0 1016 0 1 1970
box -8 -3 16 105
use FILL  FILL_1875
timestamp 1682952543
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1682952543
transform 1 0 1032 0 1 1970
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1682952543
transform 1 0 1040 0 1 1970
box -8 -3 16 105
use FILL  FILL_1881
timestamp 1682952543
transform 1 0 1048 0 1 1970
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1682952543
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1682952543
transform 1 0 1064 0 1 1970
box -8 -3 16 105
use FILL  FILL_1884
timestamp 1682952543
transform 1 0 1072 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_69
timestamp 1682952543
transform -1 0 1112 0 1 1970
box -8 -3 34 105
use FILL  FILL_1885
timestamp 1682952543
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1682952543
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_1891
timestamp 1682952543
transform 1 0 1128 0 1 1970
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1682952543
transform 1 0 1136 0 1 1970
box -8 -3 16 105
use FILL  FILL_1895
timestamp 1682952543
transform 1 0 1144 0 1 1970
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1682952543
transform 1 0 1152 0 1 1970
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1682952543
transform 1 0 1160 0 1 1970
box -8 -3 16 105
use FILL  FILL_1898
timestamp 1682952543
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1682952543
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_71
timestamp 1682952543
transform -1 0 1216 0 1 1970
box -8 -3 34 105
use FILL  FILL_1900
timestamp 1682952543
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_1901
timestamp 1682952543
transform 1 0 1224 0 1 1970
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1682952543
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use FILL  FILL_1903
timestamp 1682952543
transform 1 0 1240 0 1 1970
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1682952543
transform 1 0 1248 0 1 1970
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1682952543
transform 1 0 1256 0 1 1970
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1682952543
transform 1 0 1264 0 1 1970
box -8 -3 16 105
use FILL  FILL_1909
timestamp 1682952543
transform 1 0 1272 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_223
timestamp 1682952543
transform -1 0 1320 0 1 1970
box -8 -3 46 105
use FILL  FILL_1910
timestamp 1682952543
transform 1 0 1320 0 1 1970
box -8 -3 16 105
use FILL  FILL_1911
timestamp 1682952543
transform 1 0 1328 0 1 1970
box -8 -3 16 105
use FILL  FILL_1915
timestamp 1682952543
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1682952543
transform 1 0 1344 0 1 1970
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1682952543
transform 1 0 1352 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_367
timestamp 1682952543
transform -1 0 1376 0 1 1970
box -9 -3 26 105
use M3_M2  M3_M2_5208
timestamp 1682952543
transform 1 0 1476 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_329
timestamp 1682952543
transform -1 0 1472 0 1 1970
box -8 -3 104 105
use BUFX2  BUFX2_68
timestamp 1682952543
transform -1 0 1496 0 1 1970
box -5 -3 28 105
use M3_M2  M3_M2_5209
timestamp 1682952543
transform 1 0 1516 0 1 1975
box -3 -3 3 3
use BUFX2  BUFX2_69
timestamp 1682952543
transform 1 0 1496 0 1 1970
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_330
timestamp 1682952543
transform 1 0 1520 0 1 1970
box -8 -3 104 105
use OAI22X1  OAI22X1_225
timestamp 1682952543
transform -1 0 1656 0 1 1970
box -8 -3 46 105
use FILL  FILL_1919
timestamp 1682952543
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1682952543
transform 1 0 1664 0 1 1970
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1682952543
transform 1 0 1672 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_227
timestamp 1682952543
transform -1 0 1720 0 1 1970
box -8 -3 46 105
use FILL  FILL_1931
timestamp 1682952543
transform 1 0 1720 0 1 1970
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1682952543
transform 1 0 1728 0 1 1970
box -8 -3 16 105
use FILL  FILL_1937
timestamp 1682952543
transform 1 0 1736 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_74
timestamp 1682952543
transform 1 0 1744 0 1 1970
box -5 -3 28 105
use FILL  FILL_1939
timestamp 1682952543
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1682952543
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5210
timestamp 1682952543
transform 1 0 1812 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_229
timestamp 1682952543
transform -1 0 1824 0 1 1970
box -8 -3 46 105
use FILL  FILL_1941
timestamp 1682952543
transform 1 0 1824 0 1 1970
box -8 -3 16 105
use FILL  FILL_1942
timestamp 1682952543
transform 1 0 1832 0 1 1970
box -8 -3 16 105
use FILL  FILL_1943
timestamp 1682952543
transform 1 0 1840 0 1 1970
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1682952543
transform 1 0 1848 0 1 1970
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1682952543
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5211
timestamp 1682952543
transform 1 0 1876 0 1 1975
box -3 -3 3 3
use FILL  FILL_1946
timestamp 1682952543
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_230
timestamp 1682952543
transform 1 0 1872 0 1 1970
box -8 -3 46 105
use FILL  FILL_1949
timestamp 1682952543
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1682952543
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use FILL  FILL_1955
timestamp 1682952543
transform 1 0 1928 0 1 1970
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1682952543
transform 1 0 1936 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5212
timestamp 1682952543
transform 1 0 1956 0 1 1975
box -3 -3 3 3
use FILL  FILL_1958
timestamp 1682952543
transform 1 0 1944 0 1 1970
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1682952543
transform 1 0 1952 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_35
timestamp 1682952543
transform -1 0 1992 0 1 1970
box -8 -3 40 105
use M3_M2  M3_M2_5213
timestamp 1682952543
transform 1 0 2004 0 1 1975
box -3 -3 3 3
use FILL  FILL_1960
timestamp 1682952543
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1682952543
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_1966
timestamp 1682952543
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_370
timestamp 1682952543
transform -1 0 2032 0 1 1970
box -9 -3 26 105
use FILL  FILL_1967
timestamp 1682952543
transform 1 0 2032 0 1 1970
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1682952543
transform 1 0 2040 0 1 1970
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1682952543
transform 1 0 2048 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_76
timestamp 1682952543
transform -1 0 2080 0 1 1970
box -5 -3 28 105
use FILL  FILL_1970
timestamp 1682952543
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_1971
timestamp 1682952543
transform 1 0 2088 0 1 1970
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1682952543
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5214
timestamp 1682952543
transform 1 0 2116 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_231
timestamp 1682952543
transform 1 0 2104 0 1 1970
box -8 -3 46 105
use FILL  FILL_1973
timestamp 1682952543
transform 1 0 2144 0 1 1970
box -8 -3 16 105
use FILL  FILL_1974
timestamp 1682952543
transform 1 0 2152 0 1 1970
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1682952543
transform 1 0 2160 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_232
timestamp 1682952543
transform -1 0 2208 0 1 1970
box -8 -3 46 105
use FILL  FILL_1976
timestamp 1682952543
transform 1 0 2208 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_233
timestamp 1682952543
transform -1 0 2256 0 1 1970
box -8 -3 46 105
use NOR2X1  NOR2X1_66
timestamp 1682952543
transform 1 0 2256 0 1 1970
box -8 -3 32 105
use M3_M2  M3_M2_5215
timestamp 1682952543
transform 1 0 2356 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_333
timestamp 1682952543
transform -1 0 2376 0 1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5216
timestamp 1682952543
transform 1 0 2412 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_334
timestamp 1682952543
transform 1 0 2376 0 1 1970
box -8 -3 104 105
use OAI22X1  OAI22X1_234
timestamp 1682952543
transform 1 0 2472 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_5217
timestamp 1682952543
transform 1 0 2524 0 1 1975
box -3 -3 3 3
use NOR2X1  NOR2X1_67
timestamp 1682952543
transform 1 0 2512 0 1 1970
box -8 -3 32 105
use FILL  FILL_1977
timestamp 1682952543
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5218
timestamp 1682952543
transform 1 0 2572 0 1 1975
box -3 -3 3 3
use NOR2X1  NOR2X1_68
timestamp 1682952543
transform -1 0 2568 0 1 1970
box -8 -3 32 105
use M3_M2  M3_M2_5219
timestamp 1682952543
transform 1 0 2604 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_235
timestamp 1682952543
transform -1 0 2608 0 1 1970
box -8 -3 46 105
use FILL  FILL_1978
timestamp 1682952543
transform 1 0 2608 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_70
timestamp 1682952543
transform 1 0 2616 0 1 1970
box -8 -3 32 105
use M3_M2  M3_M2_5220
timestamp 1682952543
transform 1 0 2660 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5221
timestamp 1682952543
transform 1 0 2724 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_338
timestamp 1682952543
transform -1 0 2736 0 1 1970
box -8 -3 104 105
use AND2X2  AND2X2_47
timestamp 1682952543
transform 1 0 2736 0 1 1970
box -8 -3 40 105
use FILL  FILL_1995
timestamp 1682952543
transform 1 0 2768 0 1 1970
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1682952543
transform 1 0 2776 0 1 1970
box -8 -3 16 105
use FILL  FILL_1997
timestamp 1682952543
transform 1 0 2784 0 1 1970
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1682952543
transform 1 0 2792 0 1 1970
box -8 -3 16 105
use FILL  FILL_1999
timestamp 1682952543
transform 1 0 2800 0 1 1970
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1682952543
transform 1 0 2808 0 1 1970
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1682952543
transform 1 0 2816 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5222
timestamp 1682952543
transform 1 0 2908 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_339
timestamp 1682952543
transform -1 0 2920 0 1 1970
box -8 -3 104 105
use FILL  FILL_2002
timestamp 1682952543
transform 1 0 2920 0 1 1970
box -8 -3 16 105
use FILL  FILL_2012
timestamp 1682952543
transform 1 0 2928 0 1 1970
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1682952543
transform 1 0 2936 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_236
timestamp 1682952543
transform -1 0 2984 0 1 1970
box -8 -3 46 105
use FILL  FILL_2014
timestamp 1682952543
transform 1 0 2984 0 1 1970
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1682952543
transform 1 0 2992 0 1 1970
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1682952543
transform 1 0 3000 0 1 1970
box -8 -3 16 105
use FILL  FILL_2020
timestamp 1682952543
transform 1 0 3008 0 1 1970
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1682952543
transform 1 0 3016 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5223
timestamp 1682952543
transform 1 0 3036 0 1 1975
box -3 -3 3 3
use M3_M2  M3_M2_5224
timestamp 1682952543
transform 1 0 3052 0 1 1975
box -3 -3 3 3
use NAND3X1  NAND3X1_40
timestamp 1682952543
transform -1 0 3056 0 1 1970
box -8 -3 40 105
use FILL  FILL_2022
timestamp 1682952543
transform 1 0 3056 0 1 1970
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1682952543
transform 1 0 3064 0 1 1970
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1682952543
transform 1 0 3072 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_41
timestamp 1682952543
transform -1 0 3112 0 1 1970
box -8 -3 40 105
use FILL  FILL_2025
timestamp 1682952543
transform 1 0 3112 0 1 1970
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1682952543
transform 1 0 3120 0 1 1970
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1682952543
transform 1 0 3128 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_42
timestamp 1682952543
transform 1 0 3136 0 1 1970
box -8 -3 40 105
use FILL  FILL_2032
timestamp 1682952543
transform 1 0 3168 0 1 1970
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1682952543
transform 1 0 3176 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_77
timestamp 1682952543
transform 1 0 3184 0 1 1970
box -5 -3 28 105
use AOI22X1  AOI22X1_216
timestamp 1682952543
transform -1 0 3248 0 1 1970
box -8 -3 46 105
use FILL  FILL_2036
timestamp 1682952543
transform 1 0 3248 0 1 1970
box -8 -3 16 105
use FILL  FILL_2037
timestamp 1682952543
transform 1 0 3256 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_238
timestamp 1682952543
transform 1 0 3264 0 1 1970
box -8 -3 46 105
use FILL  FILL_2038
timestamp 1682952543
transform 1 0 3304 0 1 1970
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1682952543
transform 1 0 3312 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_343
timestamp 1682952543
transform 1 0 3320 0 1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5225
timestamp 1682952543
transform 1 0 3436 0 1 1975
box -3 -3 3 3
use INVX2  INVX2_374
timestamp 1682952543
transform 1 0 3416 0 1 1970
box -9 -3 26 105
use FILL  FILL_2044
timestamp 1682952543
transform 1 0 3432 0 1 1970
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1682952543
transform 1 0 3440 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5226
timestamp 1682952543
transform 1 0 3468 0 1 1975
box -3 -3 3 3
use NAND3X1  NAND3X1_44
timestamp 1682952543
transform -1 0 3480 0 1 1970
box -8 -3 40 105
use FILL  FILL_2046
timestamp 1682952543
transform 1 0 3480 0 1 1970
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1682952543
transform 1 0 3488 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5227
timestamp 1682952543
transform 1 0 3508 0 1 1975
box -3 -3 3 3
use AOI22X1  AOI22X1_217
timestamp 1682952543
transform 1 0 3496 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_239
timestamp 1682952543
transform 1 0 3536 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_5228
timestamp 1682952543
transform 1 0 3676 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_344
timestamp 1682952543
transform 1 0 3576 0 1 1970
box -8 -3 104 105
use FILL  FILL_2048
timestamp 1682952543
transform 1 0 3672 0 1 1970
box -8 -3 16 105
use FILL  FILL_2049
timestamp 1682952543
transform 1 0 3680 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_375
timestamp 1682952543
transform 1 0 3688 0 1 1970
box -9 -3 26 105
use FILL  FILL_2050
timestamp 1682952543
transform 1 0 3704 0 1 1970
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1682952543
transform 1 0 3712 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_78
timestamp 1682952543
transform 1 0 3720 0 1 1970
box -5 -3 28 105
use FILL  FILL_2052
timestamp 1682952543
transform 1 0 3744 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_45
timestamp 1682952543
transform -1 0 3784 0 1 1970
box -8 -3 40 105
use FILL  FILL_2053
timestamp 1682952543
transform 1 0 3784 0 1 1970
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1682952543
transform 1 0 3792 0 1 1970
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1682952543
transform 1 0 3800 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_218
timestamp 1682952543
transform 1 0 3808 0 1 1970
box -8 -3 46 105
use OAI22X1  OAI22X1_240
timestamp 1682952543
transform 1 0 3848 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_5229
timestamp 1682952543
transform 1 0 3956 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_345
timestamp 1682952543
transform 1 0 3888 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_376
timestamp 1682952543
transform 1 0 3984 0 1 1970
box -9 -3 26 105
use OAI22X1  OAI22X1_241
timestamp 1682952543
transform 1 0 4000 0 1 1970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_346
timestamp 1682952543
transform 1 0 4040 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_377
timestamp 1682952543
transform -1 0 4152 0 1 1970
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_43
timestamp 1682952543
transform 1 0 4177 0 1 1970
box -10 -3 10 3
use M3_M2  M3_M2_5263
timestamp 1682952543
transform 1 0 84 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1682952543
transform 1 0 148 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5287
timestamp 1682952543
transform 1 0 84 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5372
timestamp 1682952543
transform 1 0 124 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5354
timestamp 1682952543
transform 1 0 148 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5230
timestamp 1682952543
transform 1 0 196 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5282
timestamp 1682952543
transform 1 0 188 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5283
timestamp 1682952543
transform 1 0 212 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5288
timestamp 1682952543
transform 1 0 188 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5289
timestamp 1682952543
transform 1 0 196 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5290
timestamp 1682952543
transform 1 0 212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5373
timestamp 1682952543
transform 1 0 164 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5374
timestamp 1682952543
transform 1 0 172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1682952543
transform 1 0 188 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5355
timestamp 1682952543
transform 1 0 196 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5231
timestamp 1682952543
transform 1 0 260 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5264
timestamp 1682952543
transform 1 0 236 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5265
timestamp 1682952543
transform 1 0 276 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5266
timestamp 1682952543
transform 1 0 428 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5291
timestamp 1682952543
transform 1 0 236 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5333
timestamp 1682952543
transform 1 0 316 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5292
timestamp 1682952543
transform 1 0 332 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5334
timestamp 1682952543
transform 1 0 412 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5284
timestamp 1682952543
transform 1 0 460 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5293
timestamp 1682952543
transform 1 0 420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5294
timestamp 1682952543
transform 1 0 436 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1682952543
transform 1 0 452 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1682952543
transform 1 0 460 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1682952543
transform 1 0 204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5377
timestamp 1682952543
transform 1 0 220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5378
timestamp 1682952543
transform 1 0 268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1682952543
transform 1 0 316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5380
timestamp 1682952543
transform 1 0 364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5381
timestamp 1682952543
transform 1 0 412 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5379
timestamp 1682952543
transform 1 0 124 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1682952543
transform 1 0 172 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5381
timestamp 1682952543
transform 1 0 188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5416
timestamp 1682952543
transform 1 0 164 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5417
timestamp 1682952543
transform 1 0 212 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1682952543
transform 1 0 276 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5356
timestamp 1682952543
transform 1 0 420 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5382
timestamp 1682952543
transform 1 0 428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5383
timestamp 1682952543
transform 1 0 460 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5383
timestamp 1682952543
transform 1 0 412 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5384
timestamp 1682952543
transform 1 0 428 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1682952543
transform 1 0 452 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1682952543
transform 1 0 460 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5232
timestamp 1682952543
transform 1 0 500 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5267
timestamp 1682952543
transform 1 0 508 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5297
timestamp 1682952543
transform 1 0 500 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5335
timestamp 1682952543
transform 1 0 516 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5298
timestamp 1682952543
transform 1 0 524 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5384
timestamp 1682952543
transform 1 0 492 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5357
timestamp 1682952543
transform 1 0 500 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5385
timestamp 1682952543
transform 1 0 508 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5418
timestamp 1682952543
transform 1 0 492 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5440
timestamp 1682952543
transform 1 0 484 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1682952543
transform 1 0 508 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1682952543
transform 1 0 580 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1682952543
transform 1 0 612 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5299
timestamp 1682952543
transform 1 0 540 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5336
timestamp 1682952543
transform 1 0 620 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5358
timestamp 1682952543
transform 1 0 580 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5386
timestamp 1682952543
transform 1 0 588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5387
timestamp 1682952543
transform 1 0 620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5388
timestamp 1682952543
transform 1 0 628 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5386
timestamp 1682952543
transform 1 0 588 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5387
timestamp 1682952543
transform 1 0 628 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1682952543
transform 1 0 660 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5389
timestamp 1682952543
transform 1 0 660 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5388
timestamp 1682952543
transform 1 0 660 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1682952543
transform 1 0 700 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5300
timestamp 1682952543
transform 1 0 676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1682952543
transform 1 0 684 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1682952543
transform 1 0 700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1682952543
transform 1 0 692 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5389
timestamp 1682952543
transform 1 0 708 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5233
timestamp 1682952543
transform 1 0 724 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5282
timestamp 1682952543
transform 1 0 724 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5338
timestamp 1682952543
transform 1 0 724 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5391
timestamp 1682952543
transform 1 0 724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1682952543
transform 1 0 772 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5390
timestamp 1682952543
transform 1 0 772 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5303
timestamp 1682952543
transform 1 0 796 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5392
timestamp 1682952543
transform 1 0 788 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5234
timestamp 1682952543
transform 1 0 836 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5284
timestamp 1682952543
transform 1 0 828 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5288
timestamp 1682952543
transform 1 0 836 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5304
timestamp 1682952543
transform 1 0 836 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5441
timestamp 1682952543
transform 1 0 828 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1682952543
transform 1 0 876 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5305
timestamp 1682952543
transform 1 0 860 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1682952543
transform 1 0 868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1682952543
transform 1 0 852 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5339
timestamp 1682952543
transform 1 0 892 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5394
timestamp 1682952543
transform 1 0 868 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1682952543
transform 1 0 876 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5396
timestamp 1682952543
transform 1 0 892 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5397
timestamp 1682952543
transform 1 0 908 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5391
timestamp 1682952543
transform 1 0 892 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1682952543
transform 1 0 876 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5443
timestamp 1682952543
transform 1 0 900 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5392
timestamp 1682952543
transform 1 0 916 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5290
timestamp 1682952543
transform 1 0 972 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5307
timestamp 1682952543
transform 1 0 956 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1682952543
transform 1 0 964 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5398
timestamp 1682952543
transform 1 0 956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5399
timestamp 1682952543
transform 1 0 972 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5455
timestamp 1682952543
transform 1 0 972 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1682952543
transform 1 0 996 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1682952543
transform 1 0 1012 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5400
timestamp 1682952543
transform 1 0 1004 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1682952543
transform 1 0 1028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5310
timestamp 1682952543
transform 1 0 1036 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5292
timestamp 1682952543
transform 1 0 1060 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5311
timestamp 1682952543
transform 1 0 1068 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5293
timestamp 1682952543
transform 1 0 1092 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5312
timestamp 1682952543
transform 1 0 1092 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1682952543
transform 1 0 1060 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5359
timestamp 1682952543
transform 1 0 1068 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5360
timestamp 1682952543
transform 1 0 1084 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5480
timestamp 1682952543
transform 1 0 1068 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5393
timestamp 1682952543
transform 1 0 1084 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5402
timestamp 1682952543
transform 1 0 1100 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5236
timestamp 1682952543
transform 1 0 1116 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5294
timestamp 1682952543
transform 1 0 1116 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5394
timestamp 1682952543
transform 1 0 1116 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1682952543
transform 1 0 1172 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5296
timestamp 1682952543
transform 1 0 1188 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5313
timestamp 1682952543
transform 1 0 1156 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5361
timestamp 1682952543
transform 1 0 1156 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5403
timestamp 1682952543
transform 1 0 1188 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5395
timestamp 1682952543
transform 1 0 1188 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5396
timestamp 1682952543
transform 1 0 1228 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5444
timestamp 1682952543
transform 1 0 1156 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5445
timestamp 1682952543
transform 1 0 1196 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5237
timestamp 1682952543
transform 1 0 1260 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5404
timestamp 1682952543
transform 1 0 1260 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5362
timestamp 1682952543
transform 1 0 1276 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1682952543
transform 1 0 1268 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5314
timestamp 1682952543
transform 1 0 1284 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5405
timestamp 1682952543
transform 1 0 1284 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5238
timestamp 1682952543
transform 1 0 1316 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5297
timestamp 1682952543
transform 1 0 1308 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5315
timestamp 1682952543
transform 1 0 1308 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1682952543
transform 1 0 1332 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5406
timestamp 1682952543
transform 1 0 1300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5407
timestamp 1682952543
transform 1 0 1316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1682952543
transform 1 0 1324 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1682952543
transform 1 0 1348 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5239
timestamp 1682952543
transform 1 0 1372 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1682952543
transform 1 0 1388 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1682952543
transform 1 0 1372 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5318
timestamp 1682952543
transform 1 0 1372 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5319
timestamp 1682952543
transform 1 0 1388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5409
timestamp 1682952543
transform 1 0 1364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5410
timestamp 1682952543
transform 1 0 1380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1682952543
transform 1 0 1388 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5241
timestamp 1682952543
transform 1 0 1460 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1682952543
transform 1 0 1444 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5320
timestamp 1682952543
transform 1 0 1492 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1682952543
transform 1 0 1444 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5363
timestamp 1682952543
transform 1 0 1452 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5364
timestamp 1682952543
transform 1 0 1492 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5268
timestamp 1682952543
transform 1 0 1516 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5413
timestamp 1682952543
transform 1 0 1508 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5446
timestamp 1682952543
transform 1 0 1460 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5242
timestamp 1682952543
transform 1 0 1532 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1682952543
transform 1 0 1540 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5321
timestamp 1682952543
transform 1 0 1532 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5269
timestamp 1682952543
transform 1 0 1572 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1682952543
transform 1 0 1564 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5322
timestamp 1682952543
transform 1 0 1564 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5302
timestamp 1682952543
transform 1 0 1604 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5414
timestamp 1682952543
transform 1 0 1604 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5243
timestamp 1682952543
transform 1 0 1644 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5323
timestamp 1682952543
transform 1 0 1628 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5324
timestamp 1682952543
transform 1 0 1636 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5365
timestamp 1682952543
transform 1 0 1636 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5419
timestamp 1682952543
transform 1 0 1636 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1682952543
transform 1 0 1652 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5415
timestamp 1682952543
transform 1 0 1652 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5325
timestamp 1682952543
transform 1 0 1668 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5420
timestamp 1682952543
transform 1 0 1660 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1682952543
transform 1 0 1676 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5326
timestamp 1682952543
transform 1 0 1692 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5341
timestamp 1682952543
transform 1 0 1700 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1682952543
transform 1 0 1724 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5342
timestamp 1682952543
transform 1 0 1716 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5416
timestamp 1682952543
transform 1 0 1684 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5417
timestamp 1682952543
transform 1 0 1708 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5421
timestamp 1682952543
transform 1 0 1684 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5366
timestamp 1682952543
transform 1 0 1732 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5327
timestamp 1682952543
transform 1 0 1748 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5328
timestamp 1682952543
transform 1 0 1756 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5305
timestamp 1682952543
transform 1 0 1796 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5329
timestamp 1682952543
transform 1 0 1780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5418
timestamp 1682952543
transform 1 0 1764 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5419
timestamp 1682952543
transform 1 0 1804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5420
timestamp 1682952543
transform 1 0 1860 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5422
timestamp 1682952543
transform 1 0 1764 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5423
timestamp 1682952543
transform 1 0 1804 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5421
timestamp 1682952543
transform 1 0 1876 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5306
timestamp 1682952543
transform 1 0 1908 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5330
timestamp 1682952543
transform 1 0 1908 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1682952543
transform 1 0 1940 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1682952543
transform 1 0 1964 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5307
timestamp 1682952543
transform 1 0 1980 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5496
timestamp 1682952543
transform 1 0 1988 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5447
timestamp 1682952543
transform 1 0 1980 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5331
timestamp 1682952543
transform 1 0 1996 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5367
timestamp 1682952543
transform 1 0 1996 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5308
timestamp 1682952543
transform 1 0 2028 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5423
timestamp 1682952543
transform 1 0 2012 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1682952543
transform 1 0 2028 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1682952543
transform 1 0 2020 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5497
timestamp 1682952543
transform 1 0 2036 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5448
timestamp 1682952543
transform 1 0 2044 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5368
timestamp 1682952543
transform 1 0 2060 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5483
timestamp 1682952543
transform 1 0 2060 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1682952543
transform 1 0 2060 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1682952543
transform 1 0 2068 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5449
timestamp 1682952543
transform 1 0 2068 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5244
timestamp 1682952543
transform 1 0 2092 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5309
timestamp 1682952543
transform 1 0 2084 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5245
timestamp 1682952543
transform 1 0 2124 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5310
timestamp 1682952543
transform 1 0 2116 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5285
timestamp 1682952543
transform 1 0 2204 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1682952543
transform 1 0 2116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1682952543
transform 1 0 2084 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5369
timestamp 1682952543
transform 1 0 2100 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5370
timestamp 1682952543
transform 1 0 2116 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5333
timestamp 1682952543
transform 1 0 2212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1682952543
transform 1 0 2140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5427
timestamp 1682952543
transform 1 0 2196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5484
timestamp 1682952543
transform 1 0 2100 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5424
timestamp 1682952543
transform 1 0 2108 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5425
timestamp 1682952543
transform 1 0 2140 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1682952543
transform 1 0 2268 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5334
timestamp 1682952543
transform 1 0 2252 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5335
timestamp 1682952543
transform 1 0 2268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1682952543
transform 1 0 2220 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1682952543
transform 1 0 2228 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1682952543
transform 1 0 2244 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5426
timestamp 1682952543
transform 1 0 2244 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5371
timestamp 1682952543
transform 1 0 2268 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5431
timestamp 1682952543
transform 1 0 2300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5432
timestamp 1682952543
transform 1 0 2348 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5427
timestamp 1682952543
transform 1 0 2356 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1682952543
transform 1 0 2388 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5433
timestamp 1682952543
transform 1 0 2380 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1682952543
transform 1 0 2396 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5428
timestamp 1682952543
transform 1 0 2380 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5312
timestamp 1682952543
transform 1 0 2428 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5336
timestamp 1682952543
transform 1 0 2428 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5429
timestamp 1682952543
transform 1 0 2420 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5337
timestamp 1682952543
transform 1 0 2444 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5372
timestamp 1682952543
transform 1 0 2444 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5247
timestamp 1682952543
transform 1 0 2540 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5313
timestamp 1682952543
transform 1 0 2532 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5434
timestamp 1682952543
transform 1 0 2468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5435
timestamp 1682952543
transform 1 0 2524 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5430
timestamp 1682952543
transform 1 0 2476 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5431
timestamp 1682952543
transform 1 0 2548 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1682952543
transform 1 0 2564 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5343
timestamp 1682952543
transform 1 0 2564 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5436
timestamp 1682952543
transform 1 0 2564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1682952543
transform 1 0 2580 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1682952543
transform 1 0 2604 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1682952543
transform 1 0 2604 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5338
timestamp 1682952543
transform 1 0 2620 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5438
timestamp 1682952543
transform 1 0 2620 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5249
timestamp 1682952543
transform 1 0 2644 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5339
timestamp 1682952543
transform 1 0 2628 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5344
timestamp 1682952543
transform 1 0 2636 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1682952543
transform 1 0 2628 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5439
timestamp 1682952543
transform 1 0 2644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5440
timestamp 1682952543
transform 1 0 2652 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5250
timestamp 1682952543
transform 1 0 2708 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5251
timestamp 1682952543
transform 1 0 2740 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5314
timestamp 1682952543
transform 1 0 2748 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5340
timestamp 1682952543
transform 1 0 2748 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5345
timestamp 1682952543
transform 1 0 2764 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5374
timestamp 1682952543
transform 1 0 2684 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5441
timestamp 1682952543
transform 1 0 2724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1682952543
transform 1 0 2764 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5398
timestamp 1682952543
transform 1 0 2676 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5399
timestamp 1682952543
transform 1 0 2748 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5286
timestamp 1682952543
transform 1 0 2780 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1682952543
transform 1 0 2780 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5346
timestamp 1682952543
transform 1 0 2804 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5375
timestamp 1682952543
transform 1 0 2780 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5443
timestamp 1682952543
transform 1 0 2804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5488
timestamp 1682952543
transform 1 0 2788 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1682952543
transform 1 0 2796 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1682952543
transform 1 0 2828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1682952543
transform 1 0 2828 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5347
timestamp 1682952543
transform 1 0 2836 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5252
timestamp 1682952543
transform 1 0 2860 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5253
timestamp 1682952543
transform 1 0 2892 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5270
timestamp 1682952543
transform 1 0 2868 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5343
timestamp 1682952543
transform 1 0 2868 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5444
timestamp 1682952543
transform 1 0 2852 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1682952543
transform 1 0 2860 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5446
timestamp 1682952543
transform 1 0 2876 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5400
timestamp 1682952543
transform 1 0 2860 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5315
timestamp 1682952543
transform 1 0 2900 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5447
timestamp 1682952543
transform 1 0 2900 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5401
timestamp 1682952543
transform 1 0 2892 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5316
timestamp 1682952543
transform 1 0 2916 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5448
timestamp 1682952543
transform 1 0 2924 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5271
timestamp 1682952543
transform 1 0 2956 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5317
timestamp 1682952543
transform 1 0 2940 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5318
timestamp 1682952543
transform 1 0 2956 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5344
timestamp 1682952543
transform 1 0 2932 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1682952543
transform 1 0 2940 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1682952543
transform 1 0 2956 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1682952543
transform 1 0 2980 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1682952543
transform 1 0 2948 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1682952543
transform 1 0 2964 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5451
timestamp 1682952543
transform 1 0 2972 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5402
timestamp 1682952543
transform 1 0 2956 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1682952543
transform 1 0 2948 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1682952543
transform 1 0 2972 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5348
timestamp 1682952543
transform 1 0 3028 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5403
timestamp 1682952543
transform 1 0 3028 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1682952543
transform 1 0 3068 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5319
timestamp 1682952543
transform 1 0 3068 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1682952543
transform 1 0 3116 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5348
timestamp 1682952543
transform 1 0 3116 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5452
timestamp 1682952543
transform 1 0 3068 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5404
timestamp 1682952543
transform 1 0 3076 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1682952543
transform 1 0 3052 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5490
timestamp 1682952543
transform 1 0 3140 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5435
timestamp 1682952543
transform 1 0 3140 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5501
timestamp 1682952543
transform 1 0 3156 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5456
timestamp 1682952543
transform 1 0 3156 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5502
timestamp 1682952543
transform 1 0 3188 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5349
timestamp 1682952543
transform 1 0 3204 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5491
timestamp 1682952543
transform 1 0 3204 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5457
timestamp 1682952543
transform 1 0 3204 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5254
timestamp 1682952543
transform 1 0 3276 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5321
timestamp 1682952543
transform 1 0 3220 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5322
timestamp 1682952543
transform 1 0 3268 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5349
timestamp 1682952543
transform 1 0 3220 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1682952543
transform 1 0 3268 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5405
timestamp 1682952543
transform 1 0 3292 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5458
timestamp 1682952543
transform 1 0 3268 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5255
timestamp 1682952543
transform 1 0 3332 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1682952543
transform 1 0 3324 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5436
timestamp 1682952543
transform 1 0 3316 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5256
timestamp 1682952543
transform 1 0 3356 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5274
timestamp 1682952543
transform 1 0 3364 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1682952543
transform 1 0 3364 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5350
timestamp 1682952543
transform 1 0 3348 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1682952543
transform 1 0 3364 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1682952543
transform 1 0 3380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1682952543
transform 1 0 3388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5454
timestamp 1682952543
transform 1 0 3348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5455
timestamp 1682952543
transform 1 0 3356 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1682952543
transform 1 0 3372 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5275
timestamp 1682952543
transform 1 0 3404 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1682952543
transform 1 0 3428 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5350
timestamp 1682952543
transform 1 0 3420 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5354
timestamp 1682952543
transform 1 0 3428 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1682952543
transform 1 0 3396 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1682952543
transform 1 0 3412 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1682952543
transform 1 0 3428 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1682952543
transform 1 0 3436 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5406
timestamp 1682952543
transform 1 0 3396 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1682952543
transform 1 0 3412 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5355
timestamp 1682952543
transform 1 0 3452 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5407
timestamp 1682952543
transform 1 0 3452 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5492
timestamp 1682952543
transform 1 0 3460 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5459
timestamp 1682952543
transform 1 0 3436 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5257
timestamp 1682952543
transform 1 0 3548 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1682952543
transform 1 0 3540 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5356
timestamp 1682952543
transform 1 0 3508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5357
timestamp 1682952543
transform 1 0 3524 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5351
timestamp 1682952543
transform 1 0 3532 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5461
timestamp 1682952543
transform 1 0 3492 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5462
timestamp 1682952543
transform 1 0 3508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5463
timestamp 1682952543
transform 1 0 3532 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5408
timestamp 1682952543
transform 1 0 3484 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5493
timestamp 1682952543
transform 1 0 3500 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1682952543
transform 1 0 3484 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5450
timestamp 1682952543
transform 1 0 3484 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5464
timestamp 1682952543
transform 1 0 3548 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5409
timestamp 1682952543
transform 1 0 3540 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5358
timestamp 1682952543
transform 1 0 3556 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5276
timestamp 1682952543
transform 1 0 3572 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1682952543
transform 1 0 3572 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5352
timestamp 1682952543
transform 1 0 3564 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5410
timestamp 1682952543
transform 1 0 3556 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5451
timestamp 1682952543
transform 1 0 3548 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5359
timestamp 1682952543
transform 1 0 3588 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5411
timestamp 1682952543
transform 1 0 3612 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5353
timestamp 1682952543
transform 1 0 3636 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5376
timestamp 1682952543
transform 1 0 3636 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5465
timestamp 1682952543
transform 1 0 3644 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1682952543
transform 1 0 3628 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5327
timestamp 1682952543
transform 1 0 3716 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5360
timestamp 1682952543
transform 1 0 3668 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5377
timestamp 1682952543
transform 1 0 3668 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5466
timestamp 1682952543
transform 1 0 3716 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5495
timestamp 1682952543
transform 1 0 3652 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1682952543
transform 1 0 3636 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5438
timestamp 1682952543
transform 1 0 3644 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5452
timestamp 1682952543
transform 1 0 3708 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5460
timestamp 1682952543
transform 1 0 3740 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5258
timestamp 1682952543
transform 1 0 3836 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1682952543
transform 1 0 3828 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1682952543
transform 1 0 3852 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5361
timestamp 1682952543
transform 1 0 3828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5362
timestamp 1682952543
transform 1 0 3836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5363
timestamp 1682952543
transform 1 0 3852 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1682952543
transform 1 0 3780 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5468
timestamp 1682952543
transform 1 0 3788 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1682952543
transform 1 0 3804 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5470
timestamp 1682952543
transform 1 0 3820 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5412
timestamp 1682952543
transform 1 0 3780 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1682952543
transform 1 0 3804 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5471
timestamp 1682952543
transform 1 0 3844 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1682952543
transform 1 0 3860 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5259
timestamp 1682952543
transform 1 0 3884 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1682952543
transform 1 0 3908 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1682952543
transform 1 0 3876 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5364
timestamp 1682952543
transform 1 0 3876 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5413
timestamp 1682952543
transform 1 0 3844 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5414
timestamp 1682952543
transform 1 0 3868 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5330
timestamp 1682952543
transform 1 0 3908 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5365
timestamp 1682952543
transform 1 0 3892 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5378
timestamp 1682952543
transform 1 0 3892 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1682952543
transform 1 0 4004 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5331
timestamp 1682952543
transform 1 0 4004 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1682952543
transform 1 0 4044 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5278
timestamp 1682952543
transform 1 0 4028 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5366
timestamp 1682952543
transform 1 0 3988 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1682952543
transform 1 0 4004 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5368
timestamp 1682952543
transform 1 0 4020 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1682952543
transform 1 0 3916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5474
timestamp 1682952543
transform 1 0 3972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1682952543
transform 1 0 3980 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5415
timestamp 1682952543
transform 1 0 3916 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5476
timestamp 1682952543
transform 1 0 4012 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5369
timestamp 1682952543
transform 1 0 4036 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1682952543
transform 1 0 4028 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5279
timestamp 1682952543
transform 1 0 4052 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1682952543
transform 1 0 4132 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1682952543
transform 1 0 4092 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5370
timestamp 1682952543
transform 1 0 4052 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1682952543
transform 1 0 4068 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1682952543
transform 1 0 4092 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1682952543
transform 1 0 4148 0 1 1925
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_44
timestamp 1682952543
transform 1 0 24 0 1 1870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_322
timestamp 1682952543
transform 1 0 72 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_363
timestamp 1682952543
transform -1 0 184 0 -1 1970
box -9 -3 26 105
use AOI22X1  AOI22X1_208
timestamp 1682952543
transform 1 0 184 0 -1 1970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_325
timestamp 1682952543
transform 1 0 224 0 -1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_326
timestamp 1682952543
transform 1 0 320 0 -1 1970
box -8 -3 104 105
use OAI22X1  OAI22X1_221
timestamp 1682952543
transform -1 0 456 0 -1 1970
box -8 -3 46 105
use FILL  FILL_1820
timestamp 1682952543
transform 1 0 456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1682952543
transform 1 0 464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1682952543
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_222
timestamp 1682952543
transform -1 0 520 0 -1 1970
box -8 -3 46 105
use FILL  FILL_1823
timestamp 1682952543
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_327
timestamp 1682952543
transform 1 0 528 0 -1 1970
box -8 -3 104 105
use FILL  FILL_1824
timestamp 1682952543
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1682952543
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_364
timestamp 1682952543
transform -1 0 656 0 -1 1970
box -9 -3 26 105
use FILL  FILL_1827
timestamp 1682952543
transform 1 0 656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1829
timestamp 1682952543
transform 1 0 664 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5461
timestamp 1682952543
transform 1 0 700 0 1 1875
box -3 -3 3 3
use AOI22X1  AOI22X1_209
timestamp 1682952543
transform 1 0 672 0 -1 1970
box -8 -3 46 105
use FILL  FILL_1834
timestamp 1682952543
transform 1 0 712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1682952543
transform 1 0 720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1682952543
transform 1 0 728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1682952543
transform 1 0 736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1682952543
transform 1 0 744 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_63
timestamp 1682952543
transform 1 0 752 0 -1 1970
box -8 -3 32 105
use FILL  FILL_1845
timestamp 1682952543
transform 1 0 776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1682952543
transform 1 0 784 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_64
timestamp 1682952543
transform 1 0 792 0 -1 1970
box -8 -3 32 105
use FILL  FILL_1847
timestamp 1682952543
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1682952543
transform 1 0 824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1682952543
transform 1 0 832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1682952543
transform 1 0 840 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_65
timestamp 1682952543
transform 1 0 848 0 -1 1970
box -8 -3 32 105
use M3_M2  M3_M2_5462
timestamp 1682952543
transform 1 0 908 0 1 1875
box -3 -3 3 3
use AOI22X1  AOI22X1_212
timestamp 1682952543
transform 1 0 872 0 -1 1970
box -8 -3 46 105
use FILL  FILL_1858
timestamp 1682952543
transform 1 0 912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1860
timestamp 1682952543
transform 1 0 920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1682952543
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1682952543
transform 1 0 936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1682952543
transform 1 0 944 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_214
timestamp 1682952543
transform -1 0 992 0 -1 1970
box -8 -3 46 105
use FILL  FILL_1870
timestamp 1682952543
transform 1 0 992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1871
timestamp 1682952543
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1682952543
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1682952543
transform 1 0 1016 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1682952543
transform 1 0 1024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1682952543
transform 1 0 1032 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1682952543
transform 1 0 1040 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_365
timestamp 1682952543
transform 1 0 1048 0 -1 1970
box -9 -3 26 105
use OAI21X1  OAI21X1_70
timestamp 1682952543
transform -1 0 1096 0 -1 1970
box -8 -3 34 105
use FILL  FILL_1886
timestamp 1682952543
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1682952543
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1888
timestamp 1682952543
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1682952543
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1682952543
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1894
timestamp 1682952543
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5463
timestamp 1682952543
transform 1 0 1172 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5464
timestamp 1682952543
transform 1 0 1204 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_328
timestamp 1682952543
transform 1 0 1144 0 -1 1970
box -8 -3 104 105
use FILL  FILL_1904
timestamp 1682952543
transform 1 0 1240 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_366
timestamp 1682952543
transform 1 0 1248 0 -1 1970
box -9 -3 26 105
use FILL  FILL_1908
timestamp 1682952543
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1682952543
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1682952543
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_224
timestamp 1682952543
transform -1 0 1328 0 -1 1970
box -8 -3 46 105
use FILL  FILL_1914
timestamp 1682952543
transform 1 0 1328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1682952543
transform 1 0 1336 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5465
timestamp 1682952543
transform 1 0 1356 0 1 1875
box -3 -3 3 3
use FILL  FILL_1920
timestamp 1682952543
transform 1 0 1344 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_226
timestamp 1682952543
transform -1 0 1392 0 -1 1970
box -8 -3 46 105
use M3_M2  M3_M2_5466
timestamp 1682952543
transform 1 0 1404 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_368
timestamp 1682952543
transform -1 0 1408 0 -1 1970
box -9 -3 26 105
use M3_M2  M3_M2_5467
timestamp 1682952543
transform 1 0 1428 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1682952543
transform 1 0 1476 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_331
timestamp 1682952543
transform -1 0 1504 0 -1 1970
box -8 -3 104 105
use BUFX2  BUFX2_70
timestamp 1682952543
transform 1 0 1504 0 -1 1970
box -5 -3 28 105
use FILL  FILL_1921
timestamp 1682952543
transform 1 0 1528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1682952543
transform 1 0 1536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1682952543
transform 1 0 1544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1682952543
transform 1 0 1552 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_71
timestamp 1682952543
transform -1 0 1584 0 -1 1970
box -5 -3 28 105
use FILL  FILL_1925
timestamp 1682952543
transform 1 0 1584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1682952543
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_72
timestamp 1682952543
transform 1 0 1600 0 -1 1970
box -5 -3 28 105
use FILL  FILL_1927
timestamp 1682952543
transform 1 0 1624 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_73
timestamp 1682952543
transform -1 0 1656 0 -1 1970
box -5 -3 28 105
use M3_M2  M3_M2_5469
timestamp 1682952543
transform 1 0 1668 0 1 1875
box -3 -3 3 3
use FILL  FILL_1928
timestamp 1682952543
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1682952543
transform 1 0 1664 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_228
timestamp 1682952543
transform -1 0 1712 0 -1 1970
box -8 -3 46 105
use FILL  FILL_1933
timestamp 1682952543
transform 1 0 1712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1682952543
transform 1 0 1720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1936
timestamp 1682952543
transform 1 0 1728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1682952543
transform 1 0 1736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1682952543
transform 1 0 1744 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5470
timestamp 1682952543
transform 1 0 1780 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_369
timestamp 1682952543
transform 1 0 1752 0 -1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_332
timestamp 1682952543
transform 1 0 1768 0 -1 1970
box -8 -3 104 105
use FILL  FILL_1948
timestamp 1682952543
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1682952543
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5471
timestamp 1682952543
transform 1 0 1892 0 1 1875
box -3 -3 3 3
use BUFX2  BUFX2_75
timestamp 1682952543
transform 1 0 1880 0 -1 1970
box -5 -3 28 105
use FILL  FILL_1951
timestamp 1682952543
transform 1 0 1904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1682952543
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1682952543
transform 1 0 1920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1956
timestamp 1682952543
transform 1 0 1928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1682952543
transform 1 0 1936 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_36
timestamp 1682952543
transform -1 0 1976 0 -1 1970
box -8 -3 40 105
use M3_M2  M3_M2_5472
timestamp 1682952543
transform 1 0 1988 0 1 1875
box -3 -3 3 3
use FILL  FILL_1962
timestamp 1682952543
transform 1 0 1976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1682952543
transform 1 0 1984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1682952543
transform 1 0 1992 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_371
timestamp 1682952543
transform 1 0 2000 0 -1 1970
box -9 -3 26 105
use NAND3X1  NAND3X1_37
timestamp 1682952543
transform 1 0 2016 0 -1 1970
box -8 -3 40 105
use FILL  FILL_1979
timestamp 1682952543
transform 1 0 2048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1682952543
transform 1 0 2056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1981
timestamp 1682952543
transform 1 0 2064 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_38
timestamp 1682952543
transform 1 0 2072 0 -1 1970
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_335
timestamp 1682952543
transform 1 0 2104 0 -1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5473
timestamp 1682952543
transform 1 0 2212 0 1 1875
box -3 -3 3 3
use NOR2X1  NOR2X1_69
timestamp 1682952543
transform 1 0 2200 0 -1 1970
box -8 -3 32 105
use AND2X2  AND2X2_46
timestamp 1682952543
transform -1 0 2256 0 -1 1970
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_336
timestamp 1682952543
transform 1 0 2256 0 -1 1970
box -8 -3 104 105
use FILL  FILL_1982
timestamp 1682952543
transform 1 0 2352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1682952543
transform 1 0 2360 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_72
timestamp 1682952543
transform 1 0 2368 0 -1 1970
box -8 -3 34 105
use FILL  FILL_1984
timestamp 1682952543
transform 1 0 2400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1985
timestamp 1682952543
transform 1 0 2408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1682952543
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1987
timestamp 1682952543
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_337
timestamp 1682952543
transform 1 0 2432 0 -1 1970
box -8 -3 104 105
use FILL  FILL_1988
timestamp 1682952543
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1682952543
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1682952543
transform 1 0 2544 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_73
timestamp 1682952543
transform 1 0 2552 0 -1 1970
box -8 -3 34 105
use FILL  FILL_1991
timestamp 1682952543
transform 1 0 2584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1682952543
transform 1 0 2592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1993
timestamp 1682952543
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1682952543
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1682952543
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_74
timestamp 1682952543
transform -1 0 2656 0 -1 1970
box -8 -3 34 105
use FILL  FILL_2004
timestamp 1682952543
transform 1 0 2656 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_340
timestamp 1682952543
transform -1 0 2760 0 -1 1970
box -8 -3 104 105
use NOR2X1  NOR2X1_71
timestamp 1682952543
transform -1 0 2784 0 -1 1970
box -8 -3 32 105
use M3_M2  M3_M2_5474
timestamp 1682952543
transform 1 0 2796 0 1 1875
box -3 -3 3 3
use NAND3X1  NAND3X1_39
timestamp 1682952543
transform -1 0 2816 0 -1 1970
box -8 -3 40 105
use FILL  FILL_2005
timestamp 1682952543
transform 1 0 2816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1682952543
transform 1 0 2824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1682952543
transform 1 0 2832 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_372
timestamp 1682952543
transform 1 0 2840 0 -1 1970
box -9 -3 26 105
use AOI22X1  AOI22X1_215
timestamp 1682952543
transform -1 0 2896 0 -1 1970
box -8 -3 46 105
use FILL  FILL_2008
timestamp 1682952543
transform 1 0 2896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2009
timestamp 1682952543
transform 1 0 2904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1682952543
transform 1 0 2912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1682952543
transform 1 0 2920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2015
timestamp 1682952543
transform 1 0 2928 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_237
timestamp 1682952543
transform -1 0 2976 0 -1 1970
box -8 -3 46 105
use FILL  FILL_2016
timestamp 1682952543
transform 1 0 2976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1682952543
transform 1 0 2984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1682952543
transform 1 0 2992 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_373
timestamp 1682952543
transform -1 0 3016 0 -1 1970
box -9 -3 26 105
use FILL  FILL_2029
timestamp 1682952543
transform 1 0 3016 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5475
timestamp 1682952543
transform 1 0 3036 0 1 1875
box -3 -3 3 3
use FILL  FILL_2030
timestamp 1682952543
transform 1 0 3024 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5476
timestamp 1682952543
transform 1 0 3060 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_341
timestamp 1682952543
transform -1 0 3128 0 -1 1970
box -8 -3 104 105
use FILL  FILL_2031
timestamp 1682952543
transform 1 0 3128 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5477
timestamp 1682952543
transform 1 0 3148 0 1 1875
box -3 -3 3 3
use FILL  FILL_2034
timestamp 1682952543
transform 1 0 3136 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_43
timestamp 1682952543
transform -1 0 3176 0 -1 1970
box -8 -3 40 105
use FILL  FILL_2035
timestamp 1682952543
transform 1 0 3176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1682952543
transform 1 0 3184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1682952543
transform 1 0 3192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1682952543
transform 1 0 3200 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5478
timestamp 1682952543
transform 1 0 3244 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_342
timestamp 1682952543
transform 1 0 3208 0 -1 1970
box -8 -3 104 105
use FILL  FILL_2042
timestamp 1682952543
transform 1 0 3304 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_378
timestamp 1682952543
transform 1 0 3312 0 -1 1970
box -9 -3 26 105
use FILL  FILL_2056
timestamp 1682952543
transform 1 0 3328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1682952543
transform 1 0 3336 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_242
timestamp 1682952543
transform 1 0 3344 0 -1 1970
box -8 -3 46 105
use FILL  FILL_2058
timestamp 1682952543
transform 1 0 3384 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_219
timestamp 1682952543
transform 1 0 3392 0 -1 1970
box -8 -3 46 105
use BUFX2  BUFX2_79
timestamp 1682952543
transform 1 0 3432 0 -1 1970
box -5 -3 28 105
use FILL  FILL_2059
timestamp 1682952543
transform 1 0 3456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1682952543
transform 1 0 3464 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5479
timestamp 1682952543
transform 1 0 3500 0 1 1875
box -3 -3 3 3
use NAND3X1  NAND3X1_46
timestamp 1682952543
transform -1 0 3504 0 -1 1970
box -8 -3 40 105
use OAI22X1  OAI22X1_243
timestamp 1682952543
transform 1 0 3504 0 -1 1970
box -8 -3 46 105
use FILL  FILL_2061
timestamp 1682952543
transform 1 0 3544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1682952543
transform 1 0 3552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1682952543
transform 1 0 3560 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_379
timestamp 1682952543
transform -1 0 3584 0 -1 1970
box -9 -3 26 105
use FILL  FILL_2064
timestamp 1682952543
transform 1 0 3584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1682952543
transform 1 0 3592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1682952543
transform 1 0 3600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2067
timestamp 1682952543
transform 1 0 3608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1682952543
transform 1 0 3616 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_47
timestamp 1682952543
transform -1 0 3656 0 -1 1970
box -8 -3 40 105
use M3_M2  M3_M2_5480
timestamp 1682952543
transform 1 0 3676 0 1 1875
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1682952543
transform 1 0 3692 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_347
timestamp 1682952543
transform 1 0 3656 0 -1 1970
box -8 -3 104 105
use M3_M2  M3_M2_5482
timestamp 1682952543
transform 1 0 3764 0 1 1875
box -3 -3 3 3
use FILL  FILL_2069
timestamp 1682952543
transform 1 0 3752 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_380
timestamp 1682952543
transform 1 0 3760 0 -1 1970
box -9 -3 26 105
use FILL  FILL_2070
timestamp 1682952543
transform 1 0 3776 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_220
timestamp 1682952543
transform -1 0 3824 0 -1 1970
box -8 -3 46 105
use FILL  FILL_2071
timestamp 1682952543
transform 1 0 3824 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_244
timestamp 1682952543
transform -1 0 3872 0 -1 1970
box -8 -3 46 105
use FILL  FILL_2072
timestamp 1682952543
transform 1 0 3872 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_348
timestamp 1682952543
transform 1 0 3880 0 -1 1970
box -8 -3 104 105
use FILL  FILL_2073
timestamp 1682952543
transform 1 0 3976 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_245
timestamp 1682952543
transform 1 0 3984 0 -1 1970
box -8 -3 46 105
use FILL  FILL_2074
timestamp 1682952543
transform 1 0 4024 0 -1 1970
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1682952543
transform 1 0 4032 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_381
timestamp 1682952543
transform -1 0 4056 0 -1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_349
timestamp 1682952543
transform 1 0 4056 0 -1 1970
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_45
timestamp 1682952543
transform 1 0 4201 0 1 1870
box -10 -3 10 3
use M3_M2  M3_M2_5527
timestamp 1682952543
transform 1 0 164 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5549
timestamp 1682952543
transform 1 0 116 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5550
timestamp 1682952543
transform 1 0 172 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5537
timestamp 1682952543
transform 1 0 116 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1682952543
transform 1 0 164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5539
timestamp 1682952543
transform 1 0 172 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5639
timestamp 1682952543
transform 1 0 84 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5551
timestamp 1682952543
transform 1 0 204 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5540
timestamp 1682952543
transform 1 0 204 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5528
timestamp 1682952543
transform 1 0 220 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5541
timestamp 1682952543
transform 1 0 228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1682952543
transform 1 0 212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1682952543
transform 1 0 220 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5639
timestamp 1682952543
transform 1 0 204 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5640
timestamp 1682952543
transform 1 0 228 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5542
timestamp 1682952543
transform 1 0 252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1682952543
transform 1 0 268 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5642
timestamp 1682952543
transform 1 0 260 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5606
timestamp 1682952543
transform 1 0 260 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5552
timestamp 1682952543
transform 1 0 292 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5544
timestamp 1682952543
transform 1 0 292 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5641
timestamp 1682952543
transform 1 0 284 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5553
timestamp 1682952543
transform 1 0 308 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1682952543
transform 1 0 332 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5555
timestamp 1682952543
transform 1 0 348 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5545
timestamp 1682952543
transform 1 0 332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1682952543
transform 1 0 348 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5564
timestamp 1682952543
transform 1 0 356 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5547
timestamp 1682952543
transform 1 0 364 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5643
timestamp 1682952543
transform 1 0 316 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5644
timestamp 1682952543
transform 1 0 324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1682952543
transform 1 0 340 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5583
timestamp 1682952543
transform 1 0 348 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5607
timestamp 1682952543
transform 1 0 340 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5642
timestamp 1682952543
transform 1 0 324 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5556
timestamp 1682952543
transform 1 0 388 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5565
timestamp 1682952543
transform 1 0 380 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5548
timestamp 1682952543
transform 1 0 388 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5584
timestamp 1682952543
transform 1 0 372 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1682952543
transform 1 0 380 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1682952543
transform 1 0 444 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5549
timestamp 1682952543
transform 1 0 420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5550
timestamp 1682952543
transform 1 0 436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5646
timestamp 1682952543
transform 1 0 404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1682952543
transform 1 0 412 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1682952543
transform 1 0 428 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5609
timestamp 1682952543
transform 1 0 396 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5610
timestamp 1682952543
transform 1 0 412 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5649
timestamp 1682952543
transform 1 0 444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5551
timestamp 1682952543
transform 1 0 476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5552
timestamp 1682952543
transform 1 0 508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1682952543
transform 1 0 484 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5651
timestamp 1682952543
transform 1 0 500 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5505
timestamp 1682952543
transform 1 0 604 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5557
timestamp 1682952543
transform 1 0 580 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5553
timestamp 1682952543
transform 1 0 580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5554
timestamp 1682952543
transform 1 0 612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1682952543
transform 1 0 532 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5643
timestamp 1682952543
transform 1 0 612 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5558
timestamp 1682952543
transform 1 0 628 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5555
timestamp 1682952543
transform 1 0 628 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5566
timestamp 1682952543
transform 1 0 644 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5611
timestamp 1682952543
transform 1 0 636 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1682952543
transform 1 0 660 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5529
timestamp 1682952543
transform 1 0 660 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5556
timestamp 1682952543
transform 1 0 660 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5567
timestamp 1682952543
transform 1 0 676 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5557
timestamp 1682952543
transform 1 0 684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5653
timestamp 1682952543
transform 1 0 668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1682952543
transform 1 0 676 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5655
timestamp 1682952543
transform 1 0 692 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5644
timestamp 1682952543
transform 1 0 692 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5656
timestamp 1682952543
transform 1 0 708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5558
timestamp 1682952543
transform 1 0 724 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5530
timestamp 1682952543
transform 1 0 756 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5559
timestamp 1682952543
transform 1 0 772 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5559
timestamp 1682952543
transform 1 0 756 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5531
timestamp 1682952543
transform 1 0 796 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5516
timestamp 1682952543
transform 1 0 804 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1682952543
transform 1 0 796 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5568
timestamp 1682952543
transform 1 0 804 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5657
timestamp 1682952543
transform 1 0 788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1682952543
transform 1 0 796 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5645
timestamp 1682952543
transform 1 0 796 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5561
timestamp 1682952543
transform 1 0 820 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5585
timestamp 1682952543
transform 1 0 820 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5586
timestamp 1682952543
transform 1 0 836 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5505
timestamp 1682952543
transform 1 0 860 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_5659
timestamp 1682952543
transform 1 0 852 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1682952543
transform 1 0 900 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5587
timestamp 1682952543
transform 1 0 900 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5506
timestamp 1682952543
transform 1 0 908 0 1 1855
box -2 -2 2 2
use M3_M2  M3_M2_5532
timestamp 1682952543
transform 1 0 932 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5562
timestamp 1682952543
transform 1 0 932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5563
timestamp 1682952543
transform 1 0 948 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5660
timestamp 1682952543
transform 1 0 916 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5661
timestamp 1682952543
transform 1 0 924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1682952543
transform 1 0 940 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5506
timestamp 1682952543
transform 1 0 972 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5507
timestamp 1682952543
transform 1 0 1036 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5564
timestamp 1682952543
transform 1 0 1020 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5663
timestamp 1682952543
transform 1 0 972 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5612
timestamp 1682952543
transform 1 0 988 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1682952543
transform 1 0 1020 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1682952543
transform 1 0 1060 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5518
timestamp 1682952543
transform 1 0 1068 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5565
timestamp 1682952543
transform 1 0 1060 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5569
timestamp 1682952543
transform 1 0 1068 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5664
timestamp 1682952543
transform 1 0 1068 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5734
timestamp 1682952543
transform 1 0 1068 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5509
timestamp 1682952543
transform 1 0 1092 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5735
timestamp 1682952543
transform 1 0 1084 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1682952543
transform 1 0 1116 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1682952543
transform 1 0 1164 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5566
timestamp 1682952543
transform 1 0 1172 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5614
timestamp 1682952543
transform 1 0 1172 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5521
timestamp 1682952543
transform 1 0 1188 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5570
timestamp 1682952543
transform 1 0 1188 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1682952543
transform 1 0 1204 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5567
timestamp 1682952543
transform 1 0 1204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1682952543
transform 1 0 1188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1682952543
transform 1 0 1196 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1682952543
transform 1 0 1212 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5668
timestamp 1682952543
transform 1 0 1228 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1682952543
transform 1 0 1236 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5615
timestamp 1682952543
transform 1 0 1228 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1682952543
transform 1 0 1212 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5588
timestamp 1682952543
transform 1 0 1244 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5511
timestamp 1682952543
transform 1 0 1260 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5568
timestamp 1682952543
transform 1 0 1260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1682952543
transform 1 0 1260 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5512
timestamp 1682952543
transform 1 0 1316 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5569
timestamp 1682952543
transform 1 0 1316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1682952543
transform 1 0 1356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1682952543
transform 1 0 1276 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5616
timestamp 1682952543
transform 1 0 1324 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5513
timestamp 1682952543
transform 1 0 1396 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5571
timestamp 1682952543
transform 1 0 1372 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5571
timestamp 1682952543
transform 1 0 1380 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5572
timestamp 1682952543
transform 1 0 1396 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5672
timestamp 1682952543
transform 1 0 1364 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5589
timestamp 1682952543
transform 1 0 1380 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5673
timestamp 1682952543
transform 1 0 1388 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5514
timestamp 1682952543
transform 1 0 1412 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5573
timestamp 1682952543
transform 1 0 1412 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5590
timestamp 1682952543
transform 1 0 1412 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5736
timestamp 1682952543
transform 1 0 1412 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5574
timestamp 1682952543
transform 1 0 1492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1682952543
transform 1 0 1484 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5647
timestamp 1682952543
transform 1 0 1484 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5675
timestamp 1682952543
transform 1 0 1508 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5648
timestamp 1682952543
transform 1 0 1524 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5575
timestamp 1682952543
transform 1 0 1564 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1682952543
transform 1 0 1540 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5677
timestamp 1682952543
transform 1 0 1556 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5649
timestamp 1682952543
transform 1 0 1540 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1682952543
transform 1 0 1676 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_5576
timestamp 1682952543
transform 1 0 1588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5577
timestamp 1682952543
transform 1 0 1636 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5678
timestamp 1682952543
transform 1 0 1580 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5679
timestamp 1682952543
transform 1 0 1668 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5617
timestamp 1682952543
transform 1 0 1628 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5650
timestamp 1682952543
transform 1 0 1596 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1682952543
transform 1 0 1700 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5737
timestamp 1682952543
transform 1 0 1692 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1682952543
transform 1 0 1708 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5651
timestamp 1682952543
transform 1 0 1700 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5579
timestamp 1682952543
transform 1 0 1724 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5487
timestamp 1682952543
transform 1 0 1740 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5572
timestamp 1682952543
transform 1 0 1748 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1682952543
transform 1 0 1780 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5515
timestamp 1682952543
transform 1 0 1764 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5516
timestamp 1682952543
transform 1 0 1796 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5580
timestamp 1682952543
transform 1 0 1772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5581
timestamp 1682952543
transform 1 0 1788 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1682952543
transform 1 0 1748 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1682952543
transform 1 0 1756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1682952543
transform 1 0 1796 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5738
timestamp 1682952543
transform 1 0 1812 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5517
timestamp 1682952543
transform 1 0 1860 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5582
timestamp 1682952543
transform 1 0 1852 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5560
timestamp 1682952543
transform 1 0 1868 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5583
timestamp 1682952543
transform 1 0 1876 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5683
timestamp 1682952543
transform 1 0 1868 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5618
timestamp 1682952543
transform 1 0 1860 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1682952543
transform 1 0 1868 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5591
timestamp 1682952543
transform 1 0 1884 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5684
timestamp 1682952543
transform 1 0 1892 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1682952543
transform 1 0 1900 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5619
timestamp 1682952543
transform 1 0 1884 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1682952543
transform 1 0 2012 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5584
timestamp 1682952543
transform 1 0 1924 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1682952543
transform 1 0 1932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5586
timestamp 1682952543
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5592
timestamp 1682952543
transform 1 0 1924 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1682952543
transform 1 0 1964 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5686
timestamp 1682952543
transform 1 0 2012 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5518
timestamp 1682952543
transform 1 0 2036 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5739
timestamp 1682952543
transform 1 0 2028 0 1 1795
box -2 -2 2 2
use M3_M2  M3_M2_5519
timestamp 1682952543
transform 1 0 2060 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5587
timestamp 1682952543
transform 1 0 2060 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5520
timestamp 1682952543
transform 1 0 2076 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5687
timestamp 1682952543
transform 1 0 2076 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5688
timestamp 1682952543
transform 1 0 2092 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5620
timestamp 1682952543
transform 1 0 2092 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1682952543
transform 1 0 2116 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5491
timestamp 1682952543
transform 1 0 2140 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5588
timestamp 1682952543
transform 1 0 2108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1682952543
transform 1 0 2116 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5590
timestamp 1682952543
transform 1 0 2132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5689
timestamp 1682952543
transform 1 0 2116 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5621
timestamp 1682952543
transform 1 0 2132 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5653
timestamp 1682952543
transform 1 0 2116 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5492
timestamp 1682952543
transform 1 0 2156 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5533
timestamp 1682952543
transform 1 0 2156 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5591
timestamp 1682952543
transform 1 0 2156 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5594
timestamp 1682952543
transform 1 0 2156 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5534
timestamp 1682952543
transform 1 0 2204 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5522
timestamp 1682952543
transform 1 0 2212 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5592
timestamp 1682952543
transform 1 0 2196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1682952543
transform 1 0 2188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1682952543
transform 1 0 2220 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5535
timestamp 1682952543
transform 1 0 2252 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5593
timestamp 1682952543
transform 1 0 2252 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1682952543
transform 1 0 2252 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5654
timestamp 1682952543
transform 1 0 2252 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5523
timestamp 1682952543
transform 1 0 2276 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1682952543
transform 1 0 2292 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5655
timestamp 1682952543
transform 1 0 2284 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5594
timestamp 1682952543
transform 1 0 2300 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5595
timestamp 1682952543
transform 1 0 2316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5596
timestamp 1682952543
transform 1 0 2340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1682952543
transform 1 0 2324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1682952543
transform 1 0 2332 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1682952543
transform 1 0 2348 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5622
timestamp 1682952543
transform 1 0 2332 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1682952543
transform 1 0 2340 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5597
timestamp 1682952543
transform 1 0 2364 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5595
timestamp 1682952543
transform 1 0 2364 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5697
timestamp 1682952543
transform 1 0 2388 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5524
timestamp 1682952543
transform 1 0 2404 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1682952543
transform 1 0 2420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5599
timestamp 1682952543
transform 1 0 2468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5600
timestamp 1682952543
transform 1 0 2476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5698
timestamp 1682952543
transform 1 0 2452 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5699
timestamp 1682952543
transform 1 0 2460 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5623
timestamp 1682952543
transform 1 0 2460 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5596
timestamp 1682952543
transform 1 0 2476 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5601
timestamp 1682952543
transform 1 0 2500 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1682952543
transform 1 0 2516 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5602
timestamp 1682952543
transform 1 0 2540 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5603
timestamp 1682952543
transform 1 0 2556 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5701
timestamp 1682952543
transform 1 0 2556 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5624
timestamp 1682952543
transform 1 0 2540 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5657
timestamp 1682952543
transform 1 0 2556 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5604
timestamp 1682952543
transform 1 0 2628 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1682952543
transform 1 0 2644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1682952543
transform 1 0 2652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5703
timestamp 1682952543
transform 1 0 2660 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5704
timestamp 1682952543
transform 1 0 2668 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5625
timestamp 1682952543
transform 1 0 2644 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1682952543
transform 1 0 2668 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5507
timestamp 1682952543
transform 1 0 2692 0 1 1855
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1682952543
transform 1 0 2708 0 1 1855
box -2 -2 2 2
use M3_M2  M3_M2_5493
timestamp 1682952543
transform 1 0 2732 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5509
timestamp 1682952543
transform 1 0 2732 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5606
timestamp 1682952543
transform 1 0 2724 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1682952543
transform 1 0 2796 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1682952543
transform 1 0 2812 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1682952543
transform 1 0 2820 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5705
timestamp 1682952543
transform 1 0 2796 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1682952543
transform 1 0 2868 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1682952543
transform 1 0 2884 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1682952543
transform 1 0 2892 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5627
timestamp 1682952543
transform 1 0 2884 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5607
timestamp 1682952543
transform 1 0 2924 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5597
timestamp 1682952543
transform 1 0 2932 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5536
timestamp 1682952543
transform 1 0 2948 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1682952543
transform 1 0 2948 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5494
timestamp 1682952543
transform 1 0 3036 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1682952543
transform 1 0 3116 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5537
timestamp 1682952543
transform 1 0 2988 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1682952543
transform 1 0 3044 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1682952543
transform 1 0 3100 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5608
timestamp 1682952543
transform 1 0 2988 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5598
timestamp 1682952543
transform 1 0 2988 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5706
timestamp 1682952543
transform 1 0 3036 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5609
timestamp 1682952543
transform 1 0 3108 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1682952543
transform 1 0 3060 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5540
timestamp 1682952543
transform 1 0 3164 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5610
timestamp 1682952543
transform 1 0 3156 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5611
timestamp 1682952543
transform 1 0 3164 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5496
timestamp 1682952543
transform 1 0 3252 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5541
timestamp 1682952543
transform 1 0 3204 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5542
timestamp 1682952543
transform 1 0 3252 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5612
timestamp 1682952543
transform 1 0 3228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1682952543
transform 1 0 3252 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5497
timestamp 1682952543
transform 1 0 3276 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5529
timestamp 1682952543
transform 1 0 3268 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5543
timestamp 1682952543
transform 1 0 3284 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5512
timestamp 1682952543
transform 1 0 3300 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_5573
timestamp 1682952543
transform 1 0 3300 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5613
timestamp 1682952543
transform 1 0 3308 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1682952543
transform 1 0 3340 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1682952543
transform 1 0 3332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1682952543
transform 1 0 3372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1682952543
transform 1 0 3348 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5599
timestamp 1682952543
transform 1 0 3356 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5710
timestamp 1682952543
transform 1 0 3364 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5629
timestamp 1682952543
transform 1 0 3364 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5711
timestamp 1682952543
transform 1 0 3388 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5498
timestamp 1682952543
transform 1 0 3468 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1682952543
transform 1 0 3404 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5545
timestamp 1682952543
transform 1 0 3524 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5616
timestamp 1682952543
transform 1 0 3428 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5574
timestamp 1682952543
transform 1 0 3444 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5617
timestamp 1682952543
transform 1 0 3484 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5575
timestamp 1682952543
transform 1 0 3492 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5618
timestamp 1682952543
transform 1 0 3500 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5576
timestamp 1682952543
transform 1 0 3508 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5619
timestamp 1682952543
transform 1 0 3516 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1682952543
transform 1 0 3532 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5484
timestamp 1682952543
transform 1 0 3556 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1682952543
transform 1 0 3572 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5500
timestamp 1682952543
transform 1 0 3652 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5513
timestamp 1682952543
transform 1 0 3556 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1682952543
transform 1 0 3548 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1682952543
transform 1 0 3404 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1682952543
transform 1 0 3492 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1682952543
transform 1 0 3508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1682952543
transform 1 0 3524 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5630
timestamp 1682952543
transform 1 0 3428 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5631
timestamp 1682952543
transform 1 0 3492 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1682952543
transform 1 0 3396 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5600
timestamp 1682952543
transform 1 0 3532 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1682952543
transform 1 0 3612 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5532
timestamp 1682952543
transform 1 0 3572 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5577
timestamp 1682952543
transform 1 0 3572 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5521
timestamp 1682952543
transform 1 0 3684 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5514
timestamp 1682952543
transform 1 0 3684 0 1 1835
box -2 -2 2 2
use M3_M2  M3_M2_5547
timestamp 1682952543
transform 1 0 3692 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5533
timestamp 1682952543
transform 1 0 3676 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5621
timestamp 1682952543
transform 1 0 3580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5622
timestamp 1682952543
transform 1 0 3612 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1682952543
transform 1 0 3540 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5717
timestamp 1682952543
transform 1 0 3564 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5632
timestamp 1682952543
transform 1 0 3524 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5659
timestamp 1682952543
transform 1 0 3516 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1682952543
transform 1 0 3564 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5718
timestamp 1682952543
transform 1 0 3660 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5633
timestamp 1682952543
transform 1 0 3620 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5661
timestamp 1682952543
transform 1 0 3612 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_5515
timestamp 1682952543
transform 1 0 3716 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1682952543
transform 1 0 3700 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5535
timestamp 1682952543
transform 1 0 3708 0 1 1825
box -2 -2 2 2
use M3_M2  M3_M2_5561
timestamp 1682952543
transform 1 0 3716 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5536
timestamp 1682952543
transform 1 0 3732 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5623
timestamp 1682952543
transform 1 0 3692 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5578
timestamp 1682952543
transform 1 0 3708 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5624
timestamp 1682952543
transform 1 0 3724 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1682952543
transform 1 0 3740 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5601
timestamp 1682952543
transform 1 0 3724 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5719
timestamp 1682952543
transform 1 0 3772 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5522
timestamp 1682952543
transform 1 0 3788 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5626
timestamp 1682952543
transform 1 0 3788 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5634
timestamp 1682952543
transform 1 0 3780 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5662
timestamp 1682952543
transform 1 0 3772 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1682952543
transform 1 0 3796 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5627
timestamp 1682952543
transform 1 0 3804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5628
timestamp 1682952543
transform 1 0 3820 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1682952543
transform 1 0 3796 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5602
timestamp 1682952543
transform 1 0 3804 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5663
timestamp 1682952543
transform 1 0 3820 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1682952543
transform 1 0 3836 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5502
timestamp 1682952543
transform 1 0 3852 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5580
timestamp 1682952543
transform 1 0 3844 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1682952543
transform 1 0 3900 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5524
timestamp 1682952543
transform 1 0 3924 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5548
timestamp 1682952543
transform 1 0 3916 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5562
timestamp 1682952543
transform 1 0 3892 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5629
timestamp 1682952543
transform 1 0 3860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5630
timestamp 1682952543
transform 1 0 3876 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5563
timestamp 1682952543
transform 1 0 3940 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5631
timestamp 1682952543
transform 1 0 3900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5632
timestamp 1682952543
transform 1 0 3916 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1682952543
transform 1 0 3940 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1682952543
transform 1 0 3844 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5722
timestamp 1682952543
transform 1 0 3852 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1682952543
transform 1 0 3868 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1682952543
transform 1 0 3884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5725
timestamp 1682952543
transform 1 0 3892 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5635
timestamp 1682952543
transform 1 0 3844 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5603
timestamp 1682952543
transform 1 0 3900 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5726
timestamp 1682952543
transform 1 0 3924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5727
timestamp 1682952543
transform 1 0 3932 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5664
timestamp 1682952543
transform 1 0 3932 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1682952543
transform 1 0 3988 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5634
timestamp 1682952543
transform 1 0 3980 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1682952543
transform 1 0 3972 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5525
timestamp 1682952543
transform 1 0 4012 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1682952543
transform 1 0 4004 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5635
timestamp 1682952543
transform 1 0 4012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5729
timestamp 1682952543
transform 1 0 3988 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5730
timestamp 1682952543
transform 1 0 4004 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5604
timestamp 1682952543
transform 1 0 4012 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5731
timestamp 1682952543
transform 1 0 4020 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5636
timestamp 1682952543
transform 1 0 3988 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5526
timestamp 1682952543
transform 1 0 4140 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5636
timestamp 1682952543
transform 1 0 4076 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5582
timestamp 1682952543
transform 1 0 4124 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5637
timestamp 1682952543
transform 1 0 4132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5638
timestamp 1682952543
transform 1 0 4140 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5732
timestamp 1682952543
transform 1 0 4052 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5605
timestamp 1682952543
transform 1 0 4076 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5637
timestamp 1682952543
transform 1 0 4076 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5733
timestamp 1682952543
transform 1 0 4148 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5638
timestamp 1682952543
transform 1 0 4156 0 1 1795
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_46
timestamp 1682952543
transform 1 0 48 0 1 1770
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_350
timestamp 1682952543
transform 1 0 72 0 1 1770
box -8 -3 104 105
use FILL  FILL_2076
timestamp 1682952543
transform 1 0 168 0 1 1770
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1682952543
transform 1 0 176 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_382
timestamp 1682952543
transform -1 0 200 0 1 1770
box -9 -3 26 105
use FILL  FILL_2078
timestamp 1682952543
transform 1 0 200 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_221
timestamp 1682952543
transform -1 0 248 0 1 1770
box -8 -3 46 105
use FILL  FILL_2079
timestamp 1682952543
transform 1 0 248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2080
timestamp 1682952543
transform 1 0 256 0 1 1770
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1682952543
transform 1 0 264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1682952543
transform 1 0 272 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_383
timestamp 1682952543
transform -1 0 296 0 1 1770
box -9 -3 26 105
use FILL  FILL_2083
timestamp 1682952543
transform 1 0 296 0 1 1770
box -8 -3 16 105
use FILL  FILL_2084
timestamp 1682952543
transform 1 0 304 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_222
timestamp 1682952543
transform -1 0 352 0 1 1770
box -8 -3 46 105
use FILL  FILL_2085
timestamp 1682952543
transform 1 0 352 0 1 1770
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1682952543
transform 1 0 360 0 1 1770
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1682952543
transform 1 0 368 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_384
timestamp 1682952543
transform -1 0 392 0 1 1770
box -9 -3 26 105
use FILL  FILL_2088
timestamp 1682952543
transform 1 0 392 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_223
timestamp 1682952543
transform 1 0 400 0 1 1770
box -8 -3 46 105
use FILL  FILL_2089
timestamp 1682952543
transform 1 0 440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2090
timestamp 1682952543
transform 1 0 448 0 1 1770
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1682952543
transform 1 0 456 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_246
timestamp 1682952543
transform -1 0 504 0 1 1770
box -8 -3 46 105
use FILL  FILL_2092
timestamp 1682952543
transform 1 0 504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1682952543
transform 1 0 512 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_351
timestamp 1682952543
transform 1 0 520 0 1 1770
box -8 -3 104 105
use FILL  FILL_2094
timestamp 1682952543
transform 1 0 616 0 1 1770
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1682952543
transform 1 0 624 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_388
timestamp 1682952543
transform -1 0 648 0 1 1770
box -9 -3 26 105
use FILL  FILL_2108
timestamp 1682952543
transform 1 0 648 0 1 1770
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1682952543
transform 1 0 656 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5665
timestamp 1682952543
transform 1 0 692 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_226
timestamp 1682952543
transform 1 0 664 0 1 1770
box -8 -3 46 105
use FILL  FILL_2114
timestamp 1682952543
transform 1 0 704 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5666
timestamp 1682952543
transform 1 0 724 0 1 1775
box -3 -3 3 3
use FILL  FILL_2115
timestamp 1682952543
transform 1 0 712 0 1 1770
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1682952543
transform 1 0 720 0 1 1770
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1682952543
transform 1 0 728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2118
timestamp 1682952543
transform 1 0 736 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_75
timestamp 1682952543
transform 1 0 744 0 1 1770
box -8 -3 34 105
use FILL  FILL_2119
timestamp 1682952543
transform 1 0 776 0 1 1770
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1682952543
transform 1 0 784 0 1 1770
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1682952543
transform 1 0 792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1682952543
transform 1 0 800 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_76
timestamp 1682952543
transform 1 0 808 0 1 1770
box -8 -3 34 105
use FILL  FILL_2127
timestamp 1682952543
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_2128
timestamp 1682952543
transform 1 0 848 0 1 1770
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1682952543
transform 1 0 856 0 1 1770
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1682952543
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1682952543
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1682952543
transform 1 0 880 0 1 1770
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1682952543
transform 1 0 888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2138
timestamp 1682952543
transform 1 0 896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1682952543
transform 1 0 904 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_228
timestamp 1682952543
transform -1 0 952 0 1 1770
box -8 -3 46 105
use FILL  FILL_2140
timestamp 1682952543
transform 1 0 952 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5667
timestamp 1682952543
transform 1 0 972 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_356
timestamp 1682952543
transform 1 0 960 0 1 1770
box -8 -3 104 105
use FILL  FILL_2148
timestamp 1682952543
transform 1 0 1056 0 1 1770
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1682952543
transform 1 0 1064 0 1 1770
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1682952543
transform 1 0 1072 0 1 1770
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1682952543
transform 1 0 1080 0 1 1770
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1682952543
transform 1 0 1088 0 1 1770
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1682952543
transform 1 0 1096 0 1 1770
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1682952543
transform 1 0 1104 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_78
timestamp 1682952543
transform -1 0 1144 0 1 1770
box -8 -3 34 105
use FILL  FILL_2163
timestamp 1682952543
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1682952543
transform 1 0 1152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1682952543
transform 1 0 1160 0 1 1770
box -8 -3 16 105
use FILL  FILL_2172
timestamp 1682952543
transform 1 0 1168 0 1 1770
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1682952543
transform 1 0 1176 0 1 1770
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1682952543
transform 1 0 1184 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_248
timestamp 1682952543
transform -1 0 1232 0 1 1770
box -8 -3 46 105
use FILL  FILL_2177
timestamp 1682952543
transform 1 0 1232 0 1 1770
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1682952543
transform 1 0 1240 0 1 1770
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1682952543
transform 1 0 1248 0 1 1770
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1682952543
transform 1 0 1256 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5668
timestamp 1682952543
transform 1 0 1340 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_357
timestamp 1682952543
transform 1 0 1264 0 1 1770
box -8 -3 104 105
use FILL  FILL_2181
timestamp 1682952543
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_249
timestamp 1682952543
transform -1 0 1408 0 1 1770
box -8 -3 46 105
use FILL  FILL_2182
timestamp 1682952543
transform 1 0 1408 0 1 1770
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1682952543
transform 1 0 1416 0 1 1770
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1682952543
transform 1 0 1424 0 1 1770
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1682952543
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_394
timestamp 1682952543
transform -1 0 1456 0 1 1770
box -9 -3 26 105
use FILL  FILL_2198
timestamp 1682952543
transform 1 0 1456 0 1 1770
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1682952543
transform 1 0 1464 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5669
timestamp 1682952543
transform 1 0 1484 0 1 1775
box -3 -3 3 3
use FILL  FILL_2200
timestamp 1682952543
transform 1 0 1472 0 1 1770
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1682952543
transform 1 0 1480 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_80
timestamp 1682952543
transform 1 0 1488 0 1 1770
box -5 -3 28 105
use FILL  FILL_2202
timestamp 1682952543
transform 1 0 1512 0 1 1770
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1682952543
transform 1 0 1520 0 1 1770
box -8 -3 16 105
use FILL  FILL_2204
timestamp 1682952543
transform 1 0 1528 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5670
timestamp 1682952543
transform 1 0 1564 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_251
timestamp 1682952543
transform 1 0 1536 0 1 1770
box -8 -3 46 105
use FILL  FILL_2205
timestamp 1682952543
transform 1 0 1576 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5671
timestamp 1682952543
transform 1 0 1604 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_358
timestamp 1682952543
transform -1 0 1680 0 1 1770
box -8 -3 104 105
use FILL  FILL_2206
timestamp 1682952543
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_72
timestamp 1682952543
transform 1 0 1688 0 1 1770
box -8 -3 32 105
use FILL  FILL_2207
timestamp 1682952543
transform 1 0 1712 0 1 1770
box -8 -3 16 105
use FILL  FILL_2219
timestamp 1682952543
transform 1 0 1720 0 1 1770
box -8 -3 16 105
use FILL  FILL_2220
timestamp 1682952543
transform 1 0 1728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1682952543
transform 1 0 1736 0 1 1770
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1682952543
transform 1 0 1744 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5672
timestamp 1682952543
transform 1 0 1788 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_232
timestamp 1682952543
transform 1 0 1752 0 1 1770
box -8 -3 46 105
use FILL  FILL_2224
timestamp 1682952543
transform 1 0 1792 0 1 1770
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1682952543
transform 1 0 1800 0 1 1770
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1682952543
transform 1 0 1808 0 1 1770
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1682952543
transform 1 0 1816 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_75
timestamp 1682952543
transform 1 0 1824 0 1 1770
box -8 -3 32 105
use FILL  FILL_2234
timestamp 1682952543
transform 1 0 1848 0 1 1770
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1682952543
transform 1 0 1856 0 1 1770
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1682952543
transform 1 0 1864 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_81
timestamp 1682952543
transform 1 0 1872 0 1 1770
box -5 -3 28 105
use FILL  FILL_2239
timestamp 1682952543
transform 1 0 1896 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5673
timestamp 1682952543
transform 1 0 1916 0 1 1775
box -3 -3 3 3
use FILL  FILL_2240
timestamp 1682952543
transform 1 0 1904 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_397
timestamp 1682952543
transform 1 0 1912 0 1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_360
timestamp 1682952543
transform -1 0 2024 0 1 1770
box -8 -3 104 105
use FILL  FILL_2241
timestamp 1682952543
transform 1 0 2024 0 1 1770
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1682952543
transform 1 0 2032 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_77
timestamp 1682952543
transform 1 0 2040 0 1 1770
box -8 -3 32 105
use FILL  FILL_2252
timestamp 1682952543
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1682952543
transform 1 0 2072 0 1 1770
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1682952543
transform 1 0 2080 0 1 1770
box -8 -3 16 105
use FILL  FILL_2255
timestamp 1682952543
transform 1 0 2088 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5674
timestamp 1682952543
transform 1 0 2108 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_398
timestamp 1682952543
transform 1 0 2096 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_5675
timestamp 1682952543
transform 1 0 2156 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_234
timestamp 1682952543
transform 1 0 2112 0 1 1770
box -8 -3 46 105
use FILL  FILL_2256
timestamp 1682952543
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1682952543
transform 1 0 2160 0 1 1770
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1682952543
transform 1 0 2168 0 1 1770
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1682952543
transform 1 0 2176 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_84
timestamp 1682952543
transform 1 0 2184 0 1 1770
box -8 -3 34 105
use FILL  FILL_2260
timestamp 1682952543
transform 1 0 2216 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5676
timestamp 1682952543
transform 1 0 2236 0 1 1775
box -3 -3 3 3
use FILL  FILL_2261
timestamp 1682952543
transform 1 0 2224 0 1 1770
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1682952543
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1682952543
transform 1 0 2240 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5677
timestamp 1682952543
transform 1 0 2268 0 1 1775
box -3 -3 3 3
use OAI21X1  OAI21X1_85
timestamp 1682952543
transform 1 0 2248 0 1 1770
box -8 -3 34 105
use FILL  FILL_2264
timestamp 1682952543
transform 1 0 2280 0 1 1770
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1682952543
transform 1 0 2288 0 1 1770
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1682952543
transform 1 0 2296 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_401
timestamp 1682952543
transform -1 0 2320 0 1 1770
box -9 -3 26 105
use M3_M2  M3_M2_5678
timestamp 1682952543
transform 1 0 2356 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_236
timestamp 1682952543
transform 1 0 2320 0 1 1770
box -8 -3 46 105
use FILL  FILL_2278
timestamp 1682952543
transform 1 0 2360 0 1 1770
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1682952543
transform 1 0 2368 0 1 1770
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1682952543
transform 1 0 2376 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5679
timestamp 1682952543
transform 1 0 2396 0 1 1775
box -3 -3 3 3
use FILL  FILL_2286
timestamp 1682952543
transform 1 0 2384 0 1 1770
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1682952543
transform 1 0 2392 0 1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_86
timestamp 1682952543
transform -1 0 2432 0 1 1770
box -8 -3 34 105
use FILL  FILL_2288
timestamp 1682952543
transform 1 0 2432 0 1 1770
box -8 -3 16 105
use FILL  FILL_2289
timestamp 1682952543
transform 1 0 2440 0 1 1770
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1682952543
transform 1 0 2448 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_402
timestamp 1682952543
transform 1 0 2456 0 1 1770
box -9 -3 26 105
use FILL  FILL_2291
timestamp 1682952543
transform 1 0 2472 0 1 1770
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1682952543
transform 1 0 2480 0 1 1770
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1682952543
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1682952543
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_2296
timestamp 1682952543
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1682952543
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_238
timestamp 1682952543
transform -1 0 2560 0 1 1770
box -8 -3 46 105
use FILL  FILL_2300
timestamp 1682952543
transform 1 0 2560 0 1 1770
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1682952543
transform 1 0 2568 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5680
timestamp 1682952543
transform 1 0 2588 0 1 1775
box -3 -3 3 3
use FILL  FILL_2305
timestamp 1682952543
transform 1 0 2576 0 1 1770
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1682952543
transform 1 0 2584 0 1 1770
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1682952543
transform 1 0 2592 0 1 1770
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1682952543
transform 1 0 2600 0 1 1770
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1682952543
transform 1 0 2608 0 1 1770
box -8 -3 16 105
use FILL  FILL_2313
timestamp 1682952543
transform 1 0 2616 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5681
timestamp 1682952543
transform 1 0 2660 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_240
timestamp 1682952543
transform 1 0 2624 0 1 1770
box -8 -3 46 105
use FILL  FILL_2315
timestamp 1682952543
transform 1 0 2664 0 1 1770
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1682952543
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1682952543
transform 1 0 2680 0 1 1770
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1682952543
transform 1 0 2688 0 1 1770
box -8 -3 16 105
use FILL  FILL_2324
timestamp 1682952543
transform 1 0 2696 0 1 1770
box -8 -3 16 105
use FILL  FILL_2326
timestamp 1682952543
transform 1 0 2704 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_405
timestamp 1682952543
transform 1 0 2712 0 1 1770
box -9 -3 26 105
use FILL  FILL_2327
timestamp 1682952543
transform 1 0 2728 0 1 1770
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1682952543
transform 1 0 2736 0 1 1770
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1682952543
transform 1 0 2744 0 1 1770
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1682952543
transform 1 0 2752 0 1 1770
box -8 -3 16 105
use FILL  FILL_2334
timestamp 1682952543
transform 1 0 2760 0 1 1770
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1682952543
transform 1 0 2768 0 1 1770
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1682952543
transform 1 0 2776 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_48
timestamp 1682952543
transform 1 0 2784 0 1 1770
box -8 -3 40 105
use FILL  FILL_2337
timestamp 1682952543
transform 1 0 2816 0 1 1770
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1682952543
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_2339
timestamp 1682952543
transform 1 0 2832 0 1 1770
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1682952543
transform 1 0 2840 0 1 1770
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1682952543
transform 1 0 2848 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_49
timestamp 1682952543
transform -1 0 2888 0 1 1770
box -8 -3 40 105
use FILL  FILL_2342
timestamp 1682952543
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1682952543
transform 1 0 2896 0 1 1770
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1682952543
transform 1 0 2904 0 1 1770
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1682952543
transform 1 0 2912 0 1 1770
box -8 -3 16 105
use FILL  FILL_2358
timestamp 1682952543
transform 1 0 2920 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_407
timestamp 1682952543
transform -1 0 2944 0 1 1770
box -9 -3 26 105
use FILL  FILL_2359
timestamp 1682952543
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5682
timestamp 1682952543
transform 1 0 3004 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_363
timestamp 1682952543
transform -1 0 3048 0 1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_364
timestamp 1682952543
transform 1 0 3048 0 1 1770
box -8 -3 104 105
use FILL  FILL_2360
timestamp 1682952543
transform 1 0 3144 0 1 1770
box -8 -3 16 105
use FILL  FILL_2377
timestamp 1682952543
transform 1 0 3152 0 1 1770
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1682952543
transform 1 0 3160 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_365
timestamp 1682952543
transform -1 0 3264 0 1 1770
box -8 -3 104 105
use FILL  FILL_2380
timestamp 1682952543
transform 1 0 3264 0 1 1770
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1682952543
transform 1 0 3272 0 1 1770
box -8 -3 16 105
use FILL  FILL_2382
timestamp 1682952543
transform 1 0 3280 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_52
timestamp 1682952543
transform -1 0 3320 0 1 1770
box -8 -3 40 105
use FILL  FILL_2383
timestamp 1682952543
transform 1 0 3320 0 1 1770
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1682952543
transform 1 0 3328 0 1 1770
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1682952543
transform 1 0 3336 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_255
timestamp 1682952543
transform 1 0 3344 0 1 1770
box -8 -3 46 105
use FILL  FILL_2399
timestamp 1682952543
transform 1 0 3384 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5683
timestamp 1682952543
transform 1 0 3420 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5684
timestamp 1682952543
transform 1 0 3468 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_366
timestamp 1682952543
transform 1 0 3392 0 1 1770
box -8 -3 104 105
use M3_M2  M3_M2_5685
timestamp 1682952543
transform 1 0 3524 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_256
timestamp 1682952543
transform 1 0 3488 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_410
timestamp 1682952543
transform -1 0 3544 0 1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_53
timestamp 1682952543
transform -1 0 3576 0 1 1770
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_367
timestamp 1682952543
transform -1 0 3672 0 1 1770
box -8 -3 104 105
use NAND3X1  NAND3X1_54
timestamp 1682952543
transform -1 0 3704 0 1 1770
box -8 -3 40 105
use NAND3X1  NAND3X1_55
timestamp 1682952543
transform -1 0 3736 0 1 1770
box -8 -3 40 105
use BUFX2  BUFX2_84
timestamp 1682952543
transform 1 0 3736 0 1 1770
box -5 -3 28 105
use FILL  FILL_2400
timestamp 1682952543
transform 1 0 3760 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5686
timestamp 1682952543
transform 1 0 3780 0 1 1775
box -3 -3 3 3
use FILL  FILL_2401
timestamp 1682952543
transform 1 0 3768 0 1 1770
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1682952543
transform 1 0 3776 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5687
timestamp 1682952543
transform 1 0 3828 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_242
timestamp 1682952543
transform -1 0 3824 0 1 1770
box -8 -3 46 105
use FILL  FILL_2409
timestamp 1682952543
transform 1 0 3824 0 1 1770
box -8 -3 16 105
use FILL  FILL_2411
timestamp 1682952543
transform 1 0 3832 0 1 1770
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1682952543
transform 1 0 3840 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5688
timestamp 1682952543
transform 1 0 3884 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_258
timestamp 1682952543
transform 1 0 3848 0 1 1770
box -8 -3 46 105
use FILL  FILL_2415
timestamp 1682952543
transform 1 0 3888 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_243
timestamp 1682952543
transform -1 0 3936 0 1 1770
box -8 -3 46 105
use INVX2  INVX2_413
timestamp 1682952543
transform -1 0 3952 0 1 1770
box -9 -3 26 105
use FILL  FILL_2416
timestamp 1682952543
transform 1 0 3952 0 1 1770
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1682952543
transform 1 0 3960 0 1 1770
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1682952543
transform 1 0 3968 0 1 1770
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1682952543
transform 1 0 3976 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_260
timestamp 1682952543
transform 1 0 3984 0 1 1770
box -8 -3 46 105
use FILL  FILL_2427
timestamp 1682952543
transform 1 0 4024 0 1 1770
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1682952543
transform 1 0 4032 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_371
timestamp 1682952543
transform 1 0 4040 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_415
timestamp 1682952543
transform -1 0 4152 0 1 1770
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_47
timestamp 1682952543
transform 1 0 4177 0 1 1770
box -10 -3 10 3
use M2_M1  M2_M1_5750
timestamp 1682952543
transform 1 0 92 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1682952543
transform 1 0 140 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1682952543
transform 1 0 172 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5811
timestamp 1682952543
transform 1 0 140 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5858
timestamp 1682952543
transform 1 0 172 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_5844
timestamp 1682952543
transform 1 0 188 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5812
timestamp 1682952543
transform 1 0 188 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1682952543
transform 1 0 252 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_5751
timestamp 1682952543
transform 1 0 236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1682952543
transform 1 0 244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5753
timestamp 1682952543
transform 1 0 260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1682952543
transform 1 0 228 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5800
timestamp 1682952543
transform 1 0 244 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5690
timestamp 1682952543
transform 1 0 316 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1682952543
transform 1 0 284 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5709
timestamp 1682952543
transform 1 0 308 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5743
timestamp 1682952543
transform 1 0 364 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5754
timestamp 1682952543
transform 1 0 284 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5744
timestamp 1682952543
transform 1 0 412 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5755
timestamp 1682952543
transform 1 0 388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5756
timestamp 1682952543
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1682952543
transform 1 0 412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1682952543
transform 1 0 428 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5846
timestamp 1682952543
transform 1 0 252 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1682952543
transform 1 0 268 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1682952543
transform 1 0 332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1682952543
transform 1 0 364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5850
timestamp 1682952543
transform 1 0 372 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1682952543
transform 1 0 388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5852
timestamp 1682952543
transform 1 0 404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1682952543
transform 1 0 420 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5859
timestamp 1682952543
transform 1 0 244 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5813
timestamp 1682952543
transform 1 0 332 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5814
timestamp 1682952543
transform 1 0 372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1682952543
transform 1 0 316 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5891
timestamp 1682952543
transform 1 0 268 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1682952543
transform 1 0 388 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5691
timestamp 1682952543
transform 1 0 508 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1682952543
transform 1 0 452 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1682952543
transform 1 0 540 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1682952543
transform 1 0 492 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1682952543
transform 1 0 532 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5759
timestamp 1682952543
transform 1 0 452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1682952543
transform 1 0 436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5855
timestamp 1682952543
transform 1 0 476 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1682952543
transform 1 0 532 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5815
timestamp 1682952543
transform 1 0 436 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5816
timestamp 1682952543
transform 1 0 476 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1682952543
transform 1 0 428 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5872
timestamp 1682952543
transform 1 0 380 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5873
timestamp 1682952543
transform 1 0 396 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5874
timestamp 1682952543
transform 1 0 428 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1682952543
transform 1 0 476 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5892
timestamp 1682952543
transform 1 0 444 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_5760
timestamp 1682952543
transform 1 0 588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5761
timestamp 1682952543
transform 1 0 604 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1682952543
transform 1 0 580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1682952543
transform 1 0 596 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5801
timestamp 1682952543
transform 1 0 604 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1682952543
transform 1 0 644 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1682952543
transform 1 0 660 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5747
timestamp 1682952543
transform 1 0 668 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1682952543
transform 1 0 748 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5762
timestamp 1682952543
transform 1 0 668 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1682952543
transform 1 0 708 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5860
timestamp 1682952543
transform 1 0 748 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5861
timestamp 1682952543
transform 1 0 756 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5817
timestamp 1682952543
transform 1 0 708 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5864
timestamp 1682952543
transform 1 0 692 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5893
timestamp 1682952543
transform 1 0 724 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5818
timestamp 1682952543
transform 1 0 756 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1682952543
transform 1 0 772 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_5763
timestamp 1682952543
transform 1 0 804 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5819
timestamp 1682952543
transform 1 0 804 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5895
timestamp 1682952543
transform 1 0 804 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5712
timestamp 1682952543
transform 1 0 820 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1682952543
transform 1 0 860 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5749
timestamp 1682952543
transform 1 0 852 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5764
timestamp 1682952543
transform 1 0 820 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5784
timestamp 1682952543
transform 1 0 836 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5765
timestamp 1682952543
transform 1 0 852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5862
timestamp 1682952543
transform 1 0 820 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5863
timestamp 1682952543
transform 1 0 836 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1682952543
transform 1 0 852 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5820
timestamp 1682952543
transform 1 0 836 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1682952543
transform 1 0 852 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1682952543
transform 1 0 868 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1682952543
transform 1 0 868 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5695
timestamp 1682952543
transform 1 0 884 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1682952543
transform 1 0 900 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1682952543
transform 1 0 892 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5785
timestamp 1682952543
transform 1 0 884 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5766
timestamp 1682952543
transform 1 0 900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5865
timestamp 1682952543
transform 1 0 884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1682952543
transform 1 0 908 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5866
timestamp 1682952543
transform 1 0 924 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_5767
timestamp 1682952543
transform 1 0 972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1682952543
transform 1 0 988 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5786
timestamp 1682952543
transform 1 0 996 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5867
timestamp 1682952543
transform 1 0 980 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5802
timestamp 1682952543
transform 1 0 988 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_5868
timestamp 1682952543
transform 1 0 996 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1682952543
transform 1 0 956 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5821
timestamp 1682952543
transform 1 0 964 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5875
timestamp 1682952543
transform 1 0 964 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5876
timestamp 1682952543
transform 1 0 1004 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1682952543
transform 1 0 1020 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5869
timestamp 1682952543
transform 1 0 1028 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5769
timestamp 1682952543
transform 1 0 1068 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5870
timestamp 1682952543
transform 1 0 1084 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1682952543
transform 1 0 1100 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5867
timestamp 1682952543
transform 1 0 1084 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1682952543
transform 1 0 1116 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5770
timestamp 1682952543
transform 1 0 1140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5872
timestamp 1682952543
transform 1 0 1140 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5877
timestamp 1682952543
transform 1 0 1156 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_5771
timestamp 1682952543
transform 1 0 1172 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5772
timestamp 1682952543
transform 1 0 1180 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5822
timestamp 1682952543
transform 1 0 1180 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1682952543
transform 1 0 1212 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5717
timestamp 1682952543
transform 1 0 1236 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1682952543
transform 1 0 1204 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5788
timestamp 1682952543
transform 1 0 1196 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5878
timestamp 1682952543
transform 1 0 1196 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5753
timestamp 1682952543
transform 1 0 1260 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5773
timestamp 1682952543
transform 1 0 1236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1682952543
transform 1 0 1244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5873
timestamp 1682952543
transform 1 0 1228 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5789
timestamp 1682952543
transform 1 0 1268 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5874
timestamp 1682952543
transform 1 0 1260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5951
timestamp 1682952543
transform 1 0 1212 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5823
timestamp 1682952543
transform 1 0 1236 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5952
timestamp 1682952543
transform 1 0 1244 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5824
timestamp 1682952543
transform 1 0 1260 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5879
timestamp 1682952543
transform 1 0 1212 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5880
timestamp 1682952543
transform 1 0 1244 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5881
timestamp 1682952543
transform 1 0 1268 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5718
timestamp 1682952543
transform 1 0 1284 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5754
timestamp 1682952543
transform 1 0 1300 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5755
timestamp 1682952543
transform 1 0 1348 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5775
timestamp 1682952543
transform 1 0 1292 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5776
timestamp 1682952543
transform 1 0 1300 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5777
timestamp 1682952543
transform 1 0 1316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5778
timestamp 1682952543
transform 1 0 1332 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5719
timestamp 1682952543
transform 1 0 1380 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5779
timestamp 1682952543
transform 1 0 1356 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5780
timestamp 1682952543
transform 1 0 1364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5875
timestamp 1682952543
transform 1 0 1308 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5876
timestamp 1682952543
transform 1 0 1324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1682952543
transform 1 0 1332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1682952543
transform 1 0 1348 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5825
timestamp 1682952543
transform 1 0 1308 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5826
timestamp 1682952543
transform 1 0 1332 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5882
timestamp 1682952543
transform 1 0 1308 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5883
timestamp 1682952543
transform 1 0 1324 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5884
timestamp 1682952543
transform 1 0 1348 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5790
timestamp 1682952543
transform 1 0 1372 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5756
timestamp 1682952543
transform 1 0 1396 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1682952543
transform 1 0 1388 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5879
timestamp 1682952543
transform 1 0 1380 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5885
timestamp 1682952543
transform 1 0 1412 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_5781
timestamp 1682952543
transform 1 0 1428 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5757
timestamp 1682952543
transform 1 0 1468 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1682952543
transform 1 0 1492 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5782
timestamp 1682952543
transform 1 0 1444 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5792
timestamp 1682952543
transform 1 0 1468 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5880
timestamp 1682952543
transform 1 0 1468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1682952543
transform 1 0 1524 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1682952543
transform 1 0 1532 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5827
timestamp 1682952543
transform 1 0 1492 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1682952543
transform 1 0 1524 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1682952543
transform 1 0 1556 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5783
timestamp 1682952543
transform 1 0 1548 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1682952543
transform 1 0 1564 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1682952543
transform 1 0 1580 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1682952543
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1682952543
transform 1 0 1556 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1682952543
transform 1 0 1572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1682952543
transform 1 0 1588 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5829
timestamp 1682952543
transform 1 0 1580 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5886
timestamp 1682952543
transform 1 0 1604 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5830
timestamp 1682952543
transform 1 0 1596 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5787
timestamp 1682952543
transform 1 0 1644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1682952543
transform 1 0 1636 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5831
timestamp 1682952543
transform 1 0 1644 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5888
timestamp 1682952543
transform 1 0 1660 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5696
timestamp 1682952543
transform 1 0 1724 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_5740
timestamp 1682952543
transform 1 0 1716 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5788
timestamp 1682952543
transform 1 0 1708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5953
timestamp 1682952543
transform 1 0 1716 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5721
timestamp 1682952543
transform 1 0 1740 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5741
timestamp 1682952543
transform 1 0 1740 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_5722
timestamp 1682952543
transform 1 0 1756 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1682952543
transform 1 0 1780 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5789
timestamp 1682952543
transform 1 0 1780 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1682952543
transform 1 0 1788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5791
timestamp 1682952543
transform 1 0 1796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1682952543
transform 1 0 1772 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1682952543
transform 1 0 1796 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1682952543
transform 1 0 1804 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5886
timestamp 1682952543
transform 1 0 1812 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5723
timestamp 1682952543
transform 1 0 1860 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5792
timestamp 1682952543
transform 1 0 1852 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5832
timestamp 1682952543
transform 1 0 1836 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5793
timestamp 1682952543
transform 1 0 1860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1682952543
transform 1 0 1868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5954
timestamp 1682952543
transform 1 0 1868 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5833
timestamp 1682952543
transform 1 0 1876 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5964
timestamp 1682952543
transform 1 0 1876 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5724
timestamp 1682952543
transform 1 0 1908 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5893
timestamp 1682952543
transform 1 0 1900 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1682952543
transform 1 0 1916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1682952543
transform 1 0 1932 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1682952543
transform 1 0 1932 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5697
timestamp 1682952543
transform 1 0 1948 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_5896
timestamp 1682952543
transform 1 0 1964 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5834
timestamp 1682952543
transform 1 0 1956 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5887
timestamp 1682952543
transform 1 0 1972 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_5743
timestamp 1682952543
transform 1 0 1988 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1682952543
transform 1 0 1988 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5760
timestamp 1682952543
transform 1 0 2004 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5794
timestamp 1682952543
transform 1 0 2004 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5835
timestamp 1682952543
transform 1 0 2012 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5888
timestamp 1682952543
transform 1 0 2020 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_5795
timestamp 1682952543
transform 1 0 2044 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5889
timestamp 1682952543
transform 1 0 2044 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1682952543
transform 1 0 2068 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5761
timestamp 1682952543
transform 1 0 2060 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5796
timestamp 1682952543
transform 1 0 2068 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5897
timestamp 1682952543
transform 1 0 2060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5898
timestamp 1682952543
transform 1 0 2068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1682952543
transform 1 0 2084 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5836
timestamp 1682952543
transform 1 0 2084 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5900
timestamp 1682952543
transform 1 0 2108 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5726
timestamp 1682952543
transform 1 0 2116 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5744
timestamp 1682952543
transform 1 0 2116 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_5762
timestamp 1682952543
transform 1 0 2124 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5797
timestamp 1682952543
transform 1 0 2124 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5727
timestamp 1682952543
transform 1 0 2132 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5745
timestamp 1682952543
transform 1 0 2132 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1682952543
transform 1 0 2132 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5837
timestamp 1682952543
transform 1 0 2132 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5728
timestamp 1682952543
transform 1 0 2164 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5763
timestamp 1682952543
transform 1 0 2164 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5764
timestamp 1682952543
transform 1 0 2180 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5799
timestamp 1682952543
transform 1 0 2244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1682952543
transform 1 0 2156 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5902
timestamp 1682952543
transform 1 0 2164 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5903
timestamp 1682952543
transform 1 0 2196 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5838
timestamp 1682952543
transform 1 0 2156 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5839
timestamp 1682952543
transform 1 0 2196 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5904
timestamp 1682952543
transform 1 0 2260 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5729
timestamp 1682952543
transform 1 0 2292 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5765
timestamp 1682952543
transform 1 0 2300 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5730
timestamp 1682952543
transform 1 0 2316 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5800
timestamp 1682952543
transform 1 0 2316 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5801
timestamp 1682952543
transform 1 0 2324 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1682952543
transform 1 0 2340 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1682952543
transform 1 0 2348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5905
timestamp 1682952543
transform 1 0 2308 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5840
timestamp 1682952543
transform 1 0 2300 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5906
timestamp 1682952543
transform 1 0 2332 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5841
timestamp 1682952543
transform 1 0 2332 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5907
timestamp 1682952543
transform 1 0 2364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1682952543
transform 1 0 2364 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5731
timestamp 1682952543
transform 1 0 2452 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5804
timestamp 1682952543
transform 1 0 2388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5908
timestamp 1682952543
transform 1 0 2436 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5909
timestamp 1682952543
transform 1 0 2468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5910
timestamp 1682952543
transform 1 0 2476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5842
timestamp 1682952543
transform 1 0 2436 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5843
timestamp 1682952543
transform 1 0 2476 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1682952543
transform 1 0 2500 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5911
timestamp 1682952543
transform 1 0 2500 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5732
timestamp 1682952543
transform 1 0 2524 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5805
timestamp 1682952543
transform 1 0 2516 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5844
timestamp 1682952543
transform 1 0 2516 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5806
timestamp 1682952543
transform 1 0 2524 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1682952543
transform 1 0 2556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5912
timestamp 1682952543
transform 1 0 2548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1682952543
transform 1 0 2564 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5845
timestamp 1682952543
transform 1 0 2548 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1682952543
transform 1 0 2596 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5767
timestamp 1682952543
transform 1 0 2588 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5914
timestamp 1682952543
transform 1 0 2588 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5734
timestamp 1682952543
transform 1 0 2660 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5808
timestamp 1682952543
transform 1 0 2644 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5915
timestamp 1682952543
transform 1 0 2636 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5957
timestamp 1682952543
transform 1 0 2668 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5698
timestamp 1682952543
transform 1 0 2708 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_5809
timestamp 1682952543
transform 1 0 2700 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5810
timestamp 1682952543
transform 1 0 2708 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1682952543
transform 1 0 2700 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5768
timestamp 1682952543
transform 1 0 2732 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5958
timestamp 1682952543
transform 1 0 2748 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5868
timestamp 1682952543
transform 1 0 2756 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_5965
timestamp 1682952543
transform 1 0 2764 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5769
timestamp 1682952543
transform 1 0 2796 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5917
timestamp 1682952543
transform 1 0 2788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5959
timestamp 1682952543
transform 1 0 2796 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1682952543
transform 1 0 2804 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_5918
timestamp 1682952543
transform 1 0 2836 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5803
timestamp 1682952543
transform 1 0 2844 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_5960
timestamp 1682952543
transform 1 0 2844 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_5967
timestamp 1682952543
transform 1 0 2836 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5896
timestamp 1682952543
transform 1 0 2836 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5793
timestamp 1682952543
transform 1 0 2868 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1682952543
transform 1 0 2876 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_5811
timestamp 1682952543
transform 1 0 2916 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1682952543
transform 1 0 2932 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1682952543
transform 1 0 2948 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1682952543
transform 1 0 2924 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5920
timestamp 1682952543
transform 1 0 2964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1682952543
transform 1 0 2996 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5770
timestamp 1682952543
transform 1 0 3012 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5814
timestamp 1682952543
transform 1 0 3028 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1682952543
transform 1 0 3020 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5923
timestamp 1682952543
transform 1 0 3036 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5846
timestamp 1682952543
transform 1 0 3020 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5924
timestamp 1682952543
transform 1 0 3052 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5805
timestamp 1682952543
transform 1 0 3060 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5847
timestamp 1682952543
transform 1 0 3052 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1682952543
transform 1 0 3076 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5815
timestamp 1682952543
transform 1 0 3076 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5772
timestamp 1682952543
transform 1 0 3124 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5746
timestamp 1682952543
transform 1 0 3132 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1682952543
transform 1 0 3092 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5817
timestamp 1682952543
transform 1 0 3108 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5818
timestamp 1682952543
transform 1 0 3124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1682952543
transform 1 0 3116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5926
timestamp 1682952543
transform 1 0 3132 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5848
timestamp 1682952543
transform 1 0 3124 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1682952543
transform 1 0 3140 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5819
timestamp 1682952543
transform 1 0 3156 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5735
timestamp 1682952543
transform 1 0 3164 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5747
timestamp 1682952543
transform 1 0 3164 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_5736
timestamp 1682952543
transform 1 0 3196 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5820
timestamp 1682952543
transform 1 0 3196 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5773
timestamp 1682952543
transform 1 0 3220 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5821
timestamp 1682952543
transform 1 0 3244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1682952543
transform 1 0 3236 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1682952543
transform 1 0 3260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1682952543
transform 1 0 3276 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5699
timestamp 1682952543
transform 1 0 3324 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_5823
timestamp 1682952543
transform 1 0 3308 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5794
timestamp 1682952543
transform 1 0 3316 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5774
timestamp 1682952543
transform 1 0 3332 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5795
timestamp 1682952543
transform 1 0 3332 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5929
timestamp 1682952543
transform 1 0 3324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1682952543
transform 1 0 3332 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5737
timestamp 1682952543
transform 1 0 3348 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1682952543
transform 1 0 3372 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1682952543
transform 1 0 3404 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5776
timestamp 1682952543
transform 1 0 3404 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5824
timestamp 1682952543
transform 1 0 3372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5825
timestamp 1682952543
transform 1 0 3396 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5796
timestamp 1682952543
transform 1 0 3412 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5931
timestamp 1682952543
transform 1 0 3380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5932
timestamp 1682952543
transform 1 0 3396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5933
timestamp 1682952543
transform 1 0 3404 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5850
timestamp 1682952543
transform 1 0 3396 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5700
timestamp 1682952543
transform 1 0 3436 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5777
timestamp 1682952543
transform 1 0 3436 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5826
timestamp 1682952543
transform 1 0 3436 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5797
timestamp 1682952543
transform 1 0 3444 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5961
timestamp 1682952543
transform 1 0 3436 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5701
timestamp 1682952543
transform 1 0 3500 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5702
timestamp 1682952543
transform 1 0 3540 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1682952543
transform 1 0 3564 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1682952543
transform 1 0 3476 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5740
timestamp 1682952543
transform 1 0 3516 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_5934
timestamp 1682952543
transform 1 0 3460 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5851
timestamp 1682952543
transform 1 0 3452 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5778
timestamp 1682952543
transform 1 0 3484 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1682952543
transform 1 0 3500 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5827
timestamp 1682952543
transform 1 0 3484 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5806
timestamp 1682952543
transform 1 0 3484 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5780
timestamp 1682952543
transform 1 0 3580 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5781
timestamp 1682952543
transform 1 0 3596 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5828
timestamp 1682952543
transform 1 0 3580 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5704
timestamp 1682952543
transform 1 0 3732 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5705
timestamp 1682952543
transform 1 0 3756 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_5829
timestamp 1682952543
transform 1 0 3676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5935
timestamp 1682952543
transform 1 0 3508 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1682952543
transform 1 0 3564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1682952543
transform 1 0 3604 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5938
timestamp 1682952543
transform 1 0 3660 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5962
timestamp 1682952543
transform 1 0 3468 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5869
timestamp 1682952543
transform 1 0 3444 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_5968
timestamp 1682952543
transform 1 0 3452 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5852
timestamp 1682952543
transform 1 0 3532 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5853
timestamp 1682952543
transform 1 0 3564 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5870
timestamp 1682952543
transform 1 0 3484 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5871
timestamp 1682952543
transform 1 0 3524 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5890
timestamp 1682952543
transform 1 0 3620 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5807
timestamp 1682952543
transform 1 0 3676 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_5939
timestamp 1682952543
transform 1 0 3724 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5854
timestamp 1682952543
transform 1 0 3724 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5830
timestamp 1682952543
transform 1 0 3780 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5808
timestamp 1682952543
transform 1 0 3772 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_5940
timestamp 1682952543
transform 1 0 3780 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1682952543
transform 1 0 3804 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1682952543
transform 1 0 3820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5941
timestamp 1682952543
transform 1 0 3796 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5855
timestamp 1682952543
transform 1 0 3804 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5748
timestamp 1682952543
transform 1 0 3844 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1682952543
transform 1 0 3844 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5809
timestamp 1682952543
transform 1 0 3844 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_5834
timestamp 1682952543
transform 1 0 3876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5835
timestamp 1682952543
transform 1 0 3892 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5942
timestamp 1682952543
transform 1 0 3860 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5943
timestamp 1682952543
transform 1 0 3884 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1682952543
transform 1 0 3924 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5798
timestamp 1682952543
transform 1 0 3932 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5944
timestamp 1682952543
transform 1 0 3932 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5856
timestamp 1682952543
transform 1 0 3932 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5749
timestamp 1682952543
transform 1 0 3948 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_5837
timestamp 1682952543
transform 1 0 3948 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5810
timestamp 1682952543
transform 1 0 3948 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_5963
timestamp 1682952543
transform 1 0 3948 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5782
timestamp 1682952543
transform 1 0 3980 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5838
timestamp 1682952543
transform 1 0 3980 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1682952543
transform 1 0 3972 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5946
timestamp 1682952543
transform 1 0 3988 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5857
timestamp 1682952543
transform 1 0 3988 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_5839
timestamp 1682952543
transform 1 0 4020 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5706
timestamp 1682952543
transform 1 0 4036 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5707
timestamp 1682952543
transform 1 0 4084 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1682952543
transform 1 0 4036 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1682952543
transform 1 0 4052 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5783
timestamp 1682952543
transform 1 0 4060 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_5840
timestamp 1682952543
transform 1 0 4036 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5799
timestamp 1682952543
transform 1 0 4116 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_5841
timestamp 1682952543
transform 1 0 4132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_5947
timestamp 1682952543
transform 1 0 4060 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1682952543
transform 1 0 4116 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_5949
timestamp 1682952543
transform 1 0 4124 0 1 1725
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_48
timestamp 1682952543
transform 1 0 24 0 1 1670
box -10 -3 10 3
use FILL  FILL_2095
timestamp 1682952543
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_352
timestamp 1682952543
transform 1 0 80 0 -1 1770
box -8 -3 104 105
use FILL  FILL_2096
timestamp 1682952543
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1682952543
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1682952543
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1682952543
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1682952543
transform 1 0 208 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_385
timestamp 1682952543
transform -1 0 232 0 -1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_224
timestamp 1682952543
transform -1 0 272 0 -1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_353
timestamp 1682952543
transform 1 0 272 0 -1 1770
box -8 -3 104 105
use M3_M2  M3_M2_5897
timestamp 1682952543
transform 1 0 388 0 1 1675
box -3 -3 3 3
use INVX2  INVX2_386
timestamp 1682952543
transform -1 0 384 0 -1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_225
timestamp 1682952543
transform 1 0 384 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_387
timestamp 1682952543
transform 1 0 424 0 -1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_354
timestamp 1682952543
transform 1 0 440 0 -1 1770
box -8 -3 104 105
use FILL  FILL_2101
timestamp 1682952543
transform 1 0 536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1682952543
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2103
timestamp 1682952543
transform 1 0 552 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1682952543
transform 1 0 560 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_247
timestamp 1682952543
transform 1 0 568 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2105
timestamp 1682952543
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1682952543
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2109
timestamp 1682952543
transform 1 0 624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1682952543
transform 1 0 632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1682952543
transform 1 0 640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1682952543
transform 1 0 648 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_355
timestamp 1682952543
transform 1 0 656 0 -1 1770
box -8 -3 104 105
use FILL  FILL_2120
timestamp 1682952543
transform 1 0 752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1682952543
transform 1 0 760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1682952543
transform 1 0 768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1682952543
transform 1 0 776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2130
timestamp 1682952543
transform 1 0 784 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_389
timestamp 1682952543
transform -1 0 808 0 -1 1770
box -9 -3 26 105
use M3_M2  M3_M2_5898
timestamp 1682952543
transform 1 0 820 0 1 1675
box -3 -3 3 3
use FILL  FILL_2131
timestamp 1682952543
transform 1 0 808 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_227
timestamp 1682952543
transform 1 0 816 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2132
timestamp 1682952543
transform 1 0 856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2134
timestamp 1682952543
transform 1 0 864 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5899
timestamp 1682952543
transform 1 0 884 0 1 1675
box -3 -3 3 3
use OAI21X1  OAI21X1_77
timestamp 1682952543
transform 1 0 872 0 -1 1770
box -8 -3 34 105
use FILL  FILL_2141
timestamp 1682952543
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1682952543
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1682952543
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2144
timestamp 1682952543
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1682952543
transform 1 0 936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1682952543
transform 1 0 944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1682952543
transform 1 0 952 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_229
timestamp 1682952543
transform 1 0 960 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2149
timestamp 1682952543
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1682952543
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1682952543
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1682952543
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1682952543
transform 1 0 1032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2154
timestamp 1682952543
transform 1 0 1040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1682952543
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1682952543
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_230
timestamp 1682952543
transform 1 0 1064 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2164
timestamp 1682952543
transform 1 0 1104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1682952543
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1682952543
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1682952543
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1682952543
transform 1 0 1136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1682952543
transform 1 0 1144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2174
timestamp 1682952543
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_390
timestamp 1682952543
transform -1 0 1176 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2175
timestamp 1682952543
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1682952543
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1682952543
transform 1 0 1192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1682952543
transform 1 0 1200 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_79
timestamp 1682952543
transform -1 0 1240 0 -1 1770
box -8 -3 34 105
use OAI21X1  OAI21X1_80
timestamp 1682952543
transform -1 0 1272 0 -1 1770
box -8 -3 34 105
use FILL  FILL_2187
timestamp 1682952543
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1682952543
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1682952543
transform 1 0 1288 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5900
timestamp 1682952543
transform 1 0 1316 0 1 1675
box -3 -3 3 3
use OAI22X1  OAI22X1_250
timestamp 1682952543
transform -1 0 1336 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_391
timestamp 1682952543
transform -1 0 1352 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2190
timestamp 1682952543
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_392
timestamp 1682952543
transform 1 0 1360 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2191
timestamp 1682952543
transform 1 0 1376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1682952543
transform 1 0 1384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1682952543
transform 1 0 1392 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_393
timestamp 1682952543
transform -1 0 1416 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2194
timestamp 1682952543
transform 1 0 1416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2196
timestamp 1682952543
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_359
timestamp 1682952543
transform 1 0 1432 0 -1 1770
box -8 -3 104 105
use FILL  FILL_2208
timestamp 1682952543
transform 1 0 1528 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_395
timestamp 1682952543
transform -1 0 1552 0 -1 1770
box -9 -3 26 105
use AOI22X1  AOI22X1_231
timestamp 1682952543
transform 1 0 1552 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2209
timestamp 1682952543
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1682952543
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1682952543
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2212
timestamp 1682952543
transform 1 0 1616 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_396
timestamp 1682952543
transform 1 0 1624 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2213
timestamp 1682952543
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1682952543
transform 1 0 1648 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2215
timestamp 1682952543
transform 1 0 1656 0 -1 1770
box -8 -3 16 105
use OAI21X1  OAI21X1_81
timestamp 1682952543
transform 1 0 1664 0 -1 1770
box -8 -3 34 105
use FILL  FILL_2216
timestamp 1682952543
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1682952543
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1682952543
transform 1 0 1712 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_73
timestamp 1682952543
transform 1 0 1720 0 -1 1770
box -8 -3 32 105
use FILL  FILL_2223
timestamp 1682952543
transform 1 0 1744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1682952543
transform 1 0 1752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1682952543
transform 1 0 1760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2228
timestamp 1682952543
transform 1 0 1768 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5901
timestamp 1682952543
transform 1 0 1804 0 1 1675
box -3 -3 3 3
use NOR2X1  NOR2X1_74
timestamp 1682952543
transform 1 0 1776 0 -1 1770
box -8 -3 32 105
use FILL  FILL_2229
timestamp 1682952543
transform 1 0 1800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1682952543
transform 1 0 1808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1682952543
transform 1 0 1816 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5902
timestamp 1682952543
transform 1 0 1852 0 1 1675
box -3 -3 3 3
use OAI21X1  OAI21X1_82
timestamp 1682952543
transform 1 0 1824 0 -1 1770
box -8 -3 34 105
use FILL  FILL_2236
timestamp 1682952543
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1682952543
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1682952543
transform 1 0 1872 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_233
timestamp 1682952543
transform 1 0 1880 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2244
timestamp 1682952543
transform 1 0 1920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1682952543
transform 1 0 1928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1682952543
transform 1 0 1936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1682952543
transform 1 0 1944 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5903
timestamp 1682952543
transform 1 0 1964 0 1 1675
box -3 -3 3 3
use OAI21X1  OAI21X1_83
timestamp 1682952543
transform 1 0 1952 0 -1 1770
box -8 -3 34 105
use M3_M2  M3_M2_5904
timestamp 1682952543
transform 1 0 1996 0 1 1675
box -3 -3 3 3
use FILL  FILL_2248
timestamp 1682952543
transform 1 0 1984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1682952543
transform 1 0 1992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1682952543
transform 1 0 2000 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_76
timestamp 1682952543
transform 1 0 2008 0 -1 1770
box -8 -3 32 105
use FILL  FILL_2251
timestamp 1682952543
transform 1 0 2032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1682952543
transform 1 0 2040 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5905
timestamp 1682952543
transform 1 0 2060 0 1 1675
box -3 -3 3 3
use FILL  FILL_2266
timestamp 1682952543
transform 1 0 2048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1682952543
transform 1 0 2056 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5906
timestamp 1682952543
transform 1 0 2084 0 1 1675
box -3 -3 3 3
use AOI22X1  AOI22X1_235
timestamp 1682952543
transform 1 0 2064 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2268
timestamp 1682952543
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1682952543
transform 1 0 2112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2270
timestamp 1682952543
transform 1 0 2120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1682952543
transform 1 0 2128 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_399
timestamp 1682952543
transform 1 0 2136 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2272
timestamp 1682952543
transform 1 0 2152 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_361
timestamp 1682952543
transform -1 0 2256 0 -1 1770
box -8 -3 104 105
use FILL  FILL_2273
timestamp 1682952543
transform 1 0 2256 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_400
timestamp 1682952543
transform -1 0 2280 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2274
timestamp 1682952543
transform 1 0 2280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1682952543
transform 1 0 2288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1682952543
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1682952543
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_237
timestamp 1682952543
transform 1 0 2312 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2281
timestamp 1682952543
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1682952543
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1682952543
transform 1 0 2368 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_362
timestamp 1682952543
transform 1 0 2376 0 -1 1770
box -8 -3 104 105
use FILL  FILL_2292
timestamp 1682952543
transform 1 0 2472 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1682952543
transform 1 0 2480 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_403
timestamp 1682952543
transform -1 0 2504 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2298
timestamp 1682952543
transform 1 0 2504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1682952543
transform 1 0 2512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1682952543
transform 1 0 2520 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_239
timestamp 1682952543
transform -1 0 2568 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2304
timestamp 1682952543
transform 1 0 2568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1682952543
transform 1 0 2576 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5907
timestamp 1682952543
transform 1 0 2604 0 1 1675
box -3 -3 3 3
use INVX2  INVX2_404
timestamp 1682952543
transform 1 0 2584 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2310
timestamp 1682952543
transform 1 0 2600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1682952543
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1682952543
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1682952543
transform 1 0 2624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2318
timestamp 1682952543
transform 1 0 2632 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5908
timestamp 1682952543
transform 1 0 2668 0 1 1675
box -3 -3 3 3
use OAI21X1  OAI21X1_87
timestamp 1682952543
transform 1 0 2640 0 -1 1770
box -8 -3 34 105
use FILL  FILL_2319
timestamp 1682952543
transform 1 0 2672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1682952543
transform 1 0 2680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2323
timestamp 1682952543
transform 1 0 2688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1682952543
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_406
timestamp 1682952543
transform 1 0 2704 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2328
timestamp 1682952543
transform 1 0 2720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1682952543
transform 1 0 2728 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1682952543
transform 1 0 2736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2343
timestamp 1682952543
transform 1 0 2744 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_50
timestamp 1682952543
transform -1 0 2784 0 -1 1770
box -8 -3 40 105
use FILL  FILL_2344
timestamp 1682952543
transform 1 0 2784 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1682952543
transform 1 0 2792 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1682952543
transform 1 0 2800 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1682952543
transform 1 0 2808 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_51
timestamp 1682952543
transform -1 0 2848 0 -1 1770
box -8 -3 40 105
use FILL  FILL_2348
timestamp 1682952543
transform 1 0 2848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1682952543
transform 1 0 2856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1682952543
transform 1 0 2864 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1682952543
transform 1 0 2872 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1682952543
transform 1 0 2880 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1682952543
transform 1 0 2888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2355
timestamp 1682952543
transform 1 0 2896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1682952543
transform 1 0 2904 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_252
timestamp 1682952543
transform -1 0 2952 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2362
timestamp 1682952543
transform 1 0 2952 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1682952543
transform 1 0 2960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1682952543
transform 1 0 2968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1682952543
transform 1 0 2976 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5909
timestamp 1682952543
transform 1 0 2996 0 1 1675
box -3 -3 3 3
use FILL  FILL_2366
timestamp 1682952543
transform 1 0 2984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2367
timestamp 1682952543
transform 1 0 2992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1682952543
transform 1 0 3000 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5910
timestamp 1682952543
transform 1 0 3036 0 1 1675
box -3 -3 3 3
use OAI22X1  OAI22X1_253
timestamp 1682952543
transform 1 0 3008 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2369
timestamp 1682952543
transform 1 0 3048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2370
timestamp 1682952543
transform 1 0 3056 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1682952543
transform 1 0 3064 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1682952543
transform 1 0 3072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1682952543
transform 1 0 3080 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5911
timestamp 1682952543
transform 1 0 3116 0 1 1675
box -3 -3 3 3
use OAI22X1  OAI22X1_254
timestamp 1682952543
transform 1 0 3088 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2374
timestamp 1682952543
transform 1 0 3128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1682952543
transform 1 0 3136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1682952543
transform 1 0 3144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1682952543
transform 1 0 3152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1682952543
transform 1 0 3160 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_408
timestamp 1682952543
transform 1 0 3168 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2386
timestamp 1682952543
transform 1 0 3184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1682952543
transform 1 0 3192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2388
timestamp 1682952543
transform 1 0 3200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1682952543
transform 1 0 3208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2390
timestamp 1682952543
transform 1 0 3216 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_409
timestamp 1682952543
transform 1 0 3224 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2391
timestamp 1682952543
transform 1 0 3240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1682952543
transform 1 0 3248 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_82
timestamp 1682952543
transform -1 0 3280 0 -1 1770
box -5 -3 28 105
use FILL  FILL_2393
timestamp 1682952543
transform 1 0 3280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1682952543
transform 1 0 3288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1682952543
transform 1 0 3296 0 -1 1770
box -8 -3 16 105
use BUFX2  BUFX2_83
timestamp 1682952543
transform -1 0 3328 0 -1 1770
box -5 -3 28 105
use M3_M2  M3_M2_5912
timestamp 1682952543
transform 1 0 3340 0 1 1675
box -3 -3 3 3
use FILL  FILL_2396
timestamp 1682952543
transform 1 0 3328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2398
timestamp 1682952543
transform 1 0 3336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1682952543
transform 1 0 3344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2404
timestamp 1682952543
transform 1 0 3352 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_241
timestamp 1682952543
transform 1 0 3360 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2405
timestamp 1682952543
transform 1 0 3400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1682952543
transform 1 0 3408 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_411
timestamp 1682952543
transform -1 0 3432 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2407
timestamp 1682952543
transform 1 0 3432 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_56
timestamp 1682952543
transform -1 0 3472 0 -1 1770
box -8 -3 40 105
use M3_M2  M3_M2_5913
timestamp 1682952543
transform 1 0 3500 0 1 1675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_368
timestamp 1682952543
transform 1 0 3472 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_369
timestamp 1682952543
transform 1 0 3568 0 -1 1770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_370
timestamp 1682952543
transform 1 0 3664 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_412
timestamp 1682952543
transform 1 0 3760 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2408
timestamp 1682952543
transform 1 0 3776 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_257
timestamp 1682952543
transform -1 0 3824 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2410
timestamp 1682952543
transform 1 0 3824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1682952543
transform 1 0 3832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1682952543
transform 1 0 3840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1682952543
transform 1 0 3848 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_259
timestamp 1682952543
transform 1 0 3856 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2418
timestamp 1682952543
transform 1 0 3896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1682952543
transform 1 0 3904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2420
timestamp 1682952543
transform 1 0 3912 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_414
timestamp 1682952543
transform 1 0 3920 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2421
timestamp 1682952543
transform 1 0 3936 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1682952543
transform 1 0 3944 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1682952543
transform 1 0 3952 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_261
timestamp 1682952543
transform 1 0 3960 0 -1 1770
box -8 -3 46 105
use FILL  FILL_2429
timestamp 1682952543
transform 1 0 4000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2430
timestamp 1682952543
transform 1 0 4008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1682952543
transform 1 0 4016 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_372
timestamp 1682952543
transform 1 0 4024 0 -1 1770
box -8 -3 104 105
use FILL  FILL_2432
timestamp 1682952543
transform 1 0 4120 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_416
timestamp 1682952543
transform 1 0 4128 0 -1 1770
box -9 -3 26 105
use FILL  FILL_2433
timestamp 1682952543
transform 1 0 4144 0 -1 1770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_49
timestamp 1682952543
transform 1 0 4201 0 1 1670
box -10 -3 10 3
use M3_M2  M3_M2_5962
timestamp 1682952543
transform 1 0 188 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6002
timestamp 1682952543
transform 1 0 116 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6003
timestamp 1682952543
transform 1 0 172 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_5984
timestamp 1682952543
transform 1 0 116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1682952543
transform 1 0 164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5986
timestamp 1682952543
transform 1 0 172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5987
timestamp 1682952543
transform 1 0 188 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5988
timestamp 1682952543
transform 1 0 204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1682952543
transform 1 0 84 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6024
timestamp 1682952543
transform 1 0 212 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_6004
timestamp 1682952543
transform 1 0 284 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6005
timestamp 1682952543
transform 1 0 324 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_5989
timestamp 1682952543
transform 1 0 220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5990
timestamp 1682952543
transform 1 0 228 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1682952543
transform 1 0 284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5992
timestamp 1682952543
transform 1 0 324 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1682952543
transform 1 0 188 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6098
timestamp 1682952543
transform 1 0 196 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6099
timestamp 1682952543
transform 1 0 212 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6074
timestamp 1682952543
transform 1 0 188 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6111
timestamp 1682952543
transform 1 0 164 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6047
timestamp 1682952543
transform 1 0 228 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6100
timestamp 1682952543
transform 1 0 308 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6112
timestamp 1682952543
transform 1 0 212 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6025
timestamp 1682952543
transform 1 0 340 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_5993
timestamp 1682952543
transform 1 0 356 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5994
timestamp 1682952543
transform 1 0 372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6101
timestamp 1682952543
transform 1 0 340 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1682952543
transform 1 0 348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1682952543
transform 1 0 364 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6048
timestamp 1682952543
transform 1 0 372 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_5995
timestamp 1682952543
transform 1 0 388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1682952543
transform 1 0 380 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6075
timestamp 1682952543
transform 1 0 348 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6113
timestamp 1682952543
transform 1 0 364 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5943
timestamp 1682952543
transform 1 0 420 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5963
timestamp 1682952543
transform 1 0 436 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_5996
timestamp 1682952543
transform 1 0 404 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6026
timestamp 1682952543
transform 1 0 412 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5914
timestamp 1682952543
transform 1 0 452 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_6006
timestamp 1682952543
transform 1 0 444 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_5997
timestamp 1682952543
transform 1 0 420 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1682952543
transform 1 0 436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_5999
timestamp 1682952543
transform 1 0 444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6105
timestamp 1682952543
transform 1 0 428 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5944
timestamp 1682952543
transform 1 0 492 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6000
timestamp 1682952543
transform 1 0 476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1682952543
transform 1 0 492 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5924
timestamp 1682952543
transform 1 0 508 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6106
timestamp 1682952543
transform 1 0 508 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5915
timestamp 1682952543
transform 1 0 540 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5916
timestamp 1682952543
transform 1 0 588 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5925
timestamp 1682952543
transform 1 0 532 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5945
timestamp 1682952543
transform 1 0 572 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_6007
timestamp 1682952543
transform 1 0 548 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6008
timestamp 1682952543
transform 1 0 572 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6009
timestamp 1682952543
transform 1 0 612 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6002
timestamp 1682952543
transform 1 0 572 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1682952543
transform 1 0 604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6004
timestamp 1682952543
transform 1 0 612 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6107
timestamp 1682952543
transform 1 0 524 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6049
timestamp 1682952543
transform 1 0 612 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6076
timestamp 1682952543
transform 1 0 604 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5946
timestamp 1682952543
transform 1 0 628 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6005
timestamp 1682952543
transform 1 0 628 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6027
timestamp 1682952543
transform 1 0 644 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1682952543
transform 1 0 668 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6006
timestamp 1682952543
transform 1 0 676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6108
timestamp 1682952543
transform 1 0 660 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1682952543
transform 1 0 668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1682952543
transform 1 0 684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6111
timestamp 1682952543
transform 1 0 692 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6077
timestamp 1682952543
transform 1 0 684 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6180
timestamp 1682952543
transform 1 0 708 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_6114
timestamp 1682952543
transform 1 0 708 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5926
timestamp 1682952543
transform 1 0 740 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6007
timestamp 1682952543
transform 1 0 748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6112
timestamp 1682952543
transform 1 0 756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6008
timestamp 1682952543
transform 1 0 772 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5947
timestamp 1682952543
transform 1 0 820 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6009
timestamp 1682952543
transform 1 0 812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1682952543
transform 1 0 804 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6050
timestamp 1682952543
transform 1 0 812 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1682952543
transform 1 0 828 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6078
timestamp 1682952543
transform 1 0 804 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6010
timestamp 1682952543
transform 1 0 852 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5964
timestamp 1682952543
transform 1 0 884 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6011
timestamp 1682952543
transform 1 0 884 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6114
timestamp 1682952543
transform 1 0 876 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6052
timestamp 1682952543
transform 1 0 884 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6010
timestamp 1682952543
transform 1 0 908 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6012
timestamp 1682952543
transform 1 0 908 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6013
timestamp 1682952543
transform 1 0 924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6115
timestamp 1682952543
transform 1 0 892 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6116
timestamp 1682952543
transform 1 0 932 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6011
timestamp 1682952543
transform 1 0 948 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6117
timestamp 1682952543
transform 1 0 948 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6079
timestamp 1682952543
transform 1 0 940 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5917
timestamp 1682952543
transform 1 0 980 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6181
timestamp 1682952543
transform 1 0 980 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6014
timestamp 1682952543
transform 1 0 996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1682952543
transform 1 0 1028 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6115
timestamp 1682952543
transform 1 0 1028 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6015
timestamp 1682952543
transform 1 0 1068 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6080
timestamp 1682952543
transform 1 0 1068 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5918
timestamp 1682952543
transform 1 0 1084 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5948
timestamp 1682952543
transform 1 0 1084 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6016
timestamp 1682952543
transform 1 0 1092 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5949
timestamp 1682952543
transform 1 0 1108 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_6029
timestamp 1682952543
transform 1 0 1108 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5965
timestamp 1682952543
transform 1 0 1124 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6017
timestamp 1682952543
transform 1 0 1116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6119
timestamp 1682952543
transform 1 0 1108 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5950
timestamp 1682952543
transform 1 0 1148 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_6012
timestamp 1682952543
transform 1 0 1140 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6018
timestamp 1682952543
transform 1 0 1140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6120
timestamp 1682952543
transform 1 0 1132 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6013
timestamp 1682952543
transform 1 0 1164 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6019
timestamp 1682952543
transform 1 0 1164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1682952543
transform 1 0 1164 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6081
timestamp 1682952543
transform 1 0 1164 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_5972
timestamp 1682952543
transform 1 0 1172 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_6030
timestamp 1682952543
transform 1 0 1180 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6122
timestamp 1682952543
transform 1 0 1180 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1682952543
transform 1 0 1220 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6020
timestamp 1682952543
transform 1 0 1212 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6014
timestamp 1682952543
transform 1 0 1236 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5951
timestamp 1682952543
transform 1 0 1276 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6021
timestamp 1682952543
transform 1 0 1276 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1682952543
transform 1 0 1300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6123
timestamp 1682952543
transform 1 0 1268 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6053
timestamp 1682952543
transform 1 0 1276 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6124
timestamp 1682952543
transform 1 0 1292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1682952543
transform 1 0 1308 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6082
timestamp 1682952543
transform 1 0 1292 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5952
timestamp 1682952543
transform 1 0 1324 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5966
timestamp 1682952543
transform 1 0 1332 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6054
timestamp 1682952543
transform 1 0 1340 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1682952543
transform 1 0 1396 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_6031
timestamp 1682952543
transform 1 0 1356 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5920
timestamp 1682952543
transform 1 0 1540 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1682952543
transform 1 0 1516 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5921
timestamp 1682952543
transform 1 0 1572 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5953
timestamp 1682952543
transform 1 0 1500 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5954
timestamp 1682952543
transform 1 0 1532 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5955
timestamp 1682952543
transform 1 0 1548 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6023
timestamp 1682952543
transform 1 0 1380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1682952543
transform 1 0 1436 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6025
timestamp 1682952543
transform 1 0 1500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1682952543
transform 1 0 1356 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6083
timestamp 1682952543
transform 1 0 1380 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6084
timestamp 1682952543
transform 1 0 1396 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6032
timestamp 1682952543
transform 1 0 1524 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1682952543
transform 1 0 1548 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5968
timestamp 1682952543
transform 1 0 1564 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6015
timestamp 1682952543
transform 1 0 1556 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6026
timestamp 1682952543
transform 1 0 1532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1682952543
transform 1 0 1556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6127
timestamp 1682952543
transform 1 0 1452 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6055
timestamp 1682952543
transform 1 0 1524 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6128
timestamp 1682952543
transform 1 0 1540 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6129
timestamp 1682952543
transform 1 0 1548 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6130
timestamp 1682952543
transform 1 0 1564 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6033
timestamp 1682952543
transform 1 0 1580 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6028
timestamp 1682952543
transform 1 0 1588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6131
timestamp 1682952543
transform 1 0 1580 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6085
timestamp 1682952543
transform 1 0 1580 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1682952543
transform 1 0 1596 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6029
timestamp 1682952543
transform 1 0 1604 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5956
timestamp 1682952543
transform 1 0 1628 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5969
timestamp 1682952543
transform 1 0 1636 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6030
timestamp 1682952543
transform 1 0 1628 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1682952543
transform 1 0 1636 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5928
timestamp 1682952543
transform 1 0 1684 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6031
timestamp 1682952543
transform 1 0 1676 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6057
timestamp 1682952543
transform 1 0 1668 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6182
timestamp 1682952543
transform 1 0 1652 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_6086
timestamp 1682952543
transform 1 0 1660 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5957
timestamp 1682952543
transform 1 0 1708 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5929
timestamp 1682952543
transform 1 0 1724 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6032
timestamp 1682952543
transform 1 0 1708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1682952543
transform 1 0 1716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6133
timestamp 1682952543
transform 1 0 1700 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6087
timestamp 1682952543
transform 1 0 1716 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6034
timestamp 1682952543
transform 1 0 1732 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6134
timestamp 1682952543
transform 1 0 1732 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5970
timestamp 1682952543
transform 1 0 1756 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6135
timestamp 1682952543
transform 1 0 1772 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5922
timestamp 1682952543
transform 1 0 1788 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_5974
timestamp 1682952543
transform 1 0 1788 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6136
timestamp 1682952543
transform 1 0 1780 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6088
timestamp 1682952543
transform 1 0 1780 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5971
timestamp 1682952543
transform 1 0 1828 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6016
timestamp 1682952543
transform 1 0 1820 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6034
timestamp 1682952543
transform 1 0 1836 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6137
timestamp 1682952543
transform 1 0 1852 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5972
timestamp 1682952543
transform 1 0 1876 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6116
timestamp 1682952543
transform 1 0 1860 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1682952543
transform 1 0 1892 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5973
timestamp 1682952543
transform 1 0 2004 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6017
timestamp 1682952543
transform 1 0 1940 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6018
timestamp 1682952543
transform 1 0 1980 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6035
timestamp 1682952543
transform 1 0 1892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6036
timestamp 1682952543
transform 1 0 1900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1682952543
transform 1 0 1916 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1682952543
transform 1 0 1932 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6058
timestamp 1682952543
transform 1 0 1892 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6138
timestamp 1682952543
transform 1 0 1900 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6139
timestamp 1682952543
transform 1 0 1908 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6035
timestamp 1682952543
transform 1 0 1940 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6039
timestamp 1682952543
transform 1 0 1980 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6036
timestamp 1682952543
transform 1 0 2028 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6040
timestamp 1682952543
transform 1 0 2036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6140
timestamp 1682952543
transform 1 0 1940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1682952543
transform 1 0 1956 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6059
timestamp 1682952543
transform 1 0 1980 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6060
timestamp 1682952543
transform 1 0 1996 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6089
timestamp 1682952543
transform 1 0 2004 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6090
timestamp 1682952543
transform 1 0 2028 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5974
timestamp 1682952543
transform 1 0 2068 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_5975
timestamp 1682952543
transform 1 0 2076 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1682952543
transform 1 0 2060 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6061
timestamp 1682952543
transform 1 0 2060 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6142
timestamp 1682952543
transform 1 0 2084 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5975
timestamp 1682952543
transform 1 0 2100 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6183
timestamp 1682952543
transform 1 0 2092 0 1 1595
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1682952543
transform 1 0 2116 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5976
timestamp 1682952543
transform 1 0 2132 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1682952543
transform 1 0 2172 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5931
timestamp 1682952543
transform 1 0 2188 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6043
timestamp 1682952543
transform 1 0 2188 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6144
timestamp 1682952543
transform 1 0 2180 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5976
timestamp 1682952543
transform 1 0 2292 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6019
timestamp 1682952543
transform 1 0 2244 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6020
timestamp 1682952543
transform 1 0 2300 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6021
timestamp 1682952543
transform 1 0 2388 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6044
timestamp 1682952543
transform 1 0 2252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1682952543
transform 1 0 2284 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6046
timestamp 1682952543
transform 1 0 2348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1682952543
transform 1 0 2380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1682952543
transform 1 0 2388 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6145
timestamp 1682952543
transform 1 0 2204 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6091
timestamp 1682952543
transform 1 0 2204 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6146
timestamp 1682952543
transform 1 0 2300 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6062
timestamp 1682952543
transform 1 0 2348 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6063
timestamp 1682952543
transform 1 0 2388 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6092
timestamp 1682952543
transform 1 0 2300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6093
timestamp 1682952543
transform 1 0 2380 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6049
timestamp 1682952543
transform 1 0 2404 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6117
timestamp 1682952543
transform 1 0 2404 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6037
timestamp 1682952543
transform 1 0 2420 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6050
timestamp 1682952543
transform 1 0 2428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1682952543
transform 1 0 2420 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1682952543
transform 1 0 2428 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6094
timestamp 1682952543
transform 1 0 2428 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_5977
timestamp 1682952543
transform 1 0 2460 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6149
timestamp 1682952543
transform 1 0 2468 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6095
timestamp 1682952543
transform 1 0 2468 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6118
timestamp 1682952543
transform 1 0 2468 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5932
timestamp 1682952543
transform 1 0 2516 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6051
timestamp 1682952543
transform 1 0 2484 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1682952543
transform 1 0 2492 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6038
timestamp 1682952543
transform 1 0 2500 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6053
timestamp 1682952543
transform 1 0 2508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1682952543
transform 1 0 2524 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5977
timestamp 1682952543
transform 1 0 2540 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6039
timestamp 1682952543
transform 1 0 2548 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6150
timestamp 1682952543
transform 1 0 2548 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5933
timestamp 1682952543
transform 1 0 2564 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5978
timestamp 1682952543
transform 1 0 2580 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6055
timestamp 1682952543
transform 1 0 2572 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6040
timestamp 1682952543
transform 1 0 2580 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6056
timestamp 1682952543
transform 1 0 2588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6151
timestamp 1682952543
transform 1 0 2564 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6096
timestamp 1682952543
transform 1 0 2564 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1682952543
transform 1 0 2644 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5979
timestamp 1682952543
transform 1 0 2636 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6057
timestamp 1682952543
transform 1 0 2620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6058
timestamp 1682952543
transform 1 0 2636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1682952543
transform 1 0 2652 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6119
timestamp 1682952543
transform 1 0 2612 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6064
timestamp 1682952543
transform 1 0 2628 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6152
timestamp 1682952543
transform 1 0 2644 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1682952543
transform 1 0 2652 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6120
timestamp 1682952543
transform 1 0 2636 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5980
timestamp 1682952543
transform 1 0 2684 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6097
timestamp 1682952543
transform 1 0 2692 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5935
timestamp 1682952543
transform 1 0 2716 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5981
timestamp 1682952543
transform 1 0 2708 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5982
timestamp 1682952543
transform 1 0 2748 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5983
timestamp 1682952543
transform 1 0 2804 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6060
timestamp 1682952543
transform 1 0 2708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1682952543
transform 1 0 2716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1682952543
transform 1 0 2748 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6041
timestamp 1682952543
transform 1 0 2796 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6154
timestamp 1682952543
transform 1 0 2796 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6098
timestamp 1682952543
transform 1 0 2796 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5984
timestamp 1682952543
transform 1 0 2836 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5958
timestamp 1682952543
transform 1 0 2852 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_5969
timestamp 1682952543
transform 1 0 2852 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5985
timestamp 1682952543
transform 1 0 2860 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_5978
timestamp 1682952543
transform 1 0 2844 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1682952543
transform 1 0 2868 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6063
timestamp 1682952543
transform 1 0 2860 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1682952543
transform 1 0 2900 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6065
timestamp 1682952543
transform 1 0 2908 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5986
timestamp 1682952543
transform 1 0 2940 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5987
timestamp 1682952543
transform 1 0 2956 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6065
timestamp 1682952543
transform 1 0 2940 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1682952543
transform 1 0 2956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6155
timestamp 1682952543
transform 1 0 2932 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5988
timestamp 1682952543
transform 1 0 2988 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6156
timestamp 1682952543
transform 1 0 2996 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5936
timestamp 1682952543
transform 1 0 3012 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5937
timestamp 1682952543
transform 1 0 3060 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6067
timestamp 1682952543
transform 1 0 3036 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1682952543
transform 1 0 3012 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6066
timestamp 1682952543
transform 1 0 3076 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6067
timestamp 1682952543
transform 1 0 3092 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6099
timestamp 1682952543
transform 1 0 3012 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6068
timestamp 1682952543
transform 1 0 3116 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6068
timestamp 1682952543
transform 1 0 3116 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5989
timestamp 1682952543
transform 1 0 3140 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6069
timestamp 1682952543
transform 1 0 3140 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1682952543
transform 1 0 3156 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6158
timestamp 1682952543
transform 1 0 3132 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6100
timestamp 1682952543
transform 1 0 3148 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5990
timestamp 1682952543
transform 1 0 3212 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5991
timestamp 1682952543
transform 1 0 3244 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6071
timestamp 1682952543
transform 1 0 3212 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1682952543
transform 1 0 3220 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6073
timestamp 1682952543
transform 1 0 3236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6159
timestamp 1682952543
transform 1 0 3204 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6160
timestamp 1682952543
transform 1 0 3212 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6101
timestamp 1682952543
transform 1 0 3204 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6069
timestamp 1682952543
transform 1 0 3220 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6161
timestamp 1682952543
transform 1 0 3228 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6102
timestamp 1682952543
transform 1 0 3236 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_5980
timestamp 1682952543
transform 1 0 3252 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5938
timestamp 1682952543
transform 1 0 3276 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5959
timestamp 1682952543
transform 1 0 3268 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_5970
timestamp 1682952543
transform 1 0 3268 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5992
timestamp 1682952543
transform 1 0 3300 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_5981
timestamp 1682952543
transform 1 0 3284 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_6042
timestamp 1682952543
transform 1 0 3252 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_6043
timestamp 1682952543
transform 1 0 3268 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6074
timestamp 1682952543
transform 1 0 3276 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6044
timestamp 1682952543
transform 1 0 3292 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6075
timestamp 1682952543
transform 1 0 3300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6076
timestamp 1682952543
transform 1 0 3316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6162
timestamp 1682952543
transform 1 0 3252 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6121
timestamp 1682952543
transform 1 0 3252 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6070
timestamp 1682952543
transform 1 0 3284 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5939
timestamp 1682952543
transform 1 0 3380 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5993
timestamp 1682952543
transform 1 0 3404 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6077
timestamp 1682952543
transform 1 0 3364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6163
timestamp 1682952543
transform 1 0 3292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1682952543
transform 1 0 3308 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6165
timestamp 1682952543
transform 1 0 3324 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1682952543
transform 1 0 3340 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6103
timestamp 1682952543
transform 1 0 3308 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6071
timestamp 1682952543
transform 1 0 3372 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6104
timestamp 1682952543
transform 1 0 3364 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6105
timestamp 1682952543
transform 1 0 3404 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6122
timestamp 1682952543
transform 1 0 3388 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5940
timestamp 1682952543
transform 1 0 3436 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6078
timestamp 1682952543
transform 1 0 3436 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5994
timestamp 1682952543
transform 1 0 3468 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6079
timestamp 1682952543
transform 1 0 3460 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5995
timestamp 1682952543
transform 1 0 3524 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_5982
timestamp 1682952543
transform 1 0 3524 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1682952543
transform 1 0 3500 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1682952543
transform 1 0 3516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6167
timestamp 1682952543
transform 1 0 3492 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6106
timestamp 1682952543
transform 1 0 3508 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6168
timestamp 1682952543
transform 1 0 3532 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1682952543
transform 1 0 3620 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1682952543
transform 1 0 3628 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6045
timestamp 1682952543
transform 1 0 3636 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6083
timestamp 1682952543
transform 1 0 3644 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5941
timestamp 1682952543
transform 1 0 3676 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_5983
timestamp 1682952543
transform 1 0 3668 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5996
timestamp 1682952543
transform 1 0 3700 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6084
timestamp 1682952543
transform 1 0 3700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6169
timestamp 1682952543
transform 1 0 3676 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6170
timestamp 1682952543
transform 1 0 3692 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6107
timestamp 1682952543
transform 1 0 3668 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6072
timestamp 1682952543
transform 1 0 3700 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1682952543
transform 1 0 3732 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5997
timestamp 1682952543
transform 1 0 3724 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6085
timestamp 1682952543
transform 1 0 3716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1682952543
transform 1 0 3708 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6123
timestamp 1682952543
transform 1 0 3708 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6073
timestamp 1682952543
transform 1 0 3724 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_6108
timestamp 1682952543
transform 1 0 3724 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6172
timestamp 1682952543
transform 1 0 3740 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5961
timestamp 1682952543
transform 1 0 3764 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5942
timestamp 1682952543
transform 1 0 3852 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5998
timestamp 1682952543
transform 1 0 3812 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6086
timestamp 1682952543
transform 1 0 3812 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1682952543
transform 1 0 3772 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6124
timestamp 1682952543
transform 1 0 3860 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5999
timestamp 1682952543
transform 1 0 3876 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6087
timestamp 1682952543
transform 1 0 3884 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6088
timestamp 1682952543
transform 1 0 3892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1682952543
transform 1 0 3908 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_6046
timestamp 1682952543
transform 1 0 3916 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6090
timestamp 1682952543
transform 1 0 3924 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1682952543
transform 1 0 3940 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6174
timestamp 1682952543
transform 1 0 3932 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1682952543
transform 1 0 3940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6176
timestamp 1682952543
transform 1 0 3948 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6000
timestamp 1682952543
transform 1 0 3964 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6001
timestamp 1682952543
transform 1 0 3996 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_6022
timestamp 1682952543
transform 1 0 3996 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6092
timestamp 1682952543
transform 1 0 3980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1682952543
transform 1 0 3996 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6177
timestamp 1682952543
transform 1 0 3988 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1682952543
transform 1 0 4004 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6109
timestamp 1682952543
transform 1 0 3988 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6125
timestamp 1682952543
transform 1 0 4004 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_6126
timestamp 1682952543
transform 1 0 4020 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1682952543
transform 1 0 4076 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6094
timestamp 1682952543
transform 1 0 4076 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6179
timestamp 1682952543
transform 1 0 4052 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_6110
timestamp 1682952543
transform 1 0 4076 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_6023
timestamp 1682952543
transform 1 0 4148 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6095
timestamp 1682952543
transform 1 0 4148 0 1 1615
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_50
timestamp 1682952543
transform 1 0 48 0 1 1570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_373
timestamp 1682952543
transform 1 0 72 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_417
timestamp 1682952543
transform -1 0 184 0 1 1570
box -9 -3 26 105
use M3_M2  M3_M2_6127
timestamp 1682952543
transform 1 0 196 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_244
timestamp 1682952543
transform 1 0 184 0 1 1570
box -8 -3 46 105
use M3_M2  M3_M2_6128
timestamp 1682952543
transform 1 0 244 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6129
timestamp 1682952543
transform 1 0 260 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_375
timestamp 1682952543
transform -1 0 320 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_418
timestamp 1682952543
transform -1 0 336 0 1 1570
box -9 -3 26 105
use FILL  FILL_2434
timestamp 1682952543
transform 1 0 336 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_262
timestamp 1682952543
transform -1 0 384 0 1 1570
box -8 -3 46 105
use FILL  FILL_2435
timestamp 1682952543
transform 1 0 384 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6130
timestamp 1682952543
transform 1 0 404 0 1 1575
box -3 -3 3 3
use FILL  FILL_2436
timestamp 1682952543
transform 1 0 392 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_245
timestamp 1682952543
transform -1 0 440 0 1 1570
box -8 -3 46 105
use FILL  FILL_2437
timestamp 1682952543
transform 1 0 440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2438
timestamp 1682952543
transform 1 0 448 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_246
timestamp 1682952543
transform 1 0 456 0 1 1570
box -8 -3 46 105
use FILL  FILL_2439
timestamp 1682952543
transform 1 0 496 0 1 1570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1682952543
transform 1 0 504 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_376
timestamp 1682952543
transform 1 0 512 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_419
timestamp 1682952543
transform -1 0 624 0 1 1570
box -9 -3 26 105
use FILL  FILL_2441
timestamp 1682952543
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1682952543
transform 1 0 632 0 1 1570
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1682952543
transform 1 0 640 0 1 1570
box -8 -3 16 105
use FILL  FILL_2444
timestamp 1682952543
transform 1 0 648 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_247
timestamp 1682952543
transform 1 0 656 0 1 1570
box -8 -3 46 105
use FILL  FILL_2445
timestamp 1682952543
transform 1 0 696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1682952543
transform 1 0 704 0 1 1570
box -8 -3 16 105
use FILL  FILL_2470
timestamp 1682952543
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1682952543
transform 1 0 720 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_78
timestamp 1682952543
transform 1 0 728 0 1 1570
box -8 -3 32 105
use FILL  FILL_2472
timestamp 1682952543
transform 1 0 752 0 1 1570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1682952543
transform 1 0 760 0 1 1570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1682952543
transform 1 0 768 0 1 1570
box -8 -3 16 105
use FILL  FILL_2477
timestamp 1682952543
transform 1 0 776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1682952543
transform 1 0 784 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_251
timestamp 1682952543
transform 1 0 792 0 1 1570
box -8 -3 46 105
use FILL  FILL_2479
timestamp 1682952543
transform 1 0 832 0 1 1570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1682952543
transform 1 0 840 0 1 1570
box -8 -3 16 105
use FILL  FILL_2484
timestamp 1682952543
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1682952543
transform 1 0 856 0 1 1570
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1682952543
transform 1 0 864 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6131
timestamp 1682952543
transform 1 0 884 0 1 1575
box -3 -3 3 3
use FILL  FILL_2487
timestamp 1682952543
transform 1 0 872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1682952543
transform 1 0 880 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6132
timestamp 1682952543
transform 1 0 908 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6133
timestamp 1682952543
transform 1 0 924 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_252
timestamp 1682952543
transform 1 0 888 0 1 1570
box -8 -3 46 105
use FILL  FILL_2489
timestamp 1682952543
transform 1 0 928 0 1 1570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1682952543
transform 1 0 936 0 1 1570
box -8 -3 16 105
use FILL  FILL_2493
timestamp 1682952543
transform 1 0 944 0 1 1570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1682952543
transform 1 0 952 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_424
timestamp 1682952543
transform 1 0 960 0 1 1570
box -9 -3 26 105
use FILL  FILL_2495
timestamp 1682952543
transform 1 0 976 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6134
timestamp 1682952543
transform 1 0 996 0 1 1575
box -3 -3 3 3
use FILL  FILL_2496
timestamp 1682952543
transform 1 0 984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2497
timestamp 1682952543
transform 1 0 992 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6135
timestamp 1682952543
transform 1 0 1012 0 1 1575
box -3 -3 3 3
use FILL  FILL_2498
timestamp 1682952543
transform 1 0 1000 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_80
timestamp 1682952543
transform 1 0 1008 0 1 1570
box -8 -3 32 105
use FILL  FILL_2499
timestamp 1682952543
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1682952543
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1682952543
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use FILL  FILL_2502
timestamp 1682952543
transform 1 0 1056 0 1 1570
box -8 -3 16 105
use FILL  FILL_2503
timestamp 1682952543
transform 1 0 1064 0 1 1570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1682952543
transform 1 0 1072 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_425
timestamp 1682952543
transform -1 0 1096 0 1 1570
box -9 -3 26 105
use FILL  FILL_2507
timestamp 1682952543
transform 1 0 1096 0 1 1570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1682952543
transform 1 0 1104 0 1 1570
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1682952543
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1682952543
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1682952543
transform 1 0 1128 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_91
timestamp 1682952543
transform 1 0 1136 0 1 1570
box -8 -3 34 105
use FILL  FILL_2516
timestamp 1682952543
transform 1 0 1168 0 1 1570
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1682952543
transform 1 0 1176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1682952543
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1682952543
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_61
timestamp 1682952543
transform 1 0 1200 0 1 1570
box -8 -3 32 105
use FILL  FILL_2520
timestamp 1682952543
transform 1 0 1224 0 1 1570
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1682952543
transform 1 0 1232 0 1 1570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1682952543
transform 1 0 1240 0 1 1570
box -8 -3 16 105
use FILL  FILL_2531
timestamp 1682952543
transform 1 0 1248 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6136
timestamp 1682952543
transform 1 0 1268 0 1 1575
box -3 -3 3 3
use FILL  FILL_2533
timestamp 1682952543
transform 1 0 1256 0 1 1570
box -8 -3 16 105
use FILL  FILL_2535
timestamp 1682952543
transform 1 0 1264 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_265
timestamp 1682952543
transform 1 0 1272 0 1 1570
box -8 -3 46 105
use FILL  FILL_2536
timestamp 1682952543
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1682952543
transform 1 0 1320 0 1 1570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1682952543
transform 1 0 1328 0 1 1570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1682952543
transform 1 0 1336 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_379
timestamp 1682952543
transform 1 0 1344 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_6137
timestamp 1682952543
transform 1 0 1516 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6138
timestamp 1682952543
transform 1 0 1532 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_380
timestamp 1682952543
transform 1 0 1440 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_6139
timestamp 1682952543
transform 1 0 1564 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_255
timestamp 1682952543
transform 1 0 1536 0 1 1570
box -8 -3 46 105
use FILL  FILL_2540
timestamp 1682952543
transform 1 0 1576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1682952543
transform 1 0 1584 0 1 1570
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1682952543
transform 1 0 1592 0 1 1570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1682952543
transform 1 0 1600 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6140
timestamp 1682952543
transform 1 0 1636 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_256
timestamp 1682952543
transform -1 0 1648 0 1 1570
box -8 -3 46 105
use FILL  FILL_2544
timestamp 1682952543
transform 1 0 1648 0 1 1570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1682952543
transform 1 0 1656 0 1 1570
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1682952543
transform 1 0 1664 0 1 1570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1682952543
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1682952543
transform 1 0 1680 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_82
timestamp 1682952543
transform 1 0 1688 0 1 1570
box -8 -3 32 105
use FILL  FILL_2560
timestamp 1682952543
transform 1 0 1712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1682952543
transform 1 0 1720 0 1 1570
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1682952543
transform 1 0 1728 0 1 1570
box -8 -3 16 105
use FILL  FILL_2565
timestamp 1682952543
transform 1 0 1736 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_95
timestamp 1682952543
transform 1 0 1744 0 1 1570
box -8 -3 34 105
use FILL  FILL_2567
timestamp 1682952543
transform 1 0 1776 0 1 1570
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1682952543
transform 1 0 1784 0 1 1570
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1682952543
transform 1 0 1792 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6141
timestamp 1682952543
transform 1 0 1812 0 1 1575
box -3 -3 3 3
use BUFX2  BUFX2_85
timestamp 1682952543
transform -1 0 1824 0 1 1570
box -5 -3 28 105
use FILL  FILL_2570
timestamp 1682952543
transform 1 0 1824 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_86
timestamp 1682952543
transform 1 0 1832 0 1 1570
box -5 -3 28 105
use FILL  FILL_2571
timestamp 1682952543
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6142
timestamp 1682952543
transform 1 0 1884 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_429
timestamp 1682952543
transform -1 0 1880 0 1 1570
box -9 -3 26 105
use FILL  FILL_2572
timestamp 1682952543
transform 1 0 1880 0 1 1570
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1682952543
transform 1 0 1888 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_258
timestamp 1682952543
transform 1 0 1896 0 1 1570
box -8 -3 46 105
use FILL  FILL_2574
timestamp 1682952543
transform 1 0 1936 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_383
timestamp 1682952543
transform 1 0 1944 0 1 1570
box -8 -3 104 105
use FILL  FILL_2575
timestamp 1682952543
transform 1 0 2040 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_96
timestamp 1682952543
transform 1 0 2048 0 1 1570
box -8 -3 34 105
use FILL  FILL_2576
timestamp 1682952543
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1682952543
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1682952543
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_83
timestamp 1682952543
transform 1 0 2104 0 1 1570
box -8 -3 32 105
use FILL  FILL_2595
timestamp 1682952543
transform 1 0 2128 0 1 1570
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1682952543
transform 1 0 2136 0 1 1570
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1682952543
transform 1 0 2144 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_102
timestamp 1682952543
transform -1 0 2184 0 1 1570
box -8 -3 34 105
use FILL  FILL_2600
timestamp 1682952543
transform 1 0 2184 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6143
timestamp 1682952543
transform 1 0 2220 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6144
timestamp 1682952543
transform 1 0 2236 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6145
timestamp 1682952543
transform 1 0 2268 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_384
timestamp 1682952543
transform 1 0 2192 0 1 1570
box -8 -3 104 105
use M3_M2  M3_M2_6146
timestamp 1682952543
transform 1 0 2308 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6147
timestamp 1682952543
transform 1 0 2332 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6148
timestamp 1682952543
transform 1 0 2380 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_385
timestamp 1682952543
transform 1 0 2288 0 1 1570
box -8 -3 104 105
use FILL  FILL_2601
timestamp 1682952543
transform 1 0 2384 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_431
timestamp 1682952543
transform -1 0 2408 0 1 1570
box -9 -3 26 105
use FILL  FILL_2602
timestamp 1682952543
transform 1 0 2408 0 1 1570
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1682952543
transform 1 0 2416 0 1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_107
timestamp 1682952543
transform 1 0 2424 0 1 1570
box -8 -3 34 105
use FILL  FILL_2621
timestamp 1682952543
transform 1 0 2456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1682952543
transform 1 0 2464 0 1 1570
box -8 -3 16 105
use FILL  FILL_2625
timestamp 1682952543
transform 1 0 2472 0 1 1570
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1682952543
transform 1 0 2480 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_259
timestamp 1682952543
transform -1 0 2528 0 1 1570
box -8 -3 46 105
use FILL  FILL_2628
timestamp 1682952543
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1682952543
transform 1 0 2536 0 1 1570
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1682952543
transform 1 0 2544 0 1 1570
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1682952543
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use AND2X2  AND2X2_48
timestamp 1682952543
transform 1 0 2560 0 1 1570
box -8 -3 40 105
use FILL  FILL_2636
timestamp 1682952543
transform 1 0 2592 0 1 1570
box -8 -3 16 105
use FILL  FILL_2637
timestamp 1682952543
transform 1 0 2600 0 1 1570
box -8 -3 16 105
use FILL  FILL_2638
timestamp 1682952543
transform 1 0 2608 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_260
timestamp 1682952543
transform 1 0 2616 0 1 1570
box -8 -3 46 105
use FILL  FILL_2639
timestamp 1682952543
transform 1 0 2656 0 1 1570
box -8 -3 16 105
use FILL  FILL_2640
timestamp 1682952543
transform 1 0 2664 0 1 1570
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1682952543
transform 1 0 2672 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_432
timestamp 1682952543
transform 1 0 2680 0 1 1570
box -9 -3 26 105
use FILL  FILL_2642
timestamp 1682952543
transform 1 0 2696 0 1 1570
box -8 -3 16 105
use FILL  FILL_2651
timestamp 1682952543
transform 1 0 2704 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6149
timestamp 1682952543
transform 1 0 2756 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_386
timestamp 1682952543
transform -1 0 2808 0 1 1570
box -8 -3 104 105
use FILL  FILL_2652
timestamp 1682952543
transform 1 0 2808 0 1 1570
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1682952543
transform 1 0 2816 0 1 1570
box -8 -3 16 105
use FILL  FILL_2654
timestamp 1682952543
transform 1 0 2824 0 1 1570
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1682952543
transform 1 0 2832 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_58
timestamp 1682952543
transform -1 0 2872 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_6150
timestamp 1682952543
transform 1 0 2884 0 1 1575
box -3 -3 3 3
use FILL  FILL_2659
timestamp 1682952543
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1682952543
transform 1 0 2880 0 1 1570
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1682952543
transform 1 0 2888 0 1 1570
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1682952543
transform 1 0 2896 0 1 1570
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1682952543
transform 1 0 2904 0 1 1570
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1682952543
transform 1 0 2912 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_262
timestamp 1682952543
transform 1 0 2920 0 1 1570
box -8 -3 46 105
use FILL  FILL_2669
timestamp 1682952543
transform 1 0 2960 0 1 1570
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1682952543
transform 1 0 2968 0 1 1570
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1682952543
transform 1 0 2976 0 1 1570
box -8 -3 16 105
use FILL  FILL_2672
timestamp 1682952543
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1682952543
transform 1 0 2992 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_387
timestamp 1682952543
transform 1 0 3000 0 1 1570
box -8 -3 104 105
use FILL  FILL_2674
timestamp 1682952543
transform 1 0 3096 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6151
timestamp 1682952543
transform 1 0 3124 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_433
timestamp 1682952543
transform 1 0 3104 0 1 1570
box -9 -3 26 105
use FILL  FILL_2675
timestamp 1682952543
transform 1 0 3120 0 1 1570
box -8 -3 16 105
use FILL  FILL_2676
timestamp 1682952543
transform 1 0 3128 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6152
timestamp 1682952543
transform 1 0 3180 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_263
timestamp 1682952543
transform -1 0 3176 0 1 1570
box -8 -3 46 105
use M3_M2  M3_M2_6153
timestamp 1682952543
transform 1 0 3196 0 1 1575
box -3 -3 3 3
use FILL  FILL_2677
timestamp 1682952543
transform 1 0 3176 0 1 1570
box -8 -3 16 105
use FILL  FILL_2678
timestamp 1682952543
transform 1 0 3184 0 1 1570
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1682952543
transform 1 0 3192 0 1 1570
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1682952543
transform 1 0 3200 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6154
timestamp 1682952543
transform 1 0 3228 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_268
timestamp 1682952543
transform 1 0 3208 0 1 1570
box -8 -3 46 105
use FILL  FILL_2681
timestamp 1682952543
transform 1 0 3248 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6155
timestamp 1682952543
transform 1 0 3292 0 1 1575
box -3 -3 3 3
use NAND3X1  NAND3X1_59
timestamp 1682952543
transform -1 0 3288 0 1 1570
box -8 -3 40 105
use OAI22X1  OAI22X1_269
timestamp 1682952543
transform 1 0 3288 0 1 1570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_388
timestamp 1682952543
transform 1 0 3328 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_434
timestamp 1682952543
transform 1 0 3424 0 1 1570
box -9 -3 26 105
use FILL  FILL_2682
timestamp 1682952543
transform 1 0 3440 0 1 1570
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1682952543
transform 1 0 3448 0 1 1570
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1682952543
transform 1 0 3456 0 1 1570
box -8 -3 16 105
use FILL  FILL_2685
timestamp 1682952543
transform 1 0 3464 0 1 1570
box -8 -3 16 105
use FILL  FILL_2703
timestamp 1682952543
transform 1 0 3472 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_266
timestamp 1682952543
transform 1 0 3480 0 1 1570
box -8 -3 46 105
use FILL  FILL_2705
timestamp 1682952543
transform 1 0 3520 0 1 1570
box -8 -3 16 105
use FILL  FILL_2712
timestamp 1682952543
transform 1 0 3528 0 1 1570
box -8 -3 16 105
use FILL  FILL_2714
timestamp 1682952543
transform 1 0 3536 0 1 1570
box -8 -3 16 105
use FILL  FILL_2715
timestamp 1682952543
transform 1 0 3544 0 1 1570
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1682952543
transform 1 0 3552 0 1 1570
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1682952543
transform 1 0 3560 0 1 1570
box -8 -3 16 105
use FILL  FILL_2720
timestamp 1682952543
transform 1 0 3568 0 1 1570
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1682952543
transform 1 0 3576 0 1 1570
box -8 -3 16 105
use FILL  FILL_2723
timestamp 1682952543
transform 1 0 3584 0 1 1570
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1682952543
transform 1 0 3592 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6156
timestamp 1682952543
transform 1 0 3612 0 1 1575
box -3 -3 3 3
use FILL  FILL_2725
timestamp 1682952543
transform 1 0 3600 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_61
timestamp 1682952543
transform -1 0 3640 0 1 1570
box -8 -3 40 105
use FILL  FILL_2726
timestamp 1682952543
transform 1 0 3640 0 1 1570
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1682952543
transform 1 0 3648 0 1 1570
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1682952543
transform 1 0 3656 0 1 1570
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1682952543
transform 1 0 3664 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6157
timestamp 1682952543
transform 1 0 3708 0 1 1575
box -3 -3 3 3
use OAI22X1  OAI22X1_272
timestamp 1682952543
transform 1 0 3672 0 1 1570
box -8 -3 46 105
use FILL  FILL_2735
timestamp 1682952543
transform 1 0 3712 0 1 1570
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1682952543
transform 1 0 3720 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_438
timestamp 1682952543
transform -1 0 3744 0 1 1570
box -9 -3 26 105
use FILL  FILL_2737
timestamp 1682952543
transform 1 0 3744 0 1 1570
box -8 -3 16 105
use FILL  FILL_2738
timestamp 1682952543
transform 1 0 3752 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6158
timestamp 1682952543
transform 1 0 3788 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_6159
timestamp 1682952543
transform 1 0 3844 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_391
timestamp 1682952543
transform 1 0 3760 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_439
timestamp 1682952543
transform 1 0 3856 0 1 1570
box -9 -3 26 105
use FILL  FILL_2739
timestamp 1682952543
transform 1 0 3872 0 1 1570
box -8 -3 16 105
use FILL  FILL_2740
timestamp 1682952543
transform 1 0 3880 0 1 1570
box -8 -3 16 105
use FILL  FILL_2741
timestamp 1682952543
transform 1 0 3888 0 1 1570
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1682952543
transform 1 0 3896 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6160
timestamp 1682952543
transform 1 0 3924 0 1 1575
box -3 -3 3 3
use AOI22X1  AOI22X1_267
timestamp 1682952543
transform -1 0 3944 0 1 1570
box -8 -3 46 105
use FILL  FILL_2743
timestamp 1682952543
transform 1 0 3944 0 1 1570
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1682952543
transform 1 0 3952 0 1 1570
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1682952543
transform 1 0 3960 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_273
timestamp 1682952543
transform 1 0 3968 0 1 1570
box -8 -3 46 105
use FILL  FILL_2746
timestamp 1682952543
transform 1 0 4008 0 1 1570
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1682952543
transform 1 0 4016 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6161
timestamp 1682952543
transform 1 0 4036 0 1 1575
box -3 -3 3 3
use FILL  FILL_2748
timestamp 1682952543
transform 1 0 4024 0 1 1570
box -8 -3 16 105
use FILL  FILL_2749
timestamp 1682952543
transform 1 0 4032 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6162
timestamp 1682952543
transform 1 0 4052 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_392
timestamp 1682952543
transform 1 0 4040 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_440
timestamp 1682952543
transform 1 0 4136 0 1 1570
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_51
timestamp 1682952543
transform 1 0 4177 0 1 1570
box -10 -3 10 3
use M3_M2  M3_M2_6211
timestamp 1682952543
transform 1 0 164 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6186
timestamp 1682952543
transform 1 0 84 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6246
timestamp 1682952543
transform 1 0 116 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6299
timestamp 1682952543
transform 1 0 116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1682952543
transform 1 0 164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1682952543
transform 1 0 172 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6163
timestamp 1682952543
transform 1 0 196 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6302
timestamp 1682952543
transform 1 0 196 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6164
timestamp 1682952543
transform 1 0 220 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6212
timestamp 1682952543
transform 1 0 220 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6187
timestamp 1682952543
transform 1 0 212 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6188
timestamp 1682952543
transform 1 0 220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6189
timestamp 1682952543
transform 1 0 244 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6247
timestamp 1682952543
transform 1 0 260 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6303
timestamp 1682952543
transform 1 0 236 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1682952543
transform 1 0 252 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1682952543
transform 1 0 260 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6281
timestamp 1682952543
transform 1 0 236 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6314
timestamp 1682952543
transform 1 0 252 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6190
timestamp 1682952543
transform 1 0 276 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6282
timestamp 1682952543
transform 1 0 276 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6213
timestamp 1682952543
transform 1 0 388 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6191
timestamp 1682952543
transform 1 0 308 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6306
timestamp 1682952543
transform 1 0 356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6307
timestamp 1682952543
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6308
timestamp 1682952543
transform 1 0 396 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6283
timestamp 1682952543
transform 1 0 356 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6284
timestamp 1682952543
transform 1 0 396 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6309
timestamp 1682952543
transform 1 0 412 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6315
timestamp 1682952543
transform 1 0 412 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6185
timestamp 1682952543
transform 1 0 420 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6186
timestamp 1682952543
transform 1 0 452 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6214
timestamp 1682952543
transform 1 0 460 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6192
timestamp 1682952543
transform 1 0 436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1682952543
transform 1 0 444 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6194
timestamp 1682952543
transform 1 0 460 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6310
timestamp 1682952543
transform 1 0 452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6311
timestamp 1682952543
transform 1 0 468 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1682952543
transform 1 0 492 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6312
timestamp 1682952543
transform 1 0 484 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6165
timestamp 1682952543
transform 1 0 516 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6187
timestamp 1682952543
transform 1 0 524 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6215
timestamp 1682952543
transform 1 0 540 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6216
timestamp 1682952543
transform 1 0 564 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6196
timestamp 1682952543
transform 1 0 516 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6197
timestamp 1682952543
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1682952543
transform 1 0 540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6199
timestamp 1682952543
transform 1 0 556 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6248
timestamp 1682952543
transform 1 0 564 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6200
timestamp 1682952543
transform 1 0 572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6313
timestamp 1682952543
transform 1 0 508 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1682952543
transform 1 0 524 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6315
timestamp 1682952543
transform 1 0 540 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6285
timestamp 1682952543
transform 1 0 524 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6267
timestamp 1682952543
transform 1 0 556 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6316
timestamp 1682952543
transform 1 0 564 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6286
timestamp 1682952543
transform 1 0 556 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6287
timestamp 1682952543
transform 1 0 572 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6316
timestamp 1682952543
transform 1 0 516 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6317
timestamp 1682952543
transform 1 0 540 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6318
timestamp 1682952543
transform 1 0 556 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6355
timestamp 1682952543
transform 1 0 564 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6378
timestamp 1682952543
transform 1 0 540 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6217
timestamp 1682952543
transform 1 0 588 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6188
timestamp 1682952543
transform 1 0 620 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6201
timestamp 1682952543
transform 1 0 612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6202
timestamp 1682952543
transform 1 0 636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1682952543
transform 1 0 644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1682952543
transform 1 0 604 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6288
timestamp 1682952543
transform 1 0 596 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6319
timestamp 1682952543
transform 1 0 588 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6379
timestamp 1682952543
transform 1 0 588 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6356
timestamp 1682952543
transform 1 0 604 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6318
timestamp 1682952543
transform 1 0 628 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1682952543
transform 1 0 644 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6289
timestamp 1682952543
transform 1 0 636 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6357
timestamp 1682952543
transform 1 0 644 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6204
timestamp 1682952543
transform 1 0 684 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1682952543
transform 1 0 676 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6320
timestamp 1682952543
transform 1 0 692 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6358
timestamp 1682952543
transform 1 0 684 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6321
timestamp 1682952543
transform 1 0 708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1682952543
transform 1 0 724 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6290
timestamp 1682952543
transform 1 0 724 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6380
timestamp 1682952543
transform 1 0 740 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6184
timestamp 1682952543
transform 1 0 756 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6205
timestamp 1682952543
transform 1 0 748 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6268
timestamp 1682952543
transform 1 0 756 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6419
timestamp 1682952543
transform 1 0 756 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6359
timestamp 1682952543
transform 1 0 756 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6218
timestamp 1682952543
transform 1 0 788 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6206
timestamp 1682952543
transform 1 0 772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6207
timestamp 1682952543
transform 1 0 788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1682952543
transform 1 0 788 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6324
timestamp 1682952543
transform 1 0 796 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6291
timestamp 1682952543
transform 1 0 788 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6208
timestamp 1682952543
transform 1 0 820 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6249
timestamp 1682952543
transform 1 0 836 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6209
timestamp 1682952543
transform 1 0 844 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1682952543
transform 1 0 828 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6292
timestamp 1682952543
transform 1 0 820 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6420
timestamp 1682952543
transform 1 0 836 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6321
timestamp 1682952543
transform 1 0 828 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6250
timestamp 1682952543
transform 1 0 860 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6210
timestamp 1682952543
transform 1 0 868 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1682952543
transform 1 0 884 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1682952543
transform 1 0 892 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6166
timestamp 1682952543
transform 1 0 924 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6185
timestamp 1682952543
transform 1 0 924 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1682952543
transform 1 0 860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1682952543
transform 1 0 876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6328
timestamp 1682952543
transform 1 0 900 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1682952543
transform 1 0 916 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6293
timestamp 1682952543
transform 1 0 860 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6322
timestamp 1682952543
transform 1 0 844 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6323
timestamp 1682952543
transform 1 0 884 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6381
timestamp 1682952543
transform 1 0 860 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6219
timestamp 1682952543
transform 1 0 932 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6213
timestamp 1682952543
transform 1 0 940 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1682952543
transform 1 0 932 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1682952543
transform 1 0 964 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1682952543
transform 1 0 964 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6220
timestamp 1682952543
transform 1 0 1060 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6215
timestamp 1682952543
transform 1 0 980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6216
timestamp 1682952543
transform 1 0 1068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6332
timestamp 1682952543
transform 1 0 1012 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1682952543
transform 1 0 1060 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6324
timestamp 1682952543
transform 1 0 972 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6325
timestamp 1682952543
transform 1 0 1020 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6360
timestamp 1682952543
transform 1 0 1060 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6382
timestamp 1682952543
transform 1 0 980 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6383
timestamp 1682952543
transform 1 0 996 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6384
timestamp 1682952543
transform 1 0 1044 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6269
timestamp 1682952543
transform 1 0 1108 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6221
timestamp 1682952543
transform 1 0 1132 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6334
timestamp 1682952543
transform 1 0 1116 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1682952543
transform 1 0 1092 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6326
timestamp 1682952543
transform 1 0 1092 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6270
timestamp 1682952543
transform 1 0 1124 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6422
timestamp 1682952543
transform 1 0 1124 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6327
timestamp 1682952543
transform 1 0 1124 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6217
timestamp 1682952543
transform 1 0 1164 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1682952543
transform 1 0 1156 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6218
timestamp 1682952543
transform 1 0 1172 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6328
timestamp 1682952543
transform 1 0 1164 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6336
timestamp 1682952543
transform 1 0 1188 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6167
timestamp 1682952543
transform 1 0 1204 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6222
timestamp 1682952543
transform 1 0 1220 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6219
timestamp 1682952543
transform 1 0 1244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6337
timestamp 1682952543
transform 1 0 1260 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6385
timestamp 1682952543
transform 1 0 1260 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6168
timestamp 1682952543
transform 1 0 1356 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6189
timestamp 1682952543
transform 1 0 1300 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6190
timestamp 1682952543
transform 1 0 1316 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6220
timestamp 1682952543
transform 1 0 1276 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6251
timestamp 1682952543
transform 1 0 1316 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6338
timestamp 1682952543
transform 1 0 1316 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6386
timestamp 1682952543
transform 1 0 1284 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6387
timestamp 1682952543
transform 1 0 1308 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6221
timestamp 1682952543
transform 1 0 1380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1682952543
transform 1 0 1372 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6329
timestamp 1682952543
transform 1 0 1372 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6388
timestamp 1682952543
transform 1 0 1380 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6169
timestamp 1682952543
transform 1 0 1404 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6252
timestamp 1682952543
transform 1 0 1404 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6222
timestamp 1682952543
transform 1 0 1412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6223
timestamp 1682952543
transform 1 0 1436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1682952543
transform 1 0 1404 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6341
timestamp 1682952543
transform 1 0 1428 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6330
timestamp 1682952543
transform 1 0 1404 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6294
timestamp 1682952543
transform 1 0 1436 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6191
timestamp 1682952543
transform 1 0 1540 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6224
timestamp 1682952543
transform 1 0 1452 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6253
timestamp 1682952543
transform 1 0 1500 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6254
timestamp 1682952543
transform 1 0 1540 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6225
timestamp 1682952543
transform 1 0 1556 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1682952543
transform 1 0 1500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6343
timestamp 1682952543
transform 1 0 1532 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6344
timestamp 1682952543
transform 1 0 1540 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6345
timestamp 1682952543
transform 1 0 1548 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6331
timestamp 1682952543
transform 1 0 1452 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6389
timestamp 1682952543
transform 1 0 1516 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6192
timestamp 1682952543
transform 1 0 1564 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6193
timestamp 1682952543
transform 1 0 1580 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6346
timestamp 1682952543
transform 1 0 1572 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6347
timestamp 1682952543
transform 1 0 1588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1682952543
transform 1 0 1604 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6332
timestamp 1682952543
transform 1 0 1596 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6226
timestamp 1682952543
transform 1 0 1620 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6333
timestamp 1682952543
transform 1 0 1620 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6227
timestamp 1682952543
transform 1 0 1636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6349
timestamp 1682952543
transform 1 0 1636 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6350
timestamp 1682952543
transform 1 0 1652 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6334
timestamp 1682952543
transform 1 0 1676 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6228
timestamp 1682952543
transform 1 0 1692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1682952543
transform 1 0 1700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6423
timestamp 1682952543
transform 1 0 1692 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1682952543
transform 1 0 1724 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1682952543
transform 1 0 1708 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1682952543
transform 1 0 1724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6424
timestamp 1682952543
transform 1 0 1724 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6361
timestamp 1682952543
transform 1 0 1724 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6353
timestamp 1682952543
transform 1 0 1748 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6335
timestamp 1682952543
transform 1 0 1748 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6231
timestamp 1682952543
transform 1 0 1764 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1682952543
transform 1 0 1788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1682952543
transform 1 0 1788 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6362
timestamp 1682952543
transform 1 0 1788 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6233
timestamp 1682952543
transform 1 0 1796 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6255
timestamp 1682952543
transform 1 0 1804 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6256
timestamp 1682952543
transform 1 0 1820 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6194
timestamp 1682952543
transform 1 0 1844 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6354
timestamp 1682952543
transform 1 0 1836 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6363
timestamp 1682952543
transform 1 0 1844 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6195
timestamp 1682952543
transform 1 0 1876 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6234
timestamp 1682952543
transform 1 0 1860 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1682952543
transform 1 0 1868 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6426
timestamp 1682952543
transform 1 0 1868 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1682952543
transform 1 0 1908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6355
timestamp 1682952543
transform 1 0 1892 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6356
timestamp 1682952543
transform 1 0 1900 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6364
timestamp 1682952543
transform 1 0 1868 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6336
timestamp 1682952543
transform 1 0 1900 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6390
timestamp 1682952543
transform 1 0 1900 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6223
timestamp 1682952543
transform 1 0 1924 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6237
timestamp 1682952543
transform 1 0 1924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1682952543
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6239
timestamp 1682952543
transform 1 0 1948 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6224
timestamp 1682952543
transform 1 0 1964 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6357
timestamp 1682952543
transform 1 0 1956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6427
timestamp 1682952543
transform 1 0 1964 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6365
timestamp 1682952543
transform 1 0 1956 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6240
timestamp 1682952543
transform 1 0 1980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6241
timestamp 1682952543
transform 1 0 2004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6358
timestamp 1682952543
transform 1 0 1996 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6196
timestamp 1682952543
transform 1 0 2044 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6242
timestamp 1682952543
transform 1 0 2036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6359
timestamp 1682952543
transform 1 0 2044 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6428
timestamp 1682952543
transform 1 0 2060 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6243
timestamp 1682952543
transform 1 0 2068 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6360
timestamp 1682952543
transform 1 0 2068 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6337
timestamp 1682952543
transform 1 0 2068 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6366
timestamp 1682952543
transform 1 0 2060 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6244
timestamp 1682952543
transform 1 0 2084 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6257
timestamp 1682952543
transform 1 0 2116 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6429
timestamp 1682952543
transform 1 0 2116 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6367
timestamp 1682952543
transform 1 0 2116 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6245
timestamp 1682952543
transform 1 0 2132 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1682952543
transform 1 0 2132 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6362
timestamp 1682952543
transform 1 0 2164 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6338
timestamp 1682952543
transform 1 0 2164 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6368
timestamp 1682952543
transform 1 0 2164 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6246
timestamp 1682952543
transform 1 0 2180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1682952543
transform 1 0 2188 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6295
timestamp 1682952543
transform 1 0 2180 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6363
timestamp 1682952543
transform 1 0 2196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1682952543
transform 1 0 2212 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6339
timestamp 1682952543
transform 1 0 2188 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6340
timestamp 1682952543
transform 1 0 2212 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6248
timestamp 1682952543
transform 1 0 2228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1682952543
transform 1 0 2236 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1682952543
transform 1 0 2228 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6341
timestamp 1682952543
transform 1 0 2228 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6391
timestamp 1682952543
transform 1 0 2228 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6197
timestamp 1682952543
transform 1 0 2252 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6250
timestamp 1682952543
transform 1 0 2276 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6365
timestamp 1682952543
transform 1 0 2260 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1682952543
transform 1 0 2276 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6296
timestamp 1682952543
transform 1 0 2252 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6431
timestamp 1682952543
transform 1 0 2276 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6342
timestamp 1682952543
transform 1 0 2276 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6225
timestamp 1682952543
transform 1 0 2292 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6251
timestamp 1682952543
transform 1 0 2284 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6369
timestamp 1682952543
transform 1 0 2284 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6226
timestamp 1682952543
transform 1 0 2324 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6367
timestamp 1682952543
transform 1 0 2316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6368
timestamp 1682952543
transform 1 0 2332 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6432
timestamp 1682952543
transform 1 0 2332 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6343
timestamp 1682952543
transform 1 0 2332 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6252
timestamp 1682952543
transform 1 0 2340 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6253
timestamp 1682952543
transform 1 0 2348 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6370
timestamp 1682952543
transform 1 0 2364 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6170
timestamp 1682952543
transform 1 0 2396 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6433
timestamp 1682952543
transform 1 0 2388 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6344
timestamp 1682952543
transform 1 0 2388 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6371
timestamp 1682952543
transform 1 0 2388 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6254
timestamp 1682952543
transform 1 0 2412 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1682952543
transform 1 0 2404 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6297
timestamp 1682952543
transform 1 0 2404 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6255
timestamp 1682952543
transform 1 0 2428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6370
timestamp 1682952543
transform 1 0 2436 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6371
timestamp 1682952543
transform 1 0 2452 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1682952543
transform 1 0 2452 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6345
timestamp 1682952543
transform 1 0 2452 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6256
timestamp 1682952543
transform 1 0 2460 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6227
timestamp 1682952543
transform 1 0 2476 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6257
timestamp 1682952543
transform 1 0 2492 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6228
timestamp 1682952543
transform 1 0 2524 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6372
timestamp 1682952543
transform 1 0 2500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6373
timestamp 1682952543
transform 1 0 2516 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6435
timestamp 1682952543
transform 1 0 2516 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6346
timestamp 1682952543
transform 1 0 2516 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6258
timestamp 1682952543
transform 1 0 2540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6259
timestamp 1682952543
transform 1 0 2548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1682952543
transform 1 0 2556 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6298
timestamp 1682952543
transform 1 0 2564 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6436
timestamp 1682952543
transform 1 0 2572 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6347
timestamp 1682952543
transform 1 0 2572 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6260
timestamp 1682952543
transform 1 0 2596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1682952543
transform 1 0 2604 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6375
timestamp 1682952543
transform 1 0 2620 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6299
timestamp 1682952543
transform 1 0 2620 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6437
timestamp 1682952543
transform 1 0 2636 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6262
timestamp 1682952543
transform 1 0 2652 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6171
timestamp 1682952543
transform 1 0 2676 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6271
timestamp 1682952543
transform 1 0 2668 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6441
timestamp 1682952543
transform 1 0 2668 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_6229
timestamp 1682952543
transform 1 0 2692 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6263
timestamp 1682952543
transform 1 0 2692 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6300
timestamp 1682952543
transform 1 0 2700 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6442
timestamp 1682952543
transform 1 0 2700 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_6198
timestamp 1682952543
transform 1 0 2740 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6230
timestamp 1682952543
transform 1 0 2748 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6264
timestamp 1682952543
transform 1 0 2748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6376
timestamp 1682952543
transform 1 0 2724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1682952543
transform 1 0 2740 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1682952543
transform 1 0 2716 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6372
timestamp 1682952543
transform 1 0 2716 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6172
timestamp 1682952543
transform 1 0 2788 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6199
timestamp 1682952543
transform 1 0 2820 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6265
timestamp 1682952543
transform 1 0 2796 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6266
timestamp 1682952543
transform 1 0 2812 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1682952543
transform 1 0 2820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6378
timestamp 1682952543
transform 1 0 2764 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6379
timestamp 1682952543
transform 1 0 2780 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1682952543
transform 1 0 2788 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6272
timestamp 1682952543
transform 1 0 2796 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6381
timestamp 1682952543
transform 1 0 2804 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1682952543
transform 1 0 2820 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6301
timestamp 1682952543
transform 1 0 2820 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6200
timestamp 1682952543
transform 1 0 2844 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6201
timestamp 1682952543
transform 1 0 2868 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6231
timestamp 1682952543
transform 1 0 2868 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6268
timestamp 1682952543
transform 1 0 2868 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6269
timestamp 1682952543
transform 1 0 2884 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6273
timestamp 1682952543
transform 1 0 2852 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6383
timestamp 1682952543
transform 1 0 2860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1682952543
transform 1 0 2884 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6348
timestamp 1682952543
transform 1 0 2860 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6392
timestamp 1682952543
transform 1 0 2852 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6393
timestamp 1682952543
transform 1 0 2892 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6173
timestamp 1682952543
transform 1 0 2980 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6232
timestamp 1682952543
transform 1 0 2940 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6270
timestamp 1682952543
transform 1 0 2916 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6274
timestamp 1682952543
transform 1 0 2916 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6385
timestamp 1682952543
transform 1 0 2940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1682952543
transform 1 0 3020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6439
timestamp 1682952543
transform 1 0 3028 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6349
timestamp 1682952543
transform 1 0 3020 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6373
timestamp 1682952543
transform 1 0 3028 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6258
timestamp 1682952543
transform 1 0 3044 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6302
timestamp 1682952543
transform 1 0 3060 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6443
timestamp 1682952543
transform 1 0 3052 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_6271
timestamp 1682952543
transform 1 0 3076 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6233
timestamp 1682952543
transform 1 0 3092 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6440
timestamp 1682952543
transform 1 0 3076 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6303
timestamp 1682952543
transform 1 0 3084 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6272
timestamp 1682952543
transform 1 0 3100 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1682952543
transform 1 0 3092 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_6174
timestamp 1682952543
transform 1 0 3188 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6202
timestamp 1682952543
transform 1 0 3180 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6234
timestamp 1682952543
transform 1 0 3156 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6235
timestamp 1682952543
transform 1 0 3204 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6273
timestamp 1682952543
transform 1 0 3140 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1682952543
transform 1 0 3148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6275
timestamp 1682952543
transform 1 0 3156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6276
timestamp 1682952543
transform 1 0 3180 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1682952543
transform 1 0 3188 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1682952543
transform 1 0 3204 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1682952543
transform 1 0 3124 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6275
timestamp 1682952543
transform 1 0 3140 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6279
timestamp 1682952543
transform 1 0 3228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1682952543
transform 1 0 3148 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6389
timestamp 1682952543
transform 1 0 3164 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6390
timestamp 1682952543
transform 1 0 3180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1682952543
transform 1 0 3196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6392
timestamp 1682952543
transform 1 0 3212 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6304
timestamp 1682952543
transform 1 0 3124 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6305
timestamp 1682952543
transform 1 0 3156 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6276
timestamp 1682952543
transform 1 0 3220 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6306
timestamp 1682952543
transform 1 0 3196 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6374
timestamp 1682952543
transform 1 0 3180 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6175
timestamp 1682952543
transform 1 0 3252 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6176
timestamp 1682952543
transform 1 0 3308 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6177
timestamp 1682952543
transform 1 0 3324 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6259
timestamp 1682952543
transform 1 0 3244 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6393
timestamp 1682952543
transform 1 0 3244 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6203
timestamp 1682952543
transform 1 0 3316 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6236
timestamp 1682952543
transform 1 0 3284 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6260
timestamp 1682952543
transform 1 0 3292 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6280
timestamp 1682952543
transform 1 0 3332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6394
timestamp 1682952543
transform 1 0 3284 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6277
timestamp 1682952543
transform 1 0 3332 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6350
timestamp 1682952543
transform 1 0 3300 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6394
timestamp 1682952543
transform 1 0 3332 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6281
timestamp 1682952543
transform 1 0 3364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1682952543
transform 1 0 3396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6395
timestamp 1682952543
transform 1 0 3356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1682952543
transform 1 0 3372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6397
timestamp 1682952543
transform 1 0 3388 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6307
timestamp 1682952543
transform 1 0 3356 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6395
timestamp 1682952543
transform 1 0 3380 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6308
timestamp 1682952543
transform 1 0 3404 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6398
timestamp 1682952543
transform 1 0 3420 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6204
timestamp 1682952543
transform 1 0 3436 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6278
timestamp 1682952543
transform 1 0 3436 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6178
timestamp 1682952543
transform 1 0 3468 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6283
timestamp 1682952543
transform 1 0 3460 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6284
timestamp 1682952543
transform 1 0 3468 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1682952543
transform 1 0 3468 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6351
timestamp 1682952543
transform 1 0 3468 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6375
timestamp 1682952543
transform 1 0 3460 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6396
timestamp 1682952543
transform 1 0 3476 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6261
timestamp 1682952543
transform 1 0 3492 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6205
timestamp 1682952543
transform 1 0 3524 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6206
timestamp 1682952543
transform 1 0 3548 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6237
timestamp 1682952543
transform 1 0 3540 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6285
timestamp 1682952543
transform 1 0 3540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6400
timestamp 1682952543
transform 1 0 3548 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6397
timestamp 1682952543
transform 1 0 3556 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6286
timestamp 1682952543
transform 1 0 3564 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6179
timestamp 1682952543
transform 1 0 3588 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6238
timestamp 1682952543
transform 1 0 3612 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6287
timestamp 1682952543
transform 1 0 3596 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6262
timestamp 1682952543
transform 1 0 3604 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6288
timestamp 1682952543
transform 1 0 3612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6401
timestamp 1682952543
transform 1 0 3588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6402
timestamp 1682952543
transform 1 0 3604 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6263
timestamp 1682952543
transform 1 0 3628 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6403
timestamp 1682952543
transform 1 0 3628 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6180
timestamp 1682952543
transform 1 0 3644 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6404
timestamp 1682952543
transform 1 0 3644 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6289
timestamp 1682952543
transform 1 0 3660 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6239
timestamp 1682952543
transform 1 0 3692 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6290
timestamp 1682952543
transform 1 0 3692 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1682952543
transform 1 0 3716 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1682952543
transform 1 0 3700 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6406
timestamp 1682952543
transform 1 0 3716 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6181
timestamp 1682952543
transform 1 0 3796 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6182
timestamp 1682952543
transform 1 0 3820 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6207
timestamp 1682952543
transform 1 0 3780 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6208
timestamp 1682952543
transform 1 0 3804 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6240
timestamp 1682952543
transform 1 0 3772 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6241
timestamp 1682952543
transform 1 0 3820 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6292
timestamp 1682952543
transform 1 0 3820 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1682952543
transform 1 0 3740 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6408
timestamp 1682952543
transform 1 0 3772 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6279
timestamp 1682952543
transform 1 0 3796 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6280
timestamp 1682952543
transform 1 0 3820 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6309
timestamp 1682952543
transform 1 0 3796 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6409
timestamp 1682952543
transform 1 0 3836 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6310
timestamp 1682952543
transform 1 0 3836 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6352
timestamp 1682952543
transform 1 0 3828 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6242
timestamp 1682952543
transform 1 0 3852 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6243
timestamp 1682952543
transform 1 0 3924 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6183
timestamp 1682952543
transform 1 0 3948 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6209
timestamp 1682952543
transform 1 0 3948 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6264
timestamp 1682952543
transform 1 0 3884 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6293
timestamp 1682952543
transform 1 0 3924 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6265
timestamp 1682952543
transform 1 0 3940 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6294
timestamp 1682952543
transform 1 0 3948 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6266
timestamp 1682952543
transform 1 0 3972 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6295
timestamp 1682952543
transform 1 0 3980 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6410
timestamp 1682952543
transform 1 0 3876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6411
timestamp 1682952543
transform 1 0 3940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1682952543
transform 1 0 3956 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6413
timestamp 1682952543
transform 1 0 3972 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6353
timestamp 1682952543
transform 1 0 3876 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6376
timestamp 1682952543
transform 1 0 3844 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6377
timestamp 1682952543
transform 1 0 3956 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6210
timestamp 1682952543
transform 1 0 3996 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_6244
timestamp 1682952543
transform 1 0 4004 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6184
timestamp 1682952543
transform 1 0 4108 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_6245
timestamp 1682952543
transform 1 0 4060 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6296
timestamp 1682952543
transform 1 0 4004 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6297
timestamp 1682952543
transform 1 0 4020 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6298
timestamp 1682952543
transform 1 0 4036 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6414
timestamp 1682952543
transform 1 0 3988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1682952543
transform 1 0 3996 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6416
timestamp 1682952543
transform 1 0 4012 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6311
timestamp 1682952543
transform 1 0 3988 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6312
timestamp 1682952543
transform 1 0 4012 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6417
timestamp 1682952543
transform 1 0 4060 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6354
timestamp 1682952543
transform 1 0 4076 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6418
timestamp 1682952543
transform 1 0 4132 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6313
timestamp 1682952543
transform 1 0 4132 0 1 1515
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_52
timestamp 1682952543
transform 1 0 24 0 1 1470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_374
timestamp 1682952543
transform 1 0 72 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_420
timestamp 1682952543
transform -1 0 184 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2446
timestamp 1682952543
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1682952543
transform 1 0 192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1682952543
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1682952543
transform 1 0 208 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_248
timestamp 1682952543
transform -1 0 256 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2450
timestamp 1682952543
transform 1 0 256 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_421
timestamp 1682952543
transform -1 0 280 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2451
timestamp 1682952543
transform 1 0 280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1682952543
transform 1 0 288 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_377
timestamp 1682952543
transform 1 0 296 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_422
timestamp 1682952543
transform -1 0 408 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2453
timestamp 1682952543
transform 1 0 408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1682952543
transform 1 0 416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1682952543
transform 1 0 424 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_249
timestamp 1682952543
transform 1 0 432 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2456
timestamp 1682952543
transform 1 0 472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1682952543
transform 1 0 480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2458
timestamp 1682952543
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_263
timestamp 1682952543
transform 1 0 496 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_264
timestamp 1682952543
transform 1 0 536 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2459
timestamp 1682952543
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6398
timestamp 1682952543
transform 1 0 604 0 1 1475
box -3 -3 3 3
use FILL  FILL_2460
timestamp 1682952543
transform 1 0 584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1682952543
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2462
timestamp 1682952543
transform 1 0 600 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_250
timestamp 1682952543
transform 1 0 608 0 -1 1570
box -8 -3 46 105
use INVX2  INVX2_423
timestamp 1682952543
transform 1 0 648 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2463
timestamp 1682952543
transform 1 0 664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1682952543
transform 1 0 672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1682952543
transform 1 0 680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2466
timestamp 1682952543
transform 1 0 688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1682952543
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1682952543
transform 1 0 704 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_88
timestamp 1682952543
transform 1 0 712 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2473
timestamp 1682952543
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1682952543
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_79
timestamp 1682952543
transform 1 0 760 0 -1 1570
box -8 -3 32 105
use OAI21X1  OAI21X1_89
timestamp 1682952543
transform 1 0 784 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2480
timestamp 1682952543
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2481
timestamp 1682952543
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1682952543
transform 1 0 832 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_253
timestamp 1682952543
transform 1 0 840 0 -1 1570
box -8 -3 46 105
use AOI22X1  AOI22X1_254
timestamp 1682952543
transform 1 0 880 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2490
timestamp 1682952543
transform 1 0 920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1682952543
transform 1 0 928 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_81
timestamp 1682952543
transform 1 0 936 0 -1 1570
box -8 -3 32 105
use FILL  FILL_2504
timestamp 1682952543
transform 1 0 960 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_378
timestamp 1682952543
transform 1 0 968 0 -1 1570
box -8 -3 104 105
use FILL  FILL_2505
timestamp 1682952543
transform 1 0 1064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1682952543
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1682952543
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_90
timestamp 1682952543
transform -1 0 1120 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2513
timestamp 1682952543
transform 1 0 1120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2515
timestamp 1682952543
transform 1 0 1128 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1682952543
transform 1 0 1136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1682952543
transform 1 0 1144 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2524
timestamp 1682952543
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1682952543
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_92
timestamp 1682952543
transform -1 0 1200 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2526
timestamp 1682952543
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1682952543
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_426
timestamp 1682952543
transform -1 0 1232 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2528
timestamp 1682952543
transform 1 0 1232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1682952543
transform 1 0 1240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2532
timestamp 1682952543
transform 1 0 1248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1682952543
transform 1 0 1256 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_381
timestamp 1682952543
transform 1 0 1264 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_427
timestamp 1682952543
transform 1 0 1360 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2548
timestamp 1682952543
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2549
timestamp 1682952543
transform 1 0 1384 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_266
timestamp 1682952543
transform -1 0 1432 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2550
timestamp 1682952543
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_382
timestamp 1682952543
transform 1 0 1440 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_428
timestamp 1682952543
transform -1 0 1552 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2551
timestamp 1682952543
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1682952543
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6399
timestamp 1682952543
transform 1 0 1612 0 1 1475
box -3 -3 3 3
use AOI22X1  AOI22X1_257
timestamp 1682952543
transform 1 0 1568 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2553
timestamp 1682952543
transform 1 0 1608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1682952543
transform 1 0 1616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2555
timestamp 1682952543
transform 1 0 1624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1682952543
transform 1 0 1632 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_93
timestamp 1682952543
transform 1 0 1640 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2557
timestamp 1682952543
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2559
timestamp 1682952543
transform 1 0 1680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1682952543
transform 1 0 1688 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_94
timestamp 1682952543
transform 1 0 1696 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2564
timestamp 1682952543
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2566
timestamp 1682952543
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2577
timestamp 1682952543
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1682952543
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_97
timestamp 1682952543
transform 1 0 1760 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2579
timestamp 1682952543
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1682952543
transform 1 0 1800 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_87
timestamp 1682952543
transform -1 0 1832 0 -1 1570
box -5 -3 28 105
use FILL  FILL_2581
timestamp 1682952543
transform 1 0 1832 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_88
timestamp 1682952543
transform 1 0 1840 0 -1 1570
box -5 -3 28 105
use FILL  FILL_2582
timestamp 1682952543
transform 1 0 1864 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6400
timestamp 1682952543
transform 1 0 1892 0 1 1475
box -3 -3 3 3
use OAI21X1  OAI21X1_98
timestamp 1682952543
transform -1 0 1904 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2583
timestamp 1682952543
transform 1 0 1904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1682952543
transform 1 0 1912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1682952543
transform 1 0 1920 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_430
timestamp 1682952543
transform 1 0 1928 0 -1 1570
box -9 -3 26 105
use NAND2X1  NAND2X1_62
timestamp 1682952543
transform 1 0 1944 0 -1 1570
box -8 -3 32 105
use FILL  FILL_2586
timestamp 1682952543
transform 1 0 1968 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6401
timestamp 1682952543
transform 1 0 1996 0 1 1475
box -3 -3 3 3
use OAI21X1  OAI21X1_99
timestamp 1682952543
transform -1 0 2008 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2587
timestamp 1682952543
transform 1 0 2008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1682952543
transform 1 0 2016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2589
timestamp 1682952543
transform 1 0 2024 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_100
timestamp 1682952543
transform 1 0 2032 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2590
timestamp 1682952543
transform 1 0 2064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1682952543
transform 1 0 2072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1682952543
transform 1 0 2080 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6402
timestamp 1682952543
transform 1 0 2108 0 1 1475
box -3 -3 3 3
use OAI21X1  OAI21X1_101
timestamp 1682952543
transform 1 0 2088 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2596
timestamp 1682952543
transform 1 0 2120 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1682952543
transform 1 0 2128 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_89
timestamp 1682952543
transform 1 0 2136 0 -1 1570
box -5 -3 28 105
use FILL  FILL_2603
timestamp 1682952543
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6403
timestamp 1682952543
transform 1 0 2188 0 1 1475
box -3 -3 3 3
use FILL  FILL_2604
timestamp 1682952543
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1682952543
transform 1 0 2176 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_103
timestamp 1682952543
transform 1 0 2184 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2606
timestamp 1682952543
transform 1 0 2216 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1682952543
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1682952543
transform 1 0 2232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1682952543
transform 1 0 2240 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_104
timestamp 1682952543
transform 1 0 2248 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2610
timestamp 1682952543
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2611
timestamp 1682952543
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1682952543
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_105
timestamp 1682952543
transform 1 0 2304 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2613
timestamp 1682952543
transform 1 0 2336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1682952543
transform 1 0 2344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1682952543
transform 1 0 2352 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_106
timestamp 1682952543
transform 1 0 2360 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2616
timestamp 1682952543
transform 1 0 2392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1682952543
transform 1 0 2400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2618
timestamp 1682952543
transform 1 0 2408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1682952543
transform 1 0 2416 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_108
timestamp 1682952543
transform 1 0 2424 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2622
timestamp 1682952543
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1682952543
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1682952543
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1682952543
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_109
timestamp 1682952543
transform 1 0 2488 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2630
timestamp 1682952543
transform 1 0 2520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1682952543
transform 1 0 2528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1682952543
transform 1 0 2536 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_110
timestamp 1682952543
transform 1 0 2544 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2643
timestamp 1682952543
transform 1 0 2576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1682952543
transform 1 0 2584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1682952543
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_111
timestamp 1682952543
transform -1 0 2632 0 -1 1570
box -8 -3 34 105
use FILL  FILL_2646
timestamp 1682952543
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2647
timestamp 1682952543
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1682952543
transform 1 0 2648 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_57
timestamp 1682952543
transform -1 0 2688 0 -1 1570
box -8 -3 40 105
use FILL  FILL_2649
timestamp 1682952543
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1682952543
transform 1 0 2696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1682952543
transform 1 0 2704 0 -1 1570
box -8 -3 16 105
use AND2X2  AND2X2_49
timestamp 1682952543
transform 1 0 2712 0 -1 1570
box -8 -3 40 105
use FILL  FILL_2656
timestamp 1682952543
transform 1 0 2744 0 -1 1570
box -8 -3 16 105
use AND2X2  AND2X2_50
timestamp 1682952543
transform 1 0 2752 0 -1 1570
box -8 -3 40 105
use AOI22X1  AOI22X1_261
timestamp 1682952543
transform 1 0 2784 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2657
timestamp 1682952543
transform 1 0 2824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1682952543
transform 1 0 2832 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2663
timestamp 1682952543
transform 1 0 2840 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_267
timestamp 1682952543
transform -1 0 2888 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2664
timestamp 1682952543
transform 1 0 2888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1682952543
transform 1 0 2896 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_389
timestamp 1682952543
transform 1 0 2904 0 -1 1570
box -8 -3 104 105
use FILL  FILL_2686
timestamp 1682952543
transform 1 0 3000 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_435
timestamp 1682952543
transform 1 0 3008 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2687
timestamp 1682952543
transform 1 0 3024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2688
timestamp 1682952543
transform 1 0 3032 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_60
timestamp 1682952543
transform -1 0 3072 0 -1 1570
box -8 -3 40 105
use FILL  FILL_2689
timestamp 1682952543
transform 1 0 3072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1682952543
transform 1 0 3080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1682952543
transform 1 0 3088 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_90
timestamp 1682952543
transform -1 0 3120 0 -1 1570
box -5 -3 28 105
use M3_M2  M3_M2_6404
timestamp 1682952543
transform 1 0 3148 0 1 1475
box -3 -3 3 3
use BUFX2  BUFX2_91
timestamp 1682952543
transform 1 0 3120 0 -1 1570
box -5 -3 28 105
use AOI22X1  AOI22X1_264
timestamp 1682952543
transform -1 0 3184 0 -1 1570
box -8 -3 46 105
use OAI22X1  OAI22X1_270
timestamp 1682952543
transform -1 0 3224 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2692
timestamp 1682952543
transform 1 0 3224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1682952543
transform 1 0 3232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1682952543
transform 1 0 3240 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_390
timestamp 1682952543
transform -1 0 3344 0 -1 1570
box -8 -3 104 105
use FILL  FILL_2695
timestamp 1682952543
transform 1 0 3344 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6405
timestamp 1682952543
transform 1 0 3388 0 1 1475
box -3 -3 3 3
use AOI22X1  AOI22X1_265
timestamp 1682952543
transform 1 0 3352 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2696
timestamp 1682952543
transform 1 0 3392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1682952543
transform 1 0 3400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1682952543
transform 1 0 3408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1682952543
transform 1 0 3416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1682952543
transform 1 0 3424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1682952543
transform 1 0 3432 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_92
timestamp 1682952543
transform 1 0 3440 0 -1 1570
box -5 -3 28 105
use FILL  FILL_2702
timestamp 1682952543
transform 1 0 3464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1682952543
transform 1 0 3472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2706
timestamp 1682952543
transform 1 0 3480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1682952543
transform 1 0 3488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2708
timestamp 1682952543
transform 1 0 3496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1682952543
transform 1 0 3504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1682952543
transform 1 0 3512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1682952543
transform 1 0 3520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1682952543
transform 1 0 3528 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_436
timestamp 1682952543
transform 1 0 3536 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2717
timestamp 1682952543
transform 1 0 3552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1682952543
transform 1 0 3560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1682952543
transform 1 0 3568 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_271
timestamp 1682952543
transform 1 0 3576 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2728
timestamp 1682952543
transform 1 0 3616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1682952543
transform 1 0 3624 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6406
timestamp 1682952543
transform 1 0 3644 0 1 1475
box -3 -3 3 3
use INVX2  INVX2_437
timestamp 1682952543
transform -1 0 3648 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2730
timestamp 1682952543
transform 1 0 3648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1682952543
transform 1 0 3656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2734
timestamp 1682952543
transform 1 0 3664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1682952543
transform 1 0 3672 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_268
timestamp 1682952543
transform -1 0 3720 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2751
timestamp 1682952543
transform 1 0 3720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2752
timestamp 1682952543
transform 1 0 3728 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6407
timestamp 1682952543
transform 1 0 3764 0 1 1475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_393
timestamp 1682952543
transform -1 0 3832 0 -1 1570
box -8 -3 104 105
use FILL  FILL_2753
timestamp 1682952543
transform 1 0 3832 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6408
timestamp 1682952543
transform 1 0 3916 0 1 1475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_394
timestamp 1682952543
transform -1 0 3936 0 -1 1570
box -8 -3 104 105
use AOI22X1  AOI22X1_269
timestamp 1682952543
transform 1 0 3936 0 -1 1570
box -8 -3 46 105
use FILL  FILL_2754
timestamp 1682952543
transform 1 0 3976 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_274
timestamp 1682952543
transform 1 0 3984 0 -1 1570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_395
timestamp 1682952543
transform 1 0 4024 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_441
timestamp 1682952543
transform 1 0 4120 0 -1 1570
box -9 -3 26 105
use FILL  FILL_2755
timestamp 1682952543
transform 1 0 4136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1682952543
transform 1 0 4144 0 -1 1570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_53
timestamp 1682952543
transform 1 0 4201 0 1 1470
box -10 -3 10 3
use M3_M2  M3_M2_6489
timestamp 1682952543
transform 1 0 132 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6490
timestamp 1682952543
transform 1 0 164 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6453
timestamp 1682952543
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1682952543
transform 1 0 84 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6454
timestamp 1682952543
transform 1 0 196 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6456
timestamp 1682952543
transform 1 0 212 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6455
timestamp 1682952543
transform 1 0 220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1682952543
transform 1 0 212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1682952543
transform 1 0 236 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6456
timestamp 1682952543
transform 1 0 252 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6556
timestamp 1682952543
transform 1 0 252 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6491
timestamp 1682952543
transform 1 0 316 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6492
timestamp 1682952543
transform 1 0 356 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6531
timestamp 1682952543
transform 1 0 268 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6532
timestamp 1682952543
transform 1 0 308 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6457
timestamp 1682952543
transform 1 0 316 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6458
timestamp 1682952543
transform 1 0 348 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1682952543
transform 1 0 356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6460
timestamp 1682952543
transform 1 0 364 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1682952543
transform 1 0 268 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6557
timestamp 1682952543
transform 1 0 364 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6575
timestamp 1682952543
transform 1 0 348 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6533
timestamp 1682952543
transform 1 0 388 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6409
timestamp 1682952543
transform 1 0 412 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6436
timestamp 1682952543
transform 1 0 420 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6437
timestamp 1682952543
transform 1 0 436 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6461
timestamp 1682952543
transform 1 0 396 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6534
timestamp 1682952543
transform 1 0 404 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6462
timestamp 1682952543
transform 1 0 412 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6535
timestamp 1682952543
transform 1 0 428 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6563
timestamp 1682952543
transform 1 0 396 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1682952543
transform 1 0 404 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6565
timestamp 1682952543
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6576
timestamp 1682952543
transform 1 0 420 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6621
timestamp 1682952543
transform 1 0 420 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6463
timestamp 1682952543
transform 1 0 444 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6438
timestamp 1682952543
transform 1 0 476 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6439
timestamp 1682952543
transform 1 0 500 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6457
timestamp 1682952543
transform 1 0 532 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6493
timestamp 1682952543
transform 1 0 460 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6464
timestamp 1682952543
transform 1 0 484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6465
timestamp 1682952543
transform 1 0 540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1682952543
transform 1 0 460 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6577
timestamp 1682952543
transform 1 0 492 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6622
timestamp 1682952543
transform 1 0 460 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6494
timestamp 1682952543
transform 1 0 564 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6410
timestamp 1682952543
transform 1 0 596 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6495
timestamp 1682952543
transform 1 0 588 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6466
timestamp 1682952543
transform 1 0 588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6467
timestamp 1682952543
transform 1 0 604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1682952543
transform 1 0 596 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6623
timestamp 1682952543
transform 1 0 596 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6568
timestamp 1682952543
transform 1 0 628 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6578
timestamp 1682952543
transform 1 0 620 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6411
timestamp 1682952543
transform 1 0 708 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6412
timestamp 1682952543
transform 1 0 740 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6413
timestamp 1682952543
transform 1 0 756 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6496
timestamp 1682952543
transform 1 0 684 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6497
timestamp 1682952543
transform 1 0 732 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6536
timestamp 1682952543
transform 1 0 652 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6468
timestamp 1682952543
transform 1 0 676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6469
timestamp 1682952543
transform 1 0 732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6470
timestamp 1682952543
transform 1 0 740 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6471
timestamp 1682952543
transform 1 0 748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6569
timestamp 1682952543
transform 1 0 652 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6558
timestamp 1682952543
transform 1 0 676 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6570
timestamp 1682952543
transform 1 0 740 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6579
timestamp 1682952543
transform 1 0 652 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6580
timestamp 1682952543
transform 1 0 668 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6581
timestamp 1682952543
transform 1 0 716 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6571
timestamp 1682952543
transform 1 0 772 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6414
timestamp 1682952543
transform 1 0 796 0 1 1465
box -3 -3 3 3
use M2_M1  M2_M1_6446
timestamp 1682952543
transform 1 0 796 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6559
timestamp 1682952543
transform 1 0 796 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6572
timestamp 1682952543
transform 1 0 804 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6658
timestamp 1682952543
transform 1 0 788 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6624
timestamp 1682952543
transform 1 0 788 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6582
timestamp 1682952543
transform 1 0 804 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6458
timestamp 1682952543
transform 1 0 820 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6415
timestamp 1682952543
transform 1 0 844 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6440
timestamp 1682952543
transform 1 0 836 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6472
timestamp 1682952543
transform 1 0 828 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6416
timestamp 1682952543
transform 1 0 876 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6459
timestamp 1682952543
transform 1 0 852 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6460
timestamp 1682952543
transform 1 0 940 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6498
timestamp 1682952543
transform 1 0 908 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6537
timestamp 1682952543
transform 1 0 900 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6499
timestamp 1682952543
transform 1 0 948 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6473
timestamp 1682952543
transform 1 0 908 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6474
timestamp 1682952543
transform 1 0 940 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6475
timestamp 1682952543
transform 1 0 948 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1682952543
transform 1 0 860 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6625
timestamp 1682952543
transform 1 0 924 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6417
timestamp 1682952543
transform 1 0 956 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6538
timestamp 1682952543
transform 1 0 956 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6574
timestamp 1682952543
transform 1 0 956 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6583
timestamp 1682952543
transform 1 0 964 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6626
timestamp 1682952543
transform 1 0 956 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6418
timestamp 1682952543
transform 1 0 988 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6461
timestamp 1682952543
transform 1 0 980 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6575
timestamp 1682952543
transform 1 0 980 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6419
timestamp 1682952543
transform 1 0 1012 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6420
timestamp 1682952543
transform 1 0 1052 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6462
timestamp 1682952543
transform 1 0 1044 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6500
timestamp 1682952543
transform 1 0 1020 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6447
timestamp 1682952543
transform 1 0 1044 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1682952543
transform 1 0 1020 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6477
timestamp 1682952543
transform 1 0 1036 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6539
timestamp 1682952543
transform 1 0 1044 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6478
timestamp 1682952543
transform 1 0 1060 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6540
timestamp 1682952543
transform 1 0 1068 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6576
timestamp 1682952543
transform 1 0 1036 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1682952543
transform 1 0 1044 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6560
timestamp 1682952543
transform 1 0 1052 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6578
timestamp 1682952543
transform 1 0 1068 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6584
timestamp 1682952543
transform 1 0 1036 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6441
timestamp 1682952543
transform 1 0 1084 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6463
timestamp 1682952543
transform 1 0 1092 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6448
timestamp 1682952543
transform 1 0 1092 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1682952543
transform 1 0 1084 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6421
timestamp 1682952543
transform 1 0 1124 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6501
timestamp 1682952543
transform 1 0 1124 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6479
timestamp 1682952543
transform 1 0 1132 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6464
timestamp 1682952543
transform 1 0 1148 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6541
timestamp 1682952543
transform 1 0 1148 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6580
timestamp 1682952543
transform 1 0 1148 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6465
timestamp 1682952543
transform 1 0 1188 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6480
timestamp 1682952543
transform 1 0 1212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1682952543
transform 1 0 1244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1682952543
transform 1 0 1164 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6585
timestamp 1682952543
transform 1 0 1212 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6627
timestamp 1682952543
transform 1 0 1164 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6628
timestamp 1682952543
transform 1 0 1260 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6482
timestamp 1682952543
transform 1 0 1284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1682952543
transform 1 0 1324 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1682952543
transform 1 0 1276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1682952543
transform 1 0 1292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1682952543
transform 1 0 1308 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1682952543
transform 1 0 1316 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6586
timestamp 1682952543
transform 1 0 1292 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6629
timestamp 1682952543
transform 1 0 1276 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6630
timestamp 1682952543
transform 1 0 1316 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6484
timestamp 1682952543
transform 1 0 1348 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6561
timestamp 1682952543
transform 1 0 1348 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6502
timestamp 1682952543
transform 1 0 1372 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6485
timestamp 1682952543
transform 1 0 1372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6486
timestamp 1682952543
transform 1 0 1388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1682952543
transform 1 0 1380 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6562
timestamp 1682952543
transform 1 0 1388 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6587
timestamp 1682952543
transform 1 0 1380 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6487
timestamp 1682952543
transform 1 0 1428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1682952543
transform 1 0 1428 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6631
timestamp 1682952543
transform 1 0 1428 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6488
timestamp 1682952543
transform 1 0 1468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1682952543
transform 1 0 1444 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6588
timestamp 1682952543
transform 1 0 1468 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6632
timestamp 1682952543
transform 1 0 1508 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6428
timestamp 1682952543
transform 1 0 1540 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6429
timestamp 1682952543
transform 1 0 1564 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6442
timestamp 1682952543
transform 1 0 1556 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6466
timestamp 1682952543
transform 1 0 1564 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6503
timestamp 1682952543
transform 1 0 1548 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6489
timestamp 1682952543
transform 1 0 1548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1682952543
transform 1 0 1564 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6422
timestamp 1682952543
transform 1 0 1636 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6430
timestamp 1682952543
transform 1 0 1636 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6431
timestamp 1682952543
transform 1 0 1668 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6467
timestamp 1682952543
transform 1 0 1588 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6504
timestamp 1682952543
transform 1 0 1580 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6490
timestamp 1682952543
transform 1 0 1580 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6443
timestamp 1682952543
transform 1 0 1684 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6505
timestamp 1682952543
transform 1 0 1620 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6506
timestamp 1682952543
transform 1 0 1676 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6491
timestamp 1682952543
transform 1 0 1620 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6542
timestamp 1682952543
transform 1 0 1668 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6492
timestamp 1682952543
transform 1 0 1676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6590
timestamp 1682952543
transform 1 0 1596 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1682952543
transform 1 0 1684 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1682952543
transform 1 0 1708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1682952543
transform 1 0 1724 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1682952543
transform 1 0 1724 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6589
timestamp 1682952543
transform 1 0 1724 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6494
timestamp 1682952543
transform 1 0 1748 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6444
timestamp 1682952543
transform 1 0 1772 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6507
timestamp 1682952543
transform 1 0 1764 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6593
timestamp 1682952543
transform 1 0 1756 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1682952543
transform 1 0 1764 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6590
timestamp 1682952543
transform 1 0 1740 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6591
timestamp 1682952543
transform 1 0 1756 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6495
timestamp 1682952543
transform 1 0 1796 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1682952543
transform 1 0 1812 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6592
timestamp 1682952543
transform 1 0 1812 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6593
timestamp 1682952543
transform 1 0 1828 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6450
timestamp 1682952543
transform 1 0 1844 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6633
timestamp 1682952543
transform 1 0 1836 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6508
timestamp 1682952543
transform 1 0 1876 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6496
timestamp 1682952543
transform 1 0 1876 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1682952543
transform 1 0 1868 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6597
timestamp 1682952543
transform 1 0 1876 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6594
timestamp 1682952543
transform 1 0 1876 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6509
timestamp 1682952543
transform 1 0 1892 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6497
timestamp 1682952543
transform 1 0 1884 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6563
timestamp 1682952543
transform 1 0 1884 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6598
timestamp 1682952543
transform 1 0 1892 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6634
timestamp 1682952543
transform 1 0 1892 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6510
timestamp 1682952543
transform 1 0 1916 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6498
timestamp 1682952543
transform 1 0 1900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1682952543
transform 1 0 1924 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1682952543
transform 1 0 1988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1682952543
transform 1 0 1916 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6600
timestamp 1682952543
transform 1 0 1940 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6564
timestamp 1682952543
transform 1 0 1980 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6595
timestamp 1682952543
transform 1 0 1988 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6501
timestamp 1682952543
transform 1 0 2036 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6543
timestamp 1682952543
transform 1 0 2052 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6502
timestamp 1682952543
transform 1 0 2092 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6601
timestamp 1682952543
transform 1 0 2052 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6565
timestamp 1682952543
transform 1 0 2092 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6566
timestamp 1682952543
transform 1 0 2140 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6596
timestamp 1682952543
transform 1 0 2068 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6635
timestamp 1682952543
transform 1 0 2044 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6423
timestamp 1682952543
transform 1 0 2180 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6511
timestamp 1682952543
transform 1 0 2172 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6503
timestamp 1682952543
transform 1 0 2164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1682952543
transform 1 0 2172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6602
timestamp 1682952543
transform 1 0 2180 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6512
timestamp 1682952543
transform 1 0 2196 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6513
timestamp 1682952543
transform 1 0 2212 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6505
timestamp 1682952543
transform 1 0 2212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6603
timestamp 1682952543
transform 1 0 2204 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6597
timestamp 1682952543
transform 1 0 2204 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6604
timestamp 1682952543
transform 1 0 2228 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6567
timestamp 1682952543
transform 1 0 2244 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6468
timestamp 1682952543
transform 1 0 2260 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6506
timestamp 1682952543
transform 1 0 2284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1682952543
transform 1 0 2260 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6598
timestamp 1682952543
transform 1 0 2284 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6469
timestamp 1682952543
transform 1 0 2372 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6514
timestamp 1682952543
transform 1 0 2356 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6507
timestamp 1682952543
transform 1 0 2356 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6606
timestamp 1682952543
transform 1 0 2364 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6599
timestamp 1682952543
transform 1 0 2364 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6508
timestamp 1682952543
transform 1 0 2372 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6432
timestamp 1682952543
transform 1 0 2412 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6470
timestamp 1682952543
transform 1 0 2404 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6607
timestamp 1682952543
transform 1 0 2396 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6515
timestamp 1682952543
transform 1 0 2428 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6509
timestamp 1682952543
transform 1 0 2444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1682952543
transform 1 0 2460 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6608
timestamp 1682952543
transform 1 0 2436 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6609
timestamp 1682952543
transform 1 0 2452 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6600
timestamp 1682952543
transform 1 0 2452 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6516
timestamp 1682952543
transform 1 0 2484 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6445
timestamp 1682952543
transform 1 0 2500 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6511
timestamp 1682952543
transform 1 0 2492 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1682952543
transform 1 0 2500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1682952543
transform 1 0 2500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6513
timestamp 1682952543
transform 1 0 2516 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6568
timestamp 1682952543
transform 1 0 2524 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6514
timestamp 1682952543
transform 1 0 2556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6515
timestamp 1682952543
transform 1 0 2572 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6611
timestamp 1682952543
transform 1 0 2532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6612
timestamp 1682952543
transform 1 0 2548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6613
timestamp 1682952543
transform 1 0 2564 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6601
timestamp 1682952543
transform 1 0 2564 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6614
timestamp 1682952543
transform 1 0 2612 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6602
timestamp 1682952543
transform 1 0 2612 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6424
timestamp 1682952543
transform 1 0 2756 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6471
timestamp 1682952543
transform 1 0 2708 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6472
timestamp 1682952543
transform 1 0 2740 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6473
timestamp 1682952543
transform 1 0 2756 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6516
timestamp 1682952543
transform 1 0 2676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6615
timestamp 1682952543
transform 1 0 2628 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6603
timestamp 1682952543
transform 1 0 2660 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6604
timestamp 1682952543
transform 1 0 2676 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6517
timestamp 1682952543
transform 1 0 2732 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6517
timestamp 1682952543
transform 1 0 2732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1682952543
transform 1 0 2740 0 1 1417
box -2 -2 2 2
use M3_M2  M3_M2_6544
timestamp 1682952543
transform 1 0 2748 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6518
timestamp 1682952543
transform 1 0 2756 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1682952543
transform 1 0 2732 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6617
timestamp 1682952543
transform 1 0 2748 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6605
timestamp 1682952543
transform 1 0 2740 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6606
timestamp 1682952543
transform 1 0 2756 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6451
timestamp 1682952543
transform 1 0 2780 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1682952543
transform 1 0 2788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6618
timestamp 1682952543
transform 1 0 2780 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6607
timestamp 1682952543
transform 1 0 2788 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6660
timestamp 1682952543
transform 1 0 2788 0 1 1385
box -2 -2 2 2
use M3_M2  M3_M2_6425
timestamp 1682952543
transform 1 0 2796 0 1 1465
box -3 -3 3 3
use M2_M1  M2_M1_6445
timestamp 1682952543
transform 1 0 2796 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_6520
timestamp 1682952543
transform 1 0 2796 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6474
timestamp 1682952543
transform 1 0 2812 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6619
timestamp 1682952543
transform 1 0 2820 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6446
timestamp 1682952543
transform 1 0 2860 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6475
timestamp 1682952543
transform 1 0 2868 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6476
timestamp 1682952543
transform 1 0 2884 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6518
timestamp 1682952543
transform 1 0 2892 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6447
timestamp 1682952543
transform 1 0 2948 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6477
timestamp 1682952543
transform 1 0 2956 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6521
timestamp 1682952543
transform 1 0 2868 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6522
timestamp 1682952543
transform 1 0 2892 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6620
timestamp 1682952543
transform 1 0 2860 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6545
timestamp 1682952543
transform 1 0 2900 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6523
timestamp 1682952543
transform 1 0 2940 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6546
timestamp 1682952543
transform 1 0 2948 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6621
timestamp 1682952543
transform 1 0 2884 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6622
timestamp 1682952543
transform 1 0 2900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6623
timestamp 1682952543
transform 1 0 2916 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6608
timestamp 1682952543
transform 1 0 2884 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6609
timestamp 1682952543
transform 1 0 2940 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6519
timestamp 1682952543
transform 1 0 3020 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6524
timestamp 1682952543
transform 1 0 3020 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6520
timestamp 1682952543
transform 1 0 3116 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6547
timestamp 1682952543
transform 1 0 3036 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6525
timestamp 1682952543
transform 1 0 3068 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6548
timestamp 1682952543
transform 1 0 3100 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6624
timestamp 1682952543
transform 1 0 3036 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6610
timestamp 1682952543
transform 1 0 3036 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6611
timestamp 1682952543
transform 1 0 3068 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6478
timestamp 1682952543
transform 1 0 3140 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6521
timestamp 1682952543
transform 1 0 3148 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6526
timestamp 1682952543
transform 1 0 3132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1682952543
transform 1 0 3140 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6549
timestamp 1682952543
transform 1 0 3156 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6625
timestamp 1682952543
transform 1 0 3148 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6522
timestamp 1682952543
transform 1 0 3180 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6528
timestamp 1682952543
transform 1 0 3188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6529
timestamp 1682952543
transform 1 0 3204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6626
timestamp 1682952543
transform 1 0 3180 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6627
timestamp 1682952543
transform 1 0 3196 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6612
timestamp 1682952543
transform 1 0 3196 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6433
timestamp 1682952543
transform 1 0 3228 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6523
timestamp 1682952543
transform 1 0 3236 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6530
timestamp 1682952543
transform 1 0 3236 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6628
timestamp 1682952543
transform 1 0 3244 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6479
timestamp 1682952543
transform 1 0 3300 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6531
timestamp 1682952543
transform 1 0 3300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1682952543
transform 1 0 3300 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6613
timestamp 1682952543
transform 1 0 3308 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6434
timestamp 1682952543
transform 1 0 3340 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_6630
timestamp 1682952543
transform 1 0 3332 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6636
timestamp 1682952543
transform 1 0 3332 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6532
timestamp 1682952543
transform 1 0 3364 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6448
timestamp 1682952543
transform 1 0 3388 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6533
timestamp 1682952543
transform 1 0 3380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6631
timestamp 1682952543
transform 1 0 3356 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6632
timestamp 1682952543
transform 1 0 3372 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1682952543
transform 1 0 3380 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6614
timestamp 1682952543
transform 1 0 3372 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6634
timestamp 1682952543
transform 1 0 3404 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6435
timestamp 1682952543
transform 1 0 3516 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6449
timestamp 1682952543
transform 1 0 3452 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6450
timestamp 1682952543
transform 1 0 3484 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6451
timestamp 1682952543
transform 1 0 3516 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6480
timestamp 1682952543
transform 1 0 3420 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6534
timestamp 1682952543
transform 1 0 3420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1682952543
transform 1 0 3484 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6635
timestamp 1682952543
transform 1 0 3436 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6615
timestamp 1682952543
transform 1 0 3484 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6524
timestamp 1682952543
transform 1 0 3532 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6536
timestamp 1682952543
transform 1 0 3532 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6637
timestamp 1682952543
transform 1 0 3460 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6638
timestamp 1682952543
transform 1 0 3484 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6639
timestamp 1682952543
transform 1 0 3516 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6640
timestamp 1682952543
transform 1 0 3532 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6525
timestamp 1682952543
transform 1 0 3588 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6550
timestamp 1682952543
transform 1 0 3564 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6537
timestamp 1682952543
transform 1 0 3572 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6551
timestamp 1682952543
transform 1 0 3580 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6538
timestamp 1682952543
transform 1 0 3588 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1682952543
transform 1 0 3604 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6636
timestamp 1682952543
transform 1 0 3564 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1682952543
transform 1 0 3580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6638
timestamp 1682952543
transform 1 0 3596 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6616
timestamp 1682952543
transform 1 0 3572 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6641
timestamp 1682952543
transform 1 0 3564 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6642
timestamp 1682952543
transform 1 0 3604 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6481
timestamp 1682952543
transform 1 0 3628 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6540
timestamp 1682952543
transform 1 0 3628 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6426
timestamp 1682952543
transform 1 0 3652 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6482
timestamp 1682952543
transform 1 0 3668 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6483
timestamp 1682952543
transform 1 0 3684 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6526
timestamp 1682952543
transform 1 0 3660 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6552
timestamp 1682952543
transform 1 0 3644 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6639
timestamp 1682952543
transform 1 0 3636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6541
timestamp 1682952543
transform 1 0 3668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6640
timestamp 1682952543
transform 1 0 3660 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6569
timestamp 1682952543
transform 1 0 3676 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6527
timestamp 1682952543
transform 1 0 3700 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6528
timestamp 1682952543
transform 1 0 3716 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6542
timestamp 1682952543
transform 1 0 3700 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1682952543
transform 1 0 3708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6641
timestamp 1682952543
transform 1 0 3700 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6642
timestamp 1682952543
transform 1 0 3716 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6484
timestamp 1682952543
transform 1 0 3748 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6544
timestamp 1682952543
transform 1 0 3748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6545
timestamp 1682952543
transform 1 0 3764 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1682952543
transform 1 0 3772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6643
timestamp 1682952543
transform 1 0 3740 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6570
timestamp 1682952543
transform 1 0 3756 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6617
timestamp 1682952543
transform 1 0 3740 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6618
timestamp 1682952543
transform 1 0 3772 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6553
timestamp 1682952543
transform 1 0 3788 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6644
timestamp 1682952543
transform 1 0 3788 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6485
timestamp 1682952543
transform 1 0 3820 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6529
timestamp 1682952543
transform 1 0 3844 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6547
timestamp 1682952543
transform 1 0 3804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6548
timestamp 1682952543
transform 1 0 3820 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1682952543
transform 1 0 3836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6550
timestamp 1682952543
transform 1 0 3844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1682952543
transform 1 0 3804 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6646
timestamp 1682952543
transform 1 0 3812 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6571
timestamp 1682952543
transform 1 0 3820 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6647
timestamp 1682952543
transform 1 0 3828 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6648
timestamp 1682952543
transform 1 0 3844 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6643
timestamp 1682952543
transform 1 0 3820 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6452
timestamp 1682952543
transform 1 0 3876 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6486
timestamp 1682952543
transform 1 0 3868 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6572
timestamp 1682952543
transform 1 0 3860 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6649
timestamp 1682952543
transform 1 0 3868 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6644
timestamp 1682952543
transform 1 0 3852 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6453
timestamp 1682952543
transform 1 0 3892 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6454
timestamp 1682952543
transform 1 0 3916 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6487
timestamp 1682952543
transform 1 0 3892 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6551
timestamp 1682952543
transform 1 0 3900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1682952543
transform 1 0 3916 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6650
timestamp 1682952543
transform 1 0 3892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6651
timestamp 1682952543
transform 1 0 3908 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6619
timestamp 1682952543
transform 1 0 3892 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6427
timestamp 1682952543
transform 1 0 3940 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6530
timestamp 1682952543
transform 1 0 3932 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6553
timestamp 1682952543
transform 1 0 3932 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6455
timestamp 1682952543
transform 1 0 3972 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6554
timestamp 1682952543
transform 1 0 3956 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1682952543
transform 1 0 3972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6652
timestamp 1682952543
transform 1 0 3948 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6573
timestamp 1682952543
transform 1 0 3956 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6653
timestamp 1682952543
transform 1 0 3980 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6620
timestamp 1682952543
transform 1 0 3980 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6556
timestamp 1682952543
transform 1 0 3996 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6488
timestamp 1682952543
transform 1 0 4012 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6554
timestamp 1682952543
transform 1 0 4020 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6557
timestamp 1682952543
transform 1 0 4028 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6654
timestamp 1682952543
transform 1 0 4004 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6655
timestamp 1682952543
transform 1 0 4020 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6574
timestamp 1682952543
transform 1 0 4028 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6558
timestamp 1682952543
transform 1 0 4044 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6645
timestamp 1682952543
transform 1 0 4036 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6555
timestamp 1682952543
transform 1 0 4052 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6656
timestamp 1682952543
transform 1 0 4052 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6657
timestamp 1682952543
transform 1 0 4068 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6659
timestamp 1682952543
transform 1 0 4116 0 1 1395
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_54
timestamp 1682952543
transform 1 0 48 0 1 1370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_396
timestamp 1682952543
transform 1 0 72 0 1 1370
box -8 -3 104 105
use FILL  FILL_2757
timestamp 1682952543
transform 1 0 168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1682952543
transform 1 0 176 0 1 1370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1682952543
transform 1 0 184 0 1 1370
box -8 -3 16 105
use FILL  FILL_2761
timestamp 1682952543
transform 1 0 192 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_270
timestamp 1682952543
transform -1 0 240 0 1 1370
box -8 -3 46 105
use FILL  FILL_2762
timestamp 1682952543
transform 1 0 240 0 1 1370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1682952543
transform 1 0 248 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_398
timestamp 1682952543
transform 1 0 256 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_443
timestamp 1682952543
transform -1 0 368 0 1 1370
box -9 -3 26 105
use FILL  FILL_2767
timestamp 1682952543
transform 1 0 368 0 1 1370
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1682952543
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1682952543
transform 1 0 384 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_273
timestamp 1682952543
transform 1 0 392 0 1 1370
box -8 -3 46 105
use FILL  FILL_2777
timestamp 1682952543
transform 1 0 432 0 1 1370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1682952543
transform 1 0 440 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6646
timestamp 1682952543
transform 1 0 516 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6647
timestamp 1682952543
transform 1 0 548 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_399
timestamp 1682952543
transform 1 0 448 0 1 1370
box -8 -3 104 105
use FILL  FILL_2779
timestamp 1682952543
transform 1 0 544 0 1 1370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1682952543
transform 1 0 552 0 1 1370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1682952543
transform 1 0 560 0 1 1370
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1682952543
transform 1 0 568 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_276
timestamp 1682952543
transform 1 0 576 0 1 1370
box -8 -3 46 105
use FILL  FILL_2794
timestamp 1682952543
transform 1 0 616 0 1 1370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1682952543
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1682952543
transform 1 0 632 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6648
timestamp 1682952543
transform 1 0 660 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6649
timestamp 1682952543
transform 1 0 684 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6650
timestamp 1682952543
transform 1 0 708 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_400
timestamp 1682952543
transform 1 0 640 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_6651
timestamp 1682952543
transform 1 0 772 0 1 1375
box -3 -3 3 3
use OAI21X1  OAI21X1_112
timestamp 1682952543
transform 1 0 736 0 1 1370
box -8 -3 34 105
use FILL  FILL_2797
timestamp 1682952543
transform 1 0 768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1682952543
transform 1 0 776 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6652
timestamp 1682952543
transform 1 0 796 0 1 1375
box -3 -3 3 3
use FILL  FILL_2812
timestamp 1682952543
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1682952543
transform 1 0 792 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6653
timestamp 1682952543
transform 1 0 812 0 1 1375
box -3 -3 3 3
use NOR2X1  NOR2X1_85
timestamp 1682952543
transform 1 0 800 0 1 1370
box -8 -3 32 105
use FILL  FILL_2816
timestamp 1682952543
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1682952543
transform 1 0 832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1682952543
transform 1 0 840 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_401
timestamp 1682952543
transform 1 0 848 0 1 1370
box -8 -3 104 105
use FILL  FILL_2821
timestamp 1682952543
transform 1 0 944 0 1 1370
box -8 -3 16 105
use FILL  FILL_2830
timestamp 1682952543
transform 1 0 952 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_445
timestamp 1682952543
transform 1 0 960 0 1 1370
box -9 -3 26 105
use FILL  FILL_2832
timestamp 1682952543
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1682952543
transform 1 0 984 0 1 1370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1682952543
transform 1 0 992 0 1 1370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1682952543
transform 1 0 1000 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_114
timestamp 1682952543
transform 1 0 1008 0 1 1370
box -8 -3 34 105
use OAI21X1  OAI21X1_115
timestamp 1682952543
transform -1 0 1072 0 1 1370
box -8 -3 34 105
use FILL  FILL_2839
timestamp 1682952543
transform 1 0 1072 0 1 1370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1682952543
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1682952543
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1682952543
transform 1 0 1096 0 1 1370
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1682952543
transform 1 0 1104 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_117
timestamp 1682952543
transform -1 0 1144 0 1 1370
box -8 -3 34 105
use FILL  FILL_2854
timestamp 1682952543
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_402
timestamp 1682952543
transform 1 0 1152 0 1 1370
box -8 -3 104 105
use FILL  FILL_2855
timestamp 1682952543
transform 1 0 1248 0 1 1370
box -8 -3 16 105
use FILL  FILL_2856
timestamp 1682952543
transform 1 0 1256 0 1 1370
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1682952543
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6654
timestamp 1682952543
transform 1 0 1308 0 1 1375
box -3 -3 3 3
use OAI22X1  OAI22X1_277
timestamp 1682952543
transform -1 0 1312 0 1 1370
box -8 -3 46 105
use FILL  FILL_2858
timestamp 1682952543
transform 1 0 1312 0 1 1370
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1682952543
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use FILL  FILL_2860
timestamp 1682952543
transform 1 0 1328 0 1 1370
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1682952543
transform 1 0 1336 0 1 1370
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1682952543
transform 1 0 1344 0 1 1370
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1682952543
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_279
timestamp 1682952543
transform -1 0 1400 0 1 1370
box -8 -3 46 105
use FILL  FILL_2873
timestamp 1682952543
transform 1 0 1400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1682952543
transform 1 0 1408 0 1 1370
box -8 -3 16 105
use FILL  FILL_2875
timestamp 1682952543
transform 1 0 1416 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6655
timestamp 1682952543
transform 1 0 1436 0 1 1375
box -3 -3 3 3
use FILL  FILL_2876
timestamp 1682952543
transform 1 0 1424 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_404
timestamp 1682952543
transform 1 0 1432 0 1 1370
box -8 -3 104 105
use FILL  FILL_2877
timestamp 1682952543
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6656
timestamp 1682952543
transform 1 0 1548 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_447
timestamp 1682952543
transform 1 0 1536 0 1 1370
box -9 -3 26 105
use FILL  FILL_2878
timestamp 1682952543
transform 1 0 1552 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_450
timestamp 1682952543
transform 1 0 1560 0 1 1370
box -9 -3 26 105
use FILL  FILL_2889
timestamp 1682952543
transform 1 0 1576 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_406
timestamp 1682952543
transform 1 0 1584 0 1 1370
box -8 -3 104 105
use FILL  FILL_2890
timestamp 1682952543
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_451
timestamp 1682952543
transform 1 0 1688 0 1 1370
box -9 -3 26 105
use FILL  FILL_2893
timestamp 1682952543
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_2895
timestamp 1682952543
transform 1 0 1712 0 1 1370
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1682952543
transform 1 0 1720 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_119
timestamp 1682952543
transform -1 0 1760 0 1 1370
box -8 -3 34 105
use FILL  FILL_2898
timestamp 1682952543
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1682952543
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1682952543
transform 1 0 1776 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_120
timestamp 1682952543
transform 1 0 1784 0 1 1370
box -8 -3 34 105
use FILL  FILL_2904
timestamp 1682952543
transform 1 0 1816 0 1 1370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1682952543
transform 1 0 1824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1682952543
transform 1 0 1832 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_121
timestamp 1682952543
transform -1 0 1872 0 1 1370
box -8 -3 34 105
use INVX2  INVX2_455
timestamp 1682952543
transform 1 0 1872 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_456
timestamp 1682952543
transform 1 0 1888 0 1 1370
box -9 -3 26 105
use FILL  FILL_2911
timestamp 1682952543
transform 1 0 1904 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_457
timestamp 1682952543
transform 1 0 1912 0 1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_408
timestamp 1682952543
transform 1 0 1928 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_6657
timestamp 1682952543
transform 1 0 2036 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_458
timestamp 1682952543
transform 1 0 2024 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6658
timestamp 1682952543
transform 1 0 2060 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_409
timestamp 1682952543
transform 1 0 2040 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_6659
timestamp 1682952543
transform 1 0 2148 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_459
timestamp 1682952543
transform 1 0 2136 0 1 1370
box -9 -3 26 105
use FILL  FILL_2912
timestamp 1682952543
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use FILL  FILL_2913
timestamp 1682952543
transform 1 0 2160 0 1 1370
box -8 -3 16 105
use FILL  FILL_2929
timestamp 1682952543
transform 1 0 2168 0 1 1370
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1682952543
transform 1 0 2176 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_286
timestamp 1682952543
transform 1 0 2184 0 1 1370
box -8 -3 46 105
use FILL  FILL_2933
timestamp 1682952543
transform 1 0 2224 0 1 1370
box -8 -3 16 105
use FILL  FILL_2934
timestamp 1682952543
transform 1 0 2232 0 1 1370
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1682952543
transform 1 0 2240 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_410
timestamp 1682952543
transform 1 0 2248 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_461
timestamp 1682952543
transform 1 0 2344 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_462
timestamp 1682952543
transform 1 0 2360 0 1 1370
box -9 -3 26 105
use FILL  FILL_2939
timestamp 1682952543
transform 1 0 2376 0 1 1370
box -8 -3 16 105
use FILL  FILL_2940
timestamp 1682952543
transform 1 0 2384 0 1 1370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1682952543
transform 1 0 2392 0 1 1370
box -8 -3 16 105
use FILL  FILL_2942
timestamp 1682952543
transform 1 0 2400 0 1 1370
box -8 -3 16 105
use FILL  FILL_2954
timestamp 1682952543
transform 1 0 2408 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_289
timestamp 1682952543
transform 1 0 2416 0 1 1370
box -8 -3 46 105
use FILL  FILL_2955
timestamp 1682952543
transform 1 0 2456 0 1 1370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1682952543
transform 1 0 2464 0 1 1370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1682952543
transform 1 0 2472 0 1 1370
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1682952543
transform 1 0 2480 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_465
timestamp 1682952543
transform -1 0 2504 0 1 1370
box -9 -3 26 105
use FILL  FILL_2959
timestamp 1682952543
transform 1 0 2504 0 1 1370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1682952543
transform 1 0 2512 0 1 1370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1682952543
transform 1 0 2520 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_290
timestamp 1682952543
transform 1 0 2528 0 1 1370
box -8 -3 46 105
use FILL  FILL_2964
timestamp 1682952543
transform 1 0 2568 0 1 1370
box -8 -3 16 105
use FILL  FILL_2965
timestamp 1682952543
transform 1 0 2576 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_466
timestamp 1682952543
transform -1 0 2600 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6660
timestamp 1682952543
transform 1 0 2612 0 1 1375
box -3 -3 3 3
use FILL  FILL_2966
timestamp 1682952543
transform 1 0 2600 0 1 1370
box -8 -3 16 105
use FILL  FILL_2967
timestamp 1682952543
transform 1 0 2608 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6661
timestamp 1682952543
transform 1 0 2628 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6662
timestamp 1682952543
transform 1 0 2676 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_412
timestamp 1682952543
transform 1 0 2616 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_467
timestamp 1682952543
transform 1 0 2712 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6663
timestamp 1682952543
transform 1 0 2748 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6664
timestamp 1682952543
transform 1 0 2772 0 1 1375
box -3 -3 3 3
use OAI22X1  OAI22X1_291
timestamp 1682952543
transform 1 0 2728 0 1 1370
box -8 -3 46 105
use FILL  FILL_2968
timestamp 1682952543
transform 1 0 2768 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6665
timestamp 1682952543
transform 1 0 2788 0 1 1375
box -3 -3 3 3
use FILL  FILL_2969
timestamp 1682952543
transform 1 0 2776 0 1 1370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1682952543
transform 1 0 2784 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6666
timestamp 1682952543
transform 1 0 2804 0 1 1375
box -3 -3 3 3
use FILL  FILL_2971
timestamp 1682952543
transform 1 0 2792 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_468
timestamp 1682952543
transform 1 0 2800 0 1 1370
box -9 -3 26 105
use FILL  FILL_2972
timestamp 1682952543
transform 1 0 2816 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6667
timestamp 1682952543
transform 1 0 2836 0 1 1375
box -3 -3 3 3
use FILL  FILL_2977
timestamp 1682952543
transform 1 0 2824 0 1 1370
box -8 -3 16 105
use FILL  FILL_2979
timestamp 1682952543
transform 1 0 2832 0 1 1370
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1682952543
transform 1 0 2840 0 1 1370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1682952543
transform 1 0 2848 0 1 1370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1682952543
transform 1 0 2856 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6668
timestamp 1682952543
transform 1 0 2900 0 1 1375
box -3 -3 3 3
use OAI22X1  OAI22X1_294
timestamp 1682952543
transform 1 0 2864 0 1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_415
timestamp 1682952543
transform 1 0 2904 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_469
timestamp 1682952543
transform 1 0 3000 0 1 1370
box -9 -3 26 105
use FILL  FILL_2986
timestamp 1682952543
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6669
timestamp 1682952543
transform 1 0 3052 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_416
timestamp 1682952543
transform 1 0 3024 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_470
timestamp 1682952543
transform 1 0 3120 0 1 1370
box -9 -3 26 105
use FILL  FILL_2987
timestamp 1682952543
transform 1 0 3136 0 1 1370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1682952543
transform 1 0 3144 0 1 1370
box -8 -3 16 105
use FILL  FILL_2989
timestamp 1682952543
transform 1 0 3152 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6670
timestamp 1682952543
transform 1 0 3196 0 1 1375
box -3 -3 3 3
use OAI22X1  OAI22X1_297
timestamp 1682952543
transform 1 0 3160 0 1 1370
box -8 -3 46 105
use FILL  FILL_3003
timestamp 1682952543
transform 1 0 3200 0 1 1370
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1682952543
transform 1 0 3208 0 1 1370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1682952543
transform 1 0 3216 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_471
timestamp 1682952543
transform -1 0 3240 0 1 1370
box -9 -3 26 105
use FILL  FILL_3012
timestamp 1682952543
transform 1 0 3240 0 1 1370
box -8 -3 16 105
use FILL  FILL_3013
timestamp 1682952543
transform 1 0 3248 0 1 1370
box -8 -3 16 105
use FILL  FILL_3014
timestamp 1682952543
transform 1 0 3256 0 1 1370
box -8 -3 16 105
use FILL  FILL_3015
timestamp 1682952543
transform 1 0 3264 0 1 1370
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1682952543
transform 1 0 3272 0 1 1370
box -8 -3 16 105
use FILL  FILL_3017
timestamp 1682952543
transform 1 0 3280 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_472
timestamp 1682952543
transform -1 0 3304 0 1 1370
box -9 -3 26 105
use FILL  FILL_3018
timestamp 1682952543
transform 1 0 3304 0 1 1370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1682952543
transform 1 0 3312 0 1 1370
box -8 -3 16 105
use FILL  FILL_3022
timestamp 1682952543
transform 1 0 3320 0 1 1370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1682952543
transform 1 0 3328 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6671
timestamp 1682952543
transform 1 0 3348 0 1 1375
box -3 -3 3 3
use OAI22X1  OAI22X1_298
timestamp 1682952543
transform 1 0 3336 0 1 1370
box -8 -3 46 105
use FILL  FILL_3026
timestamp 1682952543
transform 1 0 3376 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6672
timestamp 1682952543
transform 1 0 3404 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_473
timestamp 1682952543
transform 1 0 3384 0 1 1370
box -9 -3 26 105
use BUFX2  BUFX2_93
timestamp 1682952543
transform -1 0 3424 0 1 1370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_418
timestamp 1682952543
transform 1 0 3424 0 1 1370
box -8 -3 104 105
use M3_M2  M3_M2_6673
timestamp 1682952543
transform 1 0 3540 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_474
timestamp 1682952543
transform 1 0 3520 0 1 1370
box -9 -3 26 105
use FILL  FILL_3027
timestamp 1682952543
transform 1 0 3536 0 1 1370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1682952543
transform 1 0 3544 0 1 1370
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1682952543
transform 1 0 3552 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6674
timestamp 1682952543
transform 1 0 3572 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6675
timestamp 1682952543
transform 1 0 3596 0 1 1375
box -3 -3 3 3
use OAI22X1  OAI22X1_299
timestamp 1682952543
transform 1 0 3560 0 1 1370
box -8 -3 46 105
use FILL  FILL_3030
timestamp 1682952543
transform 1 0 3600 0 1 1370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1682952543
transform 1 0 3608 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_475
timestamp 1682952543
transform -1 0 3632 0 1 1370
box -9 -3 26 105
use FILL  FILL_3032
timestamp 1682952543
transform 1 0 3632 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_94
timestamp 1682952543
transform 1 0 3640 0 1 1370
box -5 -3 28 105
use BUFX2  BUFX2_95
timestamp 1682952543
transform 1 0 3664 0 1 1370
box -5 -3 28 105
use FILL  FILL_3033
timestamp 1682952543
transform 1 0 3688 0 1 1370
box -8 -3 16 105
use FILL  FILL_3045
timestamp 1682952543
transform 1 0 3696 0 1 1370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1682952543
transform 1 0 3704 0 1 1370
box -8 -3 16 105
use FILL  FILL_3048
timestamp 1682952543
transform 1 0 3712 0 1 1370
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1682952543
transform 1 0 3720 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6676
timestamp 1682952543
transform 1 0 3740 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6677
timestamp 1682952543
transform 1 0 3764 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_283
timestamp 1682952543
transform 1 0 3728 0 1 1370
box -8 -3 46 105
use FILL  FILL_3050
timestamp 1682952543
transform 1 0 3768 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6678
timestamp 1682952543
transform 1 0 3788 0 1 1375
box -3 -3 3 3
use FILL  FILL_3051
timestamp 1682952543
transform 1 0 3776 0 1 1370
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1682952543
transform 1 0 3784 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_476
timestamp 1682952543
transform -1 0 3808 0 1 1370
box -9 -3 26 105
use OAI22X1  OAI22X1_301
timestamp 1682952543
transform -1 0 3848 0 1 1370
box -8 -3 46 105
use M3_M2  M3_M2_6679
timestamp 1682952543
transform 1 0 3860 0 1 1375
box -3 -3 3 3
use FILL  FILL_3053
timestamp 1682952543
transform 1 0 3848 0 1 1370
box -8 -3 16 105
use FILL  FILL_3054
timestamp 1682952543
transform 1 0 3856 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6680
timestamp 1682952543
transform 1 0 3876 0 1 1375
box -3 -3 3 3
use FILL  FILL_3055
timestamp 1682952543
transform 1 0 3864 0 1 1370
box -8 -3 16 105
use FILL  FILL_3056
timestamp 1682952543
transform 1 0 3872 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6681
timestamp 1682952543
transform 1 0 3900 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_284
timestamp 1682952543
transform 1 0 3880 0 1 1370
box -8 -3 46 105
use FILL  FILL_3057
timestamp 1682952543
transform 1 0 3920 0 1 1370
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1682952543
transform 1 0 3928 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6682
timestamp 1682952543
transform 1 0 3964 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6683
timestamp 1682952543
transform 1 0 3980 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_285
timestamp 1682952543
transform 1 0 3936 0 1 1370
box -8 -3 46 105
use FILL  FILL_3059
timestamp 1682952543
transform 1 0 3976 0 1 1370
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1682952543
transform 1 0 3984 0 1 1370
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1682952543
transform 1 0 3992 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_303
timestamp 1682952543
transform 1 0 4000 0 1 1370
box -8 -3 46 105
use FILL  FILL_3066
timestamp 1682952543
transform 1 0 4040 0 1 1370
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1682952543
transform 1 0 4048 0 1 1370
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1682952543
transform 1 0 4056 0 1 1370
box -8 -3 16 105
use FILL  FILL_3069
timestamp 1682952543
transform 1 0 4064 0 1 1370
box -8 -3 16 105
use FILL  FILL_3070
timestamp 1682952543
transform 1 0 4072 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_479
timestamp 1682952543
transform -1 0 4096 0 1 1370
box -9 -3 26 105
use FILL  FILL_3071
timestamp 1682952543
transform 1 0 4096 0 1 1370
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1682952543
transform 1 0 4104 0 1 1370
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1682952543
transform 1 0 4112 0 1 1370
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1682952543
transform 1 0 4120 0 1 1370
box -8 -3 16 105
use FILL  FILL_3075
timestamp 1682952543
transform 1 0 4128 0 1 1370
box -8 -3 16 105
use FILL  FILL_3076
timestamp 1682952543
transform 1 0 4136 0 1 1370
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1682952543
transform 1 0 4144 0 1 1370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_55
timestamp 1682952543
transform 1 0 4177 0 1 1370
box -10 -3 10 3
use M2_M1  M2_M1_6668
timestamp 1682952543
transform 1 0 84 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6779
timestamp 1682952543
transform 1 0 132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6780
timestamp 1682952543
transform 1 0 164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6781
timestamp 1682952543
transform 1 0 172 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6837
timestamp 1682952543
transform 1 0 132 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6838
timestamp 1682952543
transform 1 0 172 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6878
timestamp 1682952543
transform 1 0 164 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6782
timestamp 1682952543
transform 1 0 196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6669
timestamp 1682952543
transform 1 0 212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1682952543
transform 1 0 220 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6671
timestamp 1682952543
transform 1 0 236 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6783
timestamp 1682952543
transform 1 0 228 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6879
timestamp 1682952543
transform 1 0 220 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6784
timestamp 1682952543
transform 1 0 268 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6785
timestamp 1682952543
transform 1 0 276 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6905
timestamp 1682952543
transform 1 0 268 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_6672
timestamp 1682952543
transform 1 0 292 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6783
timestamp 1682952543
transform 1 0 300 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6786
timestamp 1682952543
transform 1 0 300 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6736
timestamp 1682952543
transform 1 0 340 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6684
timestamp 1682952543
transform 1 0 364 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6705
timestamp 1682952543
transform 1 0 364 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6737
timestamp 1682952543
transform 1 0 380 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6673
timestamp 1682952543
transform 1 0 340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6674
timestamp 1682952543
transform 1 0 348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6675
timestamp 1682952543
transform 1 0 364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6676
timestamp 1682952543
transform 1 0 380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6787
timestamp 1682952543
transform 1 0 340 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6839
timestamp 1682952543
transform 1 0 340 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6906
timestamp 1682952543
transform 1 0 332 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_6788
timestamp 1682952543
transform 1 0 356 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6789
timestamp 1682952543
transform 1 0 372 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6784
timestamp 1682952543
transform 1 0 388 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6790
timestamp 1682952543
transform 1 0 388 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6926
timestamp 1682952543
transform 1 0 388 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6738
timestamp 1682952543
transform 1 0 404 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6677
timestamp 1682952543
transform 1 0 404 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6685
timestamp 1682952543
transform 1 0 460 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6785
timestamp 1682952543
transform 1 0 452 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6791
timestamp 1682952543
transform 1 0 436 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6792
timestamp 1682952543
transform 1 0 452 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6840
timestamp 1682952543
transform 1 0 452 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_6678
timestamp 1682952543
transform 1 0 468 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6679
timestamp 1682952543
transform 1 0 476 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6813
timestamp 1682952543
transform 1 0 468 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6686
timestamp 1682952543
transform 1 0 500 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6786
timestamp 1682952543
transform 1 0 492 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6793
timestamp 1682952543
transform 1 0 484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6794
timestamp 1682952543
transform 1 0 492 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6841
timestamp 1682952543
transform 1 0 476 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6814
timestamp 1682952543
transform 1 0 500 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6687
timestamp 1682952543
transform 1 0 532 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6739
timestamp 1682952543
transform 1 0 540 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6680
timestamp 1682952543
transform 1 0 524 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6787
timestamp 1682952543
transform 1 0 532 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6681
timestamp 1682952543
transform 1 0 540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6795
timestamp 1682952543
transform 1 0 532 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6815
timestamp 1682952543
transform 1 0 540 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6796
timestamp 1682952543
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6842
timestamp 1682952543
transform 1 0 532 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6907
timestamp 1682952543
transform 1 0 548 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_6797
timestamp 1682952543
transform 1 0 580 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6740
timestamp 1682952543
transform 1 0 612 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6682
timestamp 1682952543
transform 1 0 612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6798
timestamp 1682952543
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6880
timestamp 1682952543
transform 1 0 628 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6706
timestamp 1682952543
transform 1 0 644 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6661
timestamp 1682952543
transform 1 0 652 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1682952543
transform 1 0 644 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_6799
timestamp 1682952543
transform 1 0 644 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6843
timestamp 1682952543
transform 1 0 644 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6688
timestamp 1682952543
transform 1 0 668 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_6662
timestamp 1682952543
transform 1 0 676 0 1 1355
box -2 -2 2 2
use M3_M2  M3_M2_6707
timestamp 1682952543
transform 1 0 684 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6683
timestamp 1682952543
transform 1 0 684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1682952543
transform 1 0 692 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6708
timestamp 1682952543
transform 1 0 724 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6709
timestamp 1682952543
transform 1 0 740 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6741
timestamp 1682952543
transform 1 0 716 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6663
timestamp 1682952543
transform 1 0 756 0 1 1355
box -2 -2 2 2
use M2_M1  M2_M1_6685
timestamp 1682952543
transform 1 0 716 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6788
timestamp 1682952543
transform 1 0 724 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6789
timestamp 1682952543
transform 1 0 748 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6686
timestamp 1682952543
transform 1 0 756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6800
timestamp 1682952543
transform 1 0 708 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6801
timestamp 1682952543
transform 1 0 716 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6802
timestamp 1682952543
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6803
timestamp 1682952543
transform 1 0 748 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6908
timestamp 1682952543
transform 1 0 716 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6844
timestamp 1682952543
transform 1 0 748 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6710
timestamp 1682952543
transform 1 0 780 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6664
timestamp 1682952543
transform 1 0 788 0 1 1355
box -2 -2 2 2
use M3_M2  M3_M2_6790
timestamp 1682952543
transform 1 0 788 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6804
timestamp 1682952543
transform 1 0 788 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6845
timestamp 1682952543
transform 1 0 796 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6742
timestamp 1682952543
transform 1 0 836 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6687
timestamp 1682952543
transform 1 0 828 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6805
timestamp 1682952543
transform 1 0 828 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6846
timestamp 1682952543
transform 1 0 812 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6927
timestamp 1682952543
transform 1 0 828 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_6688
timestamp 1682952543
transform 1 0 836 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6689
timestamp 1682952543
transform 1 0 860 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_6888
timestamp 1682952543
transform 1 0 876 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6881
timestamp 1682952543
transform 1 0 876 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6928
timestamp 1682952543
transform 1 0 876 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_6689
timestamp 1682952543
transform 1 0 892 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6791
timestamp 1682952543
transform 1 0 900 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6690
timestamp 1682952543
transform 1 0 916 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6691
timestamp 1682952543
transform 1 0 924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6692
timestamp 1682952543
transform 1 0 932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6806
timestamp 1682952543
transform 1 0 908 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6816
timestamp 1682952543
transform 1 0 924 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6711
timestamp 1682952543
transform 1 0 948 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6743
timestamp 1682952543
transform 1 0 940 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6882
timestamp 1682952543
transform 1 0 932 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6817
timestamp 1682952543
transform 1 0 972 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6744
timestamp 1682952543
transform 1 0 1012 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6818
timestamp 1682952543
transform 1 0 996 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6889
timestamp 1682952543
transform 1 0 996 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6883
timestamp 1682952543
transform 1 0 996 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6929
timestamp 1682952543
transform 1 0 996 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6745
timestamp 1682952543
transform 1 0 1028 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6792
timestamp 1682952543
transform 1 0 1020 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6693
timestamp 1682952543
transform 1 0 1028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6694
timestamp 1682952543
transform 1 0 1036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6890
timestamp 1682952543
transform 1 0 1028 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6884
timestamp 1682952543
transform 1 0 1028 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6909
timestamp 1682952543
transform 1 0 1028 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6819
timestamp 1682952543
transform 1 0 1044 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6793
timestamp 1682952543
transform 1 0 1068 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6807
timestamp 1682952543
transform 1 0 1060 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6930
timestamp 1682952543
transform 1 0 1052 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_6891
timestamp 1682952543
transform 1 0 1092 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6712
timestamp 1682952543
transform 1 0 1108 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6746
timestamp 1682952543
transform 1 0 1132 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6695
timestamp 1682952543
transform 1 0 1140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6808
timestamp 1682952543
transform 1 0 1108 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6809
timestamp 1682952543
transform 1 0 1124 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6810
timestamp 1682952543
transform 1 0 1132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6892
timestamp 1682952543
transform 1 0 1108 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6931
timestamp 1682952543
transform 1 0 1140 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6690
timestamp 1682952543
transform 1 0 1156 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6691
timestamp 1682952543
transform 1 0 1204 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6692
timestamp 1682952543
transform 1 0 1220 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6693
timestamp 1682952543
transform 1 0 1252 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6747
timestamp 1682952543
transform 1 0 1260 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6696
timestamp 1682952543
transform 1 0 1260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6811
timestamp 1682952543
transform 1 0 1212 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6910
timestamp 1682952543
transform 1 0 1196 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_6697
timestamp 1682952543
transform 1 0 1276 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6794
timestamp 1682952543
transform 1 0 1316 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6698
timestamp 1682952543
transform 1 0 1324 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6795
timestamp 1682952543
transform 1 0 1332 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6812
timestamp 1682952543
transform 1 0 1316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6813
timestamp 1682952543
transform 1 0 1332 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6847
timestamp 1682952543
transform 1 0 1316 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_6814
timestamp 1682952543
transform 1 0 1348 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1682952543
transform 1 0 1372 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6694
timestamp 1682952543
transform 1 0 1388 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6695
timestamp 1682952543
transform 1 0 1444 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6748
timestamp 1682952543
transform 1 0 1388 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6700
timestamp 1682952543
transform 1 0 1388 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6796
timestamp 1682952543
transform 1 0 1412 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6815
timestamp 1682952543
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6932
timestamp 1682952543
transform 1 0 1404 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6820
timestamp 1682952543
transform 1 0 1484 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6797
timestamp 1682952543
transform 1 0 1508 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6816
timestamp 1682952543
transform 1 0 1500 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6817
timestamp 1682952543
transform 1 0 1508 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6848
timestamp 1682952543
transform 1 0 1500 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6713
timestamp 1682952543
transform 1 0 1524 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6701
timestamp 1682952543
transform 1 0 1540 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6821
timestamp 1682952543
transform 1 0 1540 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6818
timestamp 1682952543
transform 1 0 1548 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6911
timestamp 1682952543
transform 1 0 1548 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_6702
timestamp 1682952543
transform 1 0 1556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6703
timestamp 1682952543
transform 1 0 1572 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6819
timestamp 1682952543
transform 1 0 1588 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6849
timestamp 1682952543
transform 1 0 1588 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6749
timestamp 1682952543
transform 1 0 1652 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6704
timestamp 1682952543
transform 1 0 1604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6705
timestamp 1682952543
transform 1 0 1692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6820
timestamp 1682952543
transform 1 0 1652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6821
timestamp 1682952543
transform 1 0 1684 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6912
timestamp 1682952543
transform 1 0 1636 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6933
timestamp 1682952543
transform 1 0 1676 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_6822
timestamp 1682952543
transform 1 0 1708 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6750
timestamp 1682952543
transform 1 0 1748 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6706
timestamp 1682952543
transform 1 0 1732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6707
timestamp 1682952543
transform 1 0 1748 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6798
timestamp 1682952543
transform 1 0 1756 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6708
timestamp 1682952543
transform 1 0 1764 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6822
timestamp 1682952543
transform 1 0 1732 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6823
timestamp 1682952543
transform 1 0 1740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6893
timestamp 1682952543
transform 1 0 1772 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6885
timestamp 1682952543
transform 1 0 1772 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6709
timestamp 1682952543
transform 1 0 1796 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6696
timestamp 1682952543
transform 1 0 1828 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_6710
timestamp 1682952543
transform 1 0 1820 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6850
timestamp 1682952543
transform 1 0 1820 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6913
timestamp 1682952543
transform 1 0 1820 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6751
timestamp 1682952543
transform 1 0 1852 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6714
timestamp 1682952543
transform 1 0 1876 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6711
timestamp 1682952543
transform 1 0 1852 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1682952543
transform 1 0 1868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1682952543
transform 1 0 1876 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6824
timestamp 1682952543
transform 1 0 1836 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6825
timestamp 1682952543
transform 1 0 1844 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6826
timestamp 1682952543
transform 1 0 1860 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6823
timestamp 1682952543
transform 1 0 1868 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6827
timestamp 1682952543
transform 1 0 1876 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6851
timestamp 1682952543
transform 1 0 1836 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6852
timestamp 1682952543
transform 1 0 1860 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6886
timestamp 1682952543
transform 1 0 1844 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6853
timestamp 1682952543
transform 1 0 1884 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6887
timestamp 1682952543
transform 1 0 1876 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6715
timestamp 1682952543
transform 1 0 1900 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6714
timestamp 1682952543
transform 1 0 1908 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6715
timestamp 1682952543
transform 1 0 1924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6828
timestamp 1682952543
transform 1 0 1916 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6829
timestamp 1682952543
transform 1 0 1932 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6824
timestamp 1682952543
transform 1 0 1940 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6854
timestamp 1682952543
transform 1 0 1932 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_6830
timestamp 1682952543
transform 1 0 1956 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6888
timestamp 1682952543
transform 1 0 1956 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6752
timestamp 1682952543
transform 1 0 1988 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6716
timestamp 1682952543
transform 1 0 1972 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1682952543
transform 1 0 1980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1682952543
transform 1 0 1996 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1682952543
transform 1 0 2012 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6831
timestamp 1682952543
transform 1 0 2004 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6825
timestamp 1682952543
transform 1 0 2012 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6826
timestamp 1682952543
transform 1 0 2028 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6914
timestamp 1682952543
transform 1 0 2036 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6753
timestamp 1682952543
transform 1 0 2052 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6716
timestamp 1682952543
transform 1 0 2084 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6720
timestamp 1682952543
transform 1 0 2052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1682952543
transform 1 0 2068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1682952543
transform 1 0 2084 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6827
timestamp 1682952543
transform 1 0 2052 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6832
timestamp 1682952543
transform 1 0 2060 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6833
timestamp 1682952543
transform 1 0 2076 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6855
timestamp 1682952543
transform 1 0 2084 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6889
timestamp 1682952543
transform 1 0 2076 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6915
timestamp 1682952543
transform 1 0 2076 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6697
timestamp 1682952543
transform 1 0 2100 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6698
timestamp 1682952543
transform 1 0 2124 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6754
timestamp 1682952543
transform 1 0 2116 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6755
timestamp 1682952543
transform 1 0 2156 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6723
timestamp 1682952543
transform 1 0 2124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1682952543
transform 1 0 2140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1682952543
transform 1 0 2156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6834
timestamp 1682952543
transform 1 0 2148 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6717
timestamp 1682952543
transform 1 0 2172 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6835
timestamp 1682952543
transform 1 0 2172 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6856
timestamp 1682952543
transform 1 0 2164 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6916
timestamp 1682952543
transform 1 0 2172 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6756
timestamp 1682952543
transform 1 0 2228 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6726
timestamp 1682952543
transform 1 0 2196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6727
timestamp 1682952543
transform 1 0 2212 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6728
timestamp 1682952543
transform 1 0 2228 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6857
timestamp 1682952543
transform 1 0 2188 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_6836
timestamp 1682952543
transform 1 0 2220 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6890
timestamp 1682952543
transform 1 0 2220 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6837
timestamp 1682952543
transform 1 0 2236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6729
timestamp 1682952543
transform 1 0 2316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6894
timestamp 1682952543
transform 1 0 2316 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6718
timestamp 1682952543
transform 1 0 2332 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6730
timestamp 1682952543
transform 1 0 2340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6838
timestamp 1682952543
transform 1 0 2332 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6839
timestamp 1682952543
transform 1 0 2348 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6719
timestamp 1682952543
transform 1 0 2372 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6757
timestamp 1682952543
transform 1 0 2364 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6731
timestamp 1682952543
transform 1 0 2364 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6840
timestamp 1682952543
transform 1 0 2364 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6699
timestamp 1682952543
transform 1 0 2412 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6700
timestamp 1682952543
transform 1 0 2476 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6701
timestamp 1682952543
transform 1 0 2492 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_6732
timestamp 1682952543
transform 1 0 2404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6733
timestamp 1682952543
transform 1 0 2420 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6841
timestamp 1682952543
transform 1 0 2444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6842
timestamp 1682952543
transform 1 0 2500 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6858
timestamp 1682952543
transform 1 0 2468 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6859
timestamp 1682952543
transform 1 0 2500 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6720
timestamp 1682952543
transform 1 0 2516 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6702
timestamp 1682952543
transform 1 0 2532 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6721
timestamp 1682952543
transform 1 0 2556 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6758
timestamp 1682952543
transform 1 0 2548 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6734
timestamp 1682952543
transform 1 0 2524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6735
timestamp 1682952543
transform 1 0 2540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6843
timestamp 1682952543
transform 1 0 2516 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6844
timestamp 1682952543
transform 1 0 2548 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6860
timestamp 1682952543
transform 1 0 2548 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6891
timestamp 1682952543
transform 1 0 2532 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6736
timestamp 1682952543
transform 1 0 2564 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6722
timestamp 1682952543
transform 1 0 2580 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6723
timestamp 1682952543
transform 1 0 2620 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6724
timestamp 1682952543
transform 1 0 2668 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6759
timestamp 1682952543
transform 1 0 2604 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6760
timestamp 1682952543
transform 1 0 2644 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6737
timestamp 1682952543
transform 1 0 2580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6845
timestamp 1682952543
transform 1 0 2604 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6828
timestamp 1682952543
transform 1 0 2628 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6761
timestamp 1682952543
transform 1 0 2692 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6762
timestamp 1682952543
transform 1 0 2724 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6738
timestamp 1682952543
transform 1 0 2676 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6846
timestamp 1682952543
transform 1 0 2660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6847
timestamp 1682952543
transform 1 0 2724 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6861
timestamp 1682952543
transform 1 0 2652 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6892
timestamp 1682952543
transform 1 0 2572 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6893
timestamp 1682952543
transform 1 0 2628 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6917
timestamp 1682952543
transform 1 0 2612 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6862
timestamp 1682952543
transform 1 0 2708 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6894
timestamp 1682952543
transform 1 0 2724 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6725
timestamp 1682952543
transform 1 0 2796 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6763
timestamp 1682952543
transform 1 0 2788 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6739
timestamp 1682952543
transform 1 0 2772 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6799
timestamp 1682952543
transform 1 0 2780 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6740
timestamp 1682952543
transform 1 0 2788 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6741
timestamp 1682952543
transform 1 0 2804 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6848
timestamp 1682952543
transform 1 0 2764 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6849
timestamp 1682952543
transform 1 0 2772 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6850
timestamp 1682952543
transform 1 0 2796 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6863
timestamp 1682952543
transform 1 0 2772 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6864
timestamp 1682952543
transform 1 0 2788 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6800
timestamp 1682952543
transform 1 0 2820 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6829
timestamp 1682952543
transform 1 0 2844 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6895
timestamp 1682952543
transform 1 0 2844 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6918
timestamp 1682952543
transform 1 0 2844 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6726
timestamp 1682952543
transform 1 0 2884 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6764
timestamp 1682952543
transform 1 0 2868 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6765
timestamp 1682952543
transform 1 0 2892 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6742
timestamp 1682952543
transform 1 0 2868 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6801
timestamp 1682952543
transform 1 0 2876 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6743
timestamp 1682952543
transform 1 0 2884 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6830
timestamp 1682952543
transform 1 0 2868 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6851
timestamp 1682952543
transform 1 0 2876 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6852
timestamp 1682952543
transform 1 0 2892 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6865
timestamp 1682952543
transform 1 0 2892 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6727
timestamp 1682952543
transform 1 0 2908 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6665
timestamp 1682952543
transform 1 0 2916 0 1 1355
box -2 -2 2 2
use M3_M2  M3_M2_6802
timestamp 1682952543
transform 1 0 2916 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6666
timestamp 1682952543
transform 1 0 2940 0 1 1355
box -2 -2 2 2
use M3_M2  M3_M2_6728
timestamp 1682952543
transform 1 0 2980 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6766
timestamp 1682952543
transform 1 0 2948 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6767
timestamp 1682952543
transform 1 0 2964 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6744
timestamp 1682952543
transform 1 0 2948 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6803
timestamp 1682952543
transform 1 0 2956 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6745
timestamp 1682952543
transform 1 0 2964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6746
timestamp 1682952543
transform 1 0 2980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6853
timestamp 1682952543
transform 1 0 2956 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6854
timestamp 1682952543
transform 1 0 2972 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6895
timestamp 1682952543
transform 1 0 2948 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6804
timestamp 1682952543
transform 1 0 2988 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6855
timestamp 1682952543
transform 1 0 2988 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6896
timestamp 1682952543
transform 1 0 2988 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6747
timestamp 1682952543
transform 1 0 3012 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6729
timestamp 1682952543
transform 1 0 3052 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6730
timestamp 1682952543
transform 1 0 3084 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6768
timestamp 1682952543
transform 1 0 3044 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6769
timestamp 1682952543
transform 1 0 3092 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6748
timestamp 1682952543
transform 1 0 3036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6749
timestamp 1682952543
transform 1 0 3052 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6750
timestamp 1682952543
transform 1 0 3060 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6751
timestamp 1682952543
transform 1 0 3068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6752
timestamp 1682952543
transform 1 0 3084 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6753
timestamp 1682952543
transform 1 0 3092 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6856
timestamp 1682952543
transform 1 0 3044 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6857
timestamp 1682952543
transform 1 0 3076 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6866
timestamp 1682952543
transform 1 0 3060 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6770
timestamp 1682952543
transform 1 0 3132 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6771
timestamp 1682952543
transform 1 0 3148 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6858
timestamp 1682952543
transform 1 0 3116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6859
timestamp 1682952543
transform 1 0 3132 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6860
timestamp 1682952543
transform 1 0 3148 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6867
timestamp 1682952543
transform 1 0 3148 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_6861
timestamp 1682952543
transform 1 0 3164 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6934
timestamp 1682952543
transform 1 0 3156 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6772
timestamp 1682952543
transform 1 0 3188 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6805
timestamp 1682952543
transform 1 0 3180 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6862
timestamp 1682952543
transform 1 0 3180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6754
timestamp 1682952543
transform 1 0 3204 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6731
timestamp 1682952543
transform 1 0 3236 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6773
timestamp 1682952543
transform 1 0 3220 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6755
timestamp 1682952543
transform 1 0 3220 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6806
timestamp 1682952543
transform 1 0 3244 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6863
timestamp 1682952543
transform 1 0 3244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6864
timestamp 1682952543
transform 1 0 3300 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6868
timestamp 1682952543
transform 1 0 3220 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6869
timestamp 1682952543
transform 1 0 3332 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6807
timestamp 1682952543
transform 1 0 3356 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6774
timestamp 1682952543
transform 1 0 3460 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6808
timestamp 1682952543
transform 1 0 3412 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6756
timestamp 1682952543
transform 1 0 3460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6865
timestamp 1682952543
transform 1 0 3380 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6866
timestamp 1682952543
transform 1 0 3412 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6870
timestamp 1682952543
transform 1 0 3380 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_6757
timestamp 1682952543
transform 1 0 3492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6867
timestamp 1682952543
transform 1 0 3484 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6868
timestamp 1682952543
transform 1 0 3500 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6897
timestamp 1682952543
transform 1 0 3476 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6871
timestamp 1682952543
transform 1 0 3492 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6775
timestamp 1682952543
transform 1 0 3556 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6758
timestamp 1682952543
transform 1 0 3532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6759
timestamp 1682952543
transform 1 0 3540 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6760
timestamp 1682952543
transform 1 0 3556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6761
timestamp 1682952543
transform 1 0 3572 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6831
timestamp 1682952543
transform 1 0 3532 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6869
timestamp 1682952543
transform 1 0 3540 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6870
timestamp 1682952543
transform 1 0 3548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6871
timestamp 1682952543
transform 1 0 3564 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6898
timestamp 1682952543
transform 1 0 3524 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6919
timestamp 1682952543
transform 1 0 3500 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6920
timestamp 1682952543
transform 1 0 3516 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6832
timestamp 1682952543
transform 1 0 3572 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6872
timestamp 1682952543
transform 1 0 3564 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6899
timestamp 1682952543
transform 1 0 3548 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6921
timestamp 1682952543
transform 1 0 3540 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6732
timestamp 1682952543
transform 1 0 3596 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6776
timestamp 1682952543
transform 1 0 3628 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6762
timestamp 1682952543
transform 1 0 3596 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6809
timestamp 1682952543
transform 1 0 3636 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6810
timestamp 1682952543
transform 1 0 3676 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6872
timestamp 1682952543
transform 1 0 3628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6873
timestamp 1682952543
transform 1 0 3676 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6922
timestamp 1682952543
transform 1 0 3628 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6777
timestamp 1682952543
transform 1 0 3732 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6763
timestamp 1682952543
transform 1 0 3716 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6764
timestamp 1682952543
transform 1 0 3732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6874
timestamp 1682952543
transform 1 0 3708 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6833
timestamp 1682952543
transform 1 0 3716 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6733
timestamp 1682952543
transform 1 0 3748 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_6875
timestamp 1682952543
transform 1 0 3724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6876
timestamp 1682952543
transform 1 0 3740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6877
timestamp 1682952543
transform 1 0 3748 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6778
timestamp 1682952543
transform 1 0 3756 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6900
timestamp 1682952543
transform 1 0 3748 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6923
timestamp 1682952543
transform 1 0 3740 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6779
timestamp 1682952543
transform 1 0 3780 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6765
timestamp 1682952543
transform 1 0 3764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6766
timestamp 1682952543
transform 1 0 3780 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6935
timestamp 1682952543
transform 1 0 3756 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6834
timestamp 1682952543
transform 1 0 3780 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6878
timestamp 1682952543
transform 1 0 3788 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6873
timestamp 1682952543
transform 1 0 3788 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6901
timestamp 1682952543
transform 1 0 3772 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6767
timestamp 1682952543
transform 1 0 3804 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6734
timestamp 1682952543
transform 1 0 3836 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6780
timestamp 1682952543
transform 1 0 3844 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6768
timestamp 1682952543
transform 1 0 3820 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6879
timestamp 1682952543
transform 1 0 3844 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6769
timestamp 1682952543
transform 1 0 3924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6770
timestamp 1682952543
transform 1 0 3932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6771
timestamp 1682952543
transform 1 0 3948 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6772
timestamp 1682952543
transform 1 0 3956 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6773
timestamp 1682952543
transform 1 0 3964 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6880
timestamp 1682952543
transform 1 0 3916 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6835
timestamp 1682952543
transform 1 0 3932 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6881
timestamp 1682952543
transform 1 0 3940 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6874
timestamp 1682952543
transform 1 0 3916 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6902
timestamp 1682952543
transform 1 0 3820 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6903
timestamp 1682952543
transform 1 0 3908 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6936
timestamp 1682952543
transform 1 0 3812 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6904
timestamp 1682952543
transform 1 0 3956 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_6774
timestamp 1682952543
transform 1 0 3980 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6882
timestamp 1682952543
transform 1 0 3972 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6703
timestamp 1682952543
transform 1 0 4004 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6735
timestamp 1682952543
transform 1 0 3996 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6704
timestamp 1682952543
transform 1 0 4084 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6781
timestamp 1682952543
transform 1 0 4020 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6782
timestamp 1682952543
transform 1 0 4060 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_6775
timestamp 1682952543
transform 1 0 4004 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6811
timestamp 1682952543
transform 1 0 4012 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6776
timestamp 1682952543
transform 1 0 4020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6777
timestamp 1682952543
transform 1 0 4036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_6883
timestamp 1682952543
transform 1 0 3996 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6836
timestamp 1682952543
transform 1 0 4004 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_6884
timestamp 1682952543
transform 1 0 4012 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6812
timestamp 1682952543
transform 1 0 4100 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_6885
timestamp 1682952543
transform 1 0 4060 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6886
timestamp 1682952543
transform 1 0 4116 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_6887
timestamp 1682952543
transform 1 0 4124 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6875
timestamp 1682952543
transform 1 0 4020 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6876
timestamp 1682952543
transform 1 0 4068 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6877
timestamp 1682952543
transform 1 0 4116 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6924
timestamp 1682952543
transform 1 0 4036 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6925
timestamp 1682952543
transform 1 0 4068 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_6778
timestamp 1682952543
transform 1 0 4148 0 1 1335
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_56
timestamp 1682952543
transform 1 0 24 0 1 1270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_397
timestamp 1682952543
transform 1 0 72 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_442
timestamp 1682952543
transform -1 0 184 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2760
timestamp 1682952543
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1682952543
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1682952543
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_271
timestamp 1682952543
transform -1 0 248 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2766
timestamp 1682952543
transform 1 0 248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2770
timestamp 1682952543
transform 1 0 256 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1682952543
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1682952543
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_272
timestamp 1682952543
transform 1 0 280 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2773
timestamp 1682952543
transform 1 0 320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1682952543
transform 1 0 328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1682952543
transform 1 0 336 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_275
timestamp 1682952543
transform -1 0 384 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2776
timestamp 1682952543
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1682952543
transform 1 0 392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2782
timestamp 1682952543
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1682952543
transform 1 0 408 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_274
timestamp 1682952543
transform 1 0 416 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2784
timestamp 1682952543
transform 1 0 456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2785
timestamp 1682952543
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_444
timestamp 1682952543
transform 1 0 472 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2786
timestamp 1682952543
transform 1 0 488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1682952543
transform 1 0 496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2788
timestamp 1682952543
transform 1 0 504 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_275
timestamp 1682952543
transform -1 0 552 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2789
timestamp 1682952543
transform 1 0 552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1682952543
transform 1 0 560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1682952543
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1682952543
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2799
timestamp 1682952543
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1682952543
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_276
timestamp 1682952543
transform 1 0 600 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2801
timestamp 1682952543
transform 1 0 640 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1682952543
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1682952543
transform 1 0 656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1682952543
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1682952543
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_84
timestamp 1682952543
transform 1 0 680 0 -1 1370
box -8 -3 32 105
use FILL  FILL_2806
timestamp 1682952543
transform 1 0 704 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_277
timestamp 1682952543
transform 1 0 712 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2807
timestamp 1682952543
transform 1 0 752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1682952543
transform 1 0 760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1682952543
transform 1 0 768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1682952543
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1682952543
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2815
timestamp 1682952543
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_113
timestamp 1682952543
transform 1 0 800 0 -1 1370
box -8 -3 34 105
use FILL  FILL_2818
timestamp 1682952543
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1682952543
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1682952543
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2823
timestamp 1682952543
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1682952543
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1682952543
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1682952543
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_278
timestamp 1682952543
transform 1 0 888 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2827
timestamp 1682952543
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1682952543
transform 1 0 936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2829
timestamp 1682952543
transform 1 0 944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1682952543
transform 1 0 952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1682952543
transform 1 0 960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2834
timestamp 1682952543
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1682952543
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1682952543
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_116
timestamp 1682952543
transform -1 0 1024 0 -1 1370
box -8 -3 34 105
use FILL  FILL_2841
timestamp 1682952543
transform 1 0 1024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1682952543
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1682952543
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1682952543
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2845
timestamp 1682952543
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1682952543
transform 1 0 1064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2847
timestamp 1682952543
transform 1 0 1072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1682952543
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1682952543
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1682952543
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_118
timestamp 1682952543
transform -1 0 1136 0 -1 1370
box -8 -3 34 105
use FILL  FILL_2864
timestamp 1682952543
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_446
timestamp 1682952543
transform -1 0 1160 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2865
timestamp 1682952543
transform 1 0 1160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1682952543
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_403
timestamp 1682952543
transform -1 0 1272 0 -1 1370
box -8 -3 104 105
use FILL  FILL_2867
timestamp 1682952543
transform 1 0 1272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2868
timestamp 1682952543
transform 1 0 1280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2869
timestamp 1682952543
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2870
timestamp 1682952543
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_278
timestamp 1682952543
transform -1 0 1344 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2871
timestamp 1682952543
transform 1 0 1344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1682952543
transform 1 0 1352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1682952543
transform 1 0 1360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2881
timestamp 1682952543
transform 1 0 1368 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_405
timestamp 1682952543
transform 1 0 1376 0 -1 1370
box -8 -3 104 105
use FILL  FILL_2882
timestamp 1682952543
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1682952543
transform 1 0 1480 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_448
timestamp 1682952543
transform 1 0 1488 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2884
timestamp 1682952543
transform 1 0 1504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2885
timestamp 1682952543
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2886
timestamp 1682952543
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_449
timestamp 1682952543
transform -1 0 1544 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2887
timestamp 1682952543
transform 1 0 1544 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1682952543
transform 1 0 1552 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1682952543
transform 1 0 1560 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_452
timestamp 1682952543
transform 1 0 1568 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2892
timestamp 1682952543
transform 1 0 1584 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_407
timestamp 1682952543
transform 1 0 1592 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_453
timestamp 1682952543
transform 1 0 1688 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2894
timestamp 1682952543
transform 1 0 1704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1682952543
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1682952543
transform 1 0 1720 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_280
timestamp 1682952543
transform -1 0 1768 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2901
timestamp 1682952543
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1682952543
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1682952543
transform 1 0 1784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1682952543
transform 1 0 1792 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_454
timestamp 1682952543
transform 1 0 1800 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2907
timestamp 1682952543
transform 1 0 1816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1682952543
transform 1 0 1824 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_281
timestamp 1682952543
transform 1 0 1832 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2914
timestamp 1682952543
transform 1 0 1872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2915
timestamp 1682952543
transform 1 0 1880 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_282
timestamp 1682952543
transform 1 0 1888 0 -1 1370
box -8 -3 46 105
use INVX2  INVX2_460
timestamp 1682952543
transform -1 0 1944 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2916
timestamp 1682952543
transform 1 0 1944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2917
timestamp 1682952543
transform 1 0 1952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1682952543
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1682952543
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_283
timestamp 1682952543
transform 1 0 1976 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2920
timestamp 1682952543
transform 1 0 2016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1682952543
transform 1 0 2024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1682952543
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1682952543
transform 1 0 2040 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_284
timestamp 1682952543
transform -1 0 2088 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2924
timestamp 1682952543
transform 1 0 2088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2925
timestamp 1682952543
transform 1 0 2096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1682952543
transform 1 0 2104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1682952543
transform 1 0 2112 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_285
timestamp 1682952543
transform 1 0 2120 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2928
timestamp 1682952543
transform 1 0 2160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1682952543
transform 1 0 2168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1682952543
transform 1 0 2176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1682952543
transform 1 0 2184 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_287
timestamp 1682952543
transform 1 0 2192 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2936
timestamp 1682952543
transform 1 0 2232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2938
timestamp 1682952543
transform 1 0 2240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1682952543
transform 1 0 2248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2944
timestamp 1682952543
transform 1 0 2256 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_463
timestamp 1682952543
transform -1 0 2280 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2945
timestamp 1682952543
transform 1 0 2280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2946
timestamp 1682952543
transform 1 0 2288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1682952543
transform 1 0 2296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1682952543
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1682952543
transform 1 0 2312 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_288
timestamp 1682952543
transform 1 0 2320 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2950
timestamp 1682952543
transform 1 0 2360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1682952543
transform 1 0 2368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1682952543
transform 1 0 2376 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_464
timestamp 1682952543
transform -1 0 2400 0 -1 1370
box -9 -3 26 105
use FILL  FILL_2953
timestamp 1682952543
transform 1 0 2400 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_411
timestamp 1682952543
transform 1 0 2408 0 -1 1370
box -8 -3 104 105
use FILL  FILL_2960
timestamp 1682952543
transform 1 0 2504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1682952543
transform 1 0 2512 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_292
timestamp 1682952543
transform 1 0 2520 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2973
timestamp 1682952543
transform 1 0 2560 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6937
timestamp 1682952543
transform 1 0 2636 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_413
timestamp 1682952543
transform 1 0 2568 0 -1 1370
box -8 -3 104 105
use M3_M2  M3_M2_6938
timestamp 1682952543
transform 1 0 2716 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_414
timestamp 1682952543
transform 1 0 2664 0 -1 1370
box -8 -3 104 105
use FILL  FILL_2974
timestamp 1682952543
transform 1 0 2760 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_293
timestamp 1682952543
transform 1 0 2768 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2975
timestamp 1682952543
transform 1 0 2808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1682952543
transform 1 0 2816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1682952543
transform 1 0 2824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2980
timestamp 1682952543
transform 1 0 2832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1682952543
transform 1 0 2840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2984
timestamp 1682952543
transform 1 0 2848 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_279
timestamp 1682952543
transform 1 0 2856 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2990
timestamp 1682952543
transform 1 0 2896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1682952543
transform 1 0 2904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1682952543
transform 1 0 2912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1682952543
transform 1 0 2920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1682952543
transform 1 0 2928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1682952543
transform 1 0 2936 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_295
timestamp 1682952543
transform 1 0 2944 0 -1 1370
box -8 -3 46 105
use FILL  FILL_2996
timestamp 1682952543
transform 1 0 2984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1682952543
transform 1 0 2992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1682952543
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1682952543
transform 1 0 3008 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_296
timestamp 1682952543
transform 1 0 3016 0 -1 1370
box -8 -3 46 105
use AOI22X1  AOI22X1_280
timestamp 1682952543
transform -1 0 3096 0 -1 1370
box -8 -3 46 105
use FILL  FILL_3000
timestamp 1682952543
transform 1 0 3096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1682952543
transform 1 0 3104 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_281
timestamp 1682952543
transform 1 0 3112 0 -1 1370
box -8 -3 46 105
use FILL  FILL_3002
timestamp 1682952543
transform 1 0 3152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1682952543
transform 1 0 3160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1682952543
transform 1 0 3168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1682952543
transform 1 0 3176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1682952543
transform 1 0 3184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1682952543
transform 1 0 3192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1682952543
transform 1 0 3200 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_417
timestamp 1682952543
transform 1 0 3208 0 -1 1370
box -8 -3 104 105
use FILL  FILL_3019
timestamp 1682952543
transform 1 0 3304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1682952543
transform 1 0 3312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1682952543
transform 1 0 3320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1682952543
transform 1 0 3328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1682952543
transform 1 0 3336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1682952543
transform 1 0 3344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1682952543
transform 1 0 3352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3037
timestamp 1682952543
transform 1 0 3360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3038
timestamp 1682952543
transform 1 0 3368 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_419
timestamp 1682952543
transform -1 0 3472 0 -1 1370
box -8 -3 104 105
use FILL  FILL_3039
timestamp 1682952543
transform 1 0 3472 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_282
timestamp 1682952543
transform 1 0 3480 0 -1 1370
box -8 -3 46 105
use FILL  FILL_3040
timestamp 1682952543
transform 1 0 3520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1682952543
transform 1 0 3528 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_300
timestamp 1682952543
transform 1 0 3536 0 -1 1370
box -8 -3 46 105
use FILL  FILL_3042
timestamp 1682952543
transform 1 0 3576 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_420
timestamp 1682952543
transform 1 0 3584 0 -1 1370
box -8 -3 104 105
use FILL  FILL_3043
timestamp 1682952543
transform 1 0 3680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3044
timestamp 1682952543
transform 1 0 3688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1682952543
transform 1 0 3696 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_286
timestamp 1682952543
transform 1 0 3704 0 -1 1370
box -8 -3 46 105
use FILL  FILL_3060
timestamp 1682952543
transform 1 0 3744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1682952543
transform 1 0 3752 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_302
timestamp 1682952543
transform 1 0 3760 0 -1 1370
box -8 -3 46 105
use FILL  FILL_3062
timestamp 1682952543
transform 1 0 3800 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_421
timestamp 1682952543
transform 1 0 3808 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_477
timestamp 1682952543
transform 1 0 3904 0 -1 1370
box -9 -3 26 105
use AOI22X1  AOI22X1_287
timestamp 1682952543
transform 1 0 3920 0 -1 1370
box -8 -3 46 105
use INVX2  INVX2_478
timestamp 1682952543
transform 1 0 3960 0 -1 1370
box -9 -3 26 105
use FILL  FILL_3063
timestamp 1682952543
transform 1 0 3976 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_304
timestamp 1682952543
transform 1 0 3984 0 -1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_422
timestamp 1682952543
transform 1 0 4024 0 -1 1370
box -8 -3 104 105
use INVX2  INVX2_480
timestamp 1682952543
transform -1 0 4136 0 -1 1370
box -9 -3 26 105
use FILL  FILL_3077
timestamp 1682952543
transform 1 0 4136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1682952543
transform 1 0 4144 0 -1 1370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_57
timestamp 1682952543
transform 1 0 4201 0 1 1270
box -10 -3 10 3
use M3_M2  M3_M2_6969
timestamp 1682952543
transform 1 0 100 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_7009
timestamp 1682952543
transform 1 0 92 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6896
timestamp 1682952543
transform 1 0 108 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_6900
timestamp 1682952543
transform 1 0 100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6999
timestamp 1682952543
transform 1 0 92 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7010
timestamp 1682952543
transform 1 0 140 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6901
timestamp 1682952543
transform 1 0 140 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7000
timestamp 1682952543
transform 1 0 132 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7083
timestamp 1682952543
transform 1 0 140 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6948
timestamp 1682952543
transform 1 0 172 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_6902
timestamp 1682952543
transform 1 0 172 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7084
timestamp 1682952543
transform 1 0 164 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7001
timestamp 1682952543
transform 1 0 172 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7104
timestamp 1682952543
transform 1 0 172 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6970
timestamp 1682952543
transform 1 0 196 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_7011
timestamp 1682952543
transform 1 0 188 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7002
timestamp 1682952543
transform 1 0 188 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6985
timestamp 1682952543
transform 1 0 212 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6949
timestamp 1682952543
transform 1 0 252 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6971
timestamp 1682952543
transform 1 0 244 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_7012
timestamp 1682952543
transform 1 0 228 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6903
timestamp 1682952543
transform 1 0 212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6904
timestamp 1682952543
transform 1 0 228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6905
timestamp 1682952543
transform 1 0 244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7003
timestamp 1682952543
transform 1 0 212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7004
timestamp 1682952543
transform 1 0 220 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7105
timestamp 1682952543
transform 1 0 220 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7005
timestamp 1682952543
transform 1 0 260 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7106
timestamp 1682952543
transform 1 0 260 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6950
timestamp 1682952543
transform 1 0 276 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7013
timestamp 1682952543
transform 1 0 284 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7014
timestamp 1682952543
transform 1 0 324 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7054
timestamp 1682952543
transform 1 0 276 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6906
timestamp 1682952543
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7055
timestamp 1682952543
transform 1 0 300 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6972
timestamp 1682952543
transform 1 0 396 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6986
timestamp 1682952543
transform 1 0 388 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6907
timestamp 1682952543
transform 1 0 324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6908
timestamp 1682952543
transform 1 0 380 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7006
timestamp 1682952543
transform 1 0 276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7007
timestamp 1682952543
transform 1 0 300 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7085
timestamp 1682952543
transform 1 0 348 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7150
timestamp 1682952543
transform 1 0 300 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7056
timestamp 1682952543
transform 1 0 388 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6973
timestamp 1682952543
transform 1 0 436 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_7015
timestamp 1682952543
transform 1 0 404 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7016
timestamp 1682952543
transform 1 0 444 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6909
timestamp 1682952543
transform 1 0 404 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7057
timestamp 1682952543
transform 1 0 420 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6910
timestamp 1682952543
transform 1 0 444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6911
timestamp 1682952543
transform 1 0 500 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7008
timestamp 1682952543
transform 1 0 396 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7151
timestamp 1682952543
transform 1 0 388 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7009
timestamp 1682952543
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7152
timestamp 1682952543
transform 1 0 420 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7153
timestamp 1682952543
transform 1 0 508 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_6912
timestamp 1682952543
transform 1 0 524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6913
timestamp 1682952543
transform 1 0 540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7010
timestamp 1682952543
transform 1 0 532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7011
timestamp 1682952543
transform 1 0 548 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7107
timestamp 1682952543
transform 1 0 548 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7154
timestamp 1682952543
transform 1 0 532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6951
timestamp 1682952543
transform 1 0 580 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7058
timestamp 1682952543
transform 1 0 580 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_7086
timestamp 1682952543
transform 1 0 572 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7012
timestamp 1682952543
transform 1 0 580 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7017
timestamp 1682952543
transform 1 0 604 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6914
timestamp 1682952543
transform 1 0 604 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7087
timestamp 1682952543
transform 1 0 604 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6939
timestamp 1682952543
transform 1 0 660 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_7018
timestamp 1682952543
transform 1 0 644 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7019
timestamp 1682952543
transform 1 0 684 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7020
timestamp 1682952543
transform 1 0 700 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7059
timestamp 1682952543
transform 1 0 620 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6915
timestamp 1682952543
transform 1 0 644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6916
timestamp 1682952543
transform 1 0 700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6917
timestamp 1682952543
transform 1 0 708 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7013
timestamp 1682952543
transform 1 0 620 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7108
timestamp 1682952543
transform 1 0 620 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7109
timestamp 1682952543
transform 1 0 668 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7014
timestamp 1682952543
transform 1 0 732 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6952
timestamp 1682952543
transform 1 0 876 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7021
timestamp 1682952543
transform 1 0 828 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7022
timestamp 1682952543
transform 1 0 868 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6918
timestamp 1682952543
transform 1 0 828 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7060
timestamp 1682952543
transform 1 0 852 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6919
timestamp 1682952543
transform 1 0 860 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6920
timestamp 1682952543
transform 1 0 868 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7015
timestamp 1682952543
transform 1 0 780 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7088
timestamp 1682952543
transform 1 0 844 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7110
timestamp 1682952543
transform 1 0 780 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7111
timestamp 1682952543
transform 1 0 860 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7092
timestamp 1682952543
transform 1 0 892 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_7155
timestamp 1682952543
transform 1 0 892 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_6921
timestamp 1682952543
transform 1 0 908 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7061
timestamp 1682952543
transform 1 0 916 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_7089
timestamp 1682952543
transform 1 0 908 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7062
timestamp 1682952543
transform 1 0 932 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7016
timestamp 1682952543
transform 1 0 924 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7017
timestamp 1682952543
transform 1 0 932 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7112
timestamp 1682952543
transform 1 0 948 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7023
timestamp 1682952543
transform 1 0 988 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6922
timestamp 1682952543
transform 1 0 980 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7113
timestamp 1682952543
transform 1 0 980 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7156
timestamp 1682952543
transform 1 0 980 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_6923
timestamp 1682952543
transform 1 0 996 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7018
timestamp 1682952543
transform 1 0 1012 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7114
timestamp 1682952543
transform 1 0 1012 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7157
timestamp 1682952543
transform 1 0 996 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_6897
timestamp 1682952543
transform 1 0 1068 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_7024
timestamp 1682952543
transform 1 0 1076 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7063
timestamp 1682952543
transform 1 0 1068 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7019
timestamp 1682952543
transform 1 0 1076 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7115
timestamp 1682952543
transform 1 0 1076 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6974
timestamp 1682952543
transform 1 0 1092 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_6898
timestamp 1682952543
transform 1 0 1108 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_6924
timestamp 1682952543
transform 1 0 1092 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7064
timestamp 1682952543
transform 1 0 1100 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_7025
timestamp 1682952543
transform 1 0 1132 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6925
timestamp 1682952543
transform 1 0 1124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7020
timestamp 1682952543
transform 1 0 1100 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7116
timestamp 1682952543
transform 1 0 1100 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_6926
timestamp 1682952543
transform 1 0 1140 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7117
timestamp 1682952543
transform 1 0 1132 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7090
timestamp 1682952543
transform 1 0 1148 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6940
timestamp 1682952543
transform 1 0 1188 0 1 1265
box -3 -3 3 3
use M2_M1  M2_M1_7021
timestamp 1682952543
transform 1 0 1172 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7022
timestamp 1682952543
transform 1 0 1180 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7158
timestamp 1682952543
transform 1 0 1172 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6975
timestamp 1682952543
transform 1 0 1228 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_7026
timestamp 1682952543
transform 1 0 1204 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6927
timestamp 1682952543
transform 1 0 1188 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7065
timestamp 1682952543
transform 1 0 1196 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6928
timestamp 1682952543
transform 1 0 1204 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7023
timestamp 1682952543
transform 1 0 1196 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7091
timestamp 1682952543
transform 1 0 1204 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7027
timestamp 1682952543
transform 1 0 1244 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7066
timestamp 1682952543
transform 1 0 1236 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6929
timestamp 1682952543
transform 1 0 1244 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7024
timestamp 1682952543
transform 1 0 1212 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7025
timestamp 1682952543
transform 1 0 1228 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7026
timestamp 1682952543
transform 1 0 1236 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7118
timestamp 1682952543
transform 1 0 1220 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7159
timestamp 1682952543
transform 1 0 1220 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6987
timestamp 1682952543
transform 1 0 1260 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7067
timestamp 1682952543
transform 1 0 1276 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7027
timestamp 1682952543
transform 1 0 1276 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7160
timestamp 1682952543
transform 1 0 1284 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6988
timestamp 1682952543
transform 1 0 1300 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7028
timestamp 1682952543
transform 1 0 1316 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6930
timestamp 1682952543
transform 1 0 1300 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6931
timestamp 1682952543
transform 1 0 1316 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7029
timestamp 1682952543
transform 1 0 1332 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7068
timestamp 1682952543
transform 1 0 1332 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7028
timestamp 1682952543
transform 1 0 1308 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7029
timestamp 1682952543
transform 1 0 1324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7030
timestamp 1682952543
transform 1 0 1332 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7119
timestamp 1682952543
transform 1 0 1324 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7092
timestamp 1682952543
transform 1 0 1372 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6976
timestamp 1682952543
transform 1 0 1404 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_7030
timestamp 1682952543
transform 1 0 1428 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6932
timestamp 1682952543
transform 1 0 1404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6933
timestamp 1682952543
transform 1 0 1428 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7093
timestamp 1682952543
transform 1 0 1404 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7031
timestamp 1682952543
transform 1 0 1412 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7161
timestamp 1682952543
transform 1 0 1404 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6953
timestamp 1682952543
transform 1 0 1460 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7031
timestamp 1682952543
transform 1 0 1452 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6934
timestamp 1682952543
transform 1 0 1444 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7120
timestamp 1682952543
transform 1 0 1444 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_6935
timestamp 1682952543
transform 1 0 1460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7032
timestamp 1682952543
transform 1 0 1460 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6977
timestamp 1682952543
transform 1 0 1468 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6978
timestamp 1682952543
transform 1 0 1484 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6989
timestamp 1682952543
transform 1 0 1476 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7033
timestamp 1682952543
transform 1 0 1476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_6936
timestamp 1682952543
transform 1 0 1492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6937
timestamp 1682952543
transform 1 0 1524 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7121
timestamp 1682952543
transform 1 0 1532 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7034
timestamp 1682952543
transform 1 0 1548 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6941
timestamp 1682952543
transform 1 0 1644 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_7069
timestamp 1682952543
transform 1 0 1580 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_7070
timestamp 1682952543
transform 1 0 1604 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6938
timestamp 1682952543
transform 1 0 1620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7035
timestamp 1682952543
transform 1 0 1564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7036
timestamp 1682952543
transform 1 0 1580 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7094
timestamp 1682952543
transform 1 0 1620 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7122
timestamp 1682952543
transform 1 0 1612 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7032
timestamp 1682952543
transform 1 0 1676 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7071
timestamp 1682952543
transform 1 0 1668 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6939
timestamp 1682952543
transform 1 0 1684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6940
timestamp 1682952543
transform 1 0 1692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7037
timestamp 1682952543
transform 1 0 1676 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7072
timestamp 1682952543
transform 1 0 1700 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6941
timestamp 1682952543
transform 1 0 1708 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7095
timestamp 1682952543
transform 1 0 1692 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7038
timestamp 1682952543
transform 1 0 1700 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7123
timestamp 1682952543
transform 1 0 1692 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7039
timestamp 1682952543
transform 1 0 1732 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7124
timestamp 1682952543
transform 1 0 1724 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_6942
timestamp 1682952543
transform 1 0 1756 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7073
timestamp 1682952543
transform 1 0 1764 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6943
timestamp 1682952543
transform 1 0 1772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7040
timestamp 1682952543
transform 1 0 1764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7041
timestamp 1682952543
transform 1 0 1780 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6990
timestamp 1682952543
transform 1 0 1828 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6991
timestamp 1682952543
transform 1 0 1852 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6992
timestamp 1682952543
transform 1 0 1892 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6944
timestamp 1682952543
transform 1 0 1796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6945
timestamp 1682952543
transform 1 0 1844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7042
timestamp 1682952543
transform 1 0 1876 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7125
timestamp 1682952543
transform 1 0 1860 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7126
timestamp 1682952543
transform 1 0 1876 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_6946
timestamp 1682952543
transform 1 0 1924 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7074
timestamp 1682952543
transform 1 0 1948 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6947
timestamp 1682952543
transform 1 0 1980 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7043
timestamp 1682952543
transform 1 0 1900 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7127
timestamp 1682952543
transform 1 0 1900 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7128
timestamp 1682952543
transform 1 0 1924 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7129
timestamp 1682952543
transform 1 0 1948 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_6948
timestamp 1682952543
transform 1 0 2004 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7044
timestamp 1682952543
transform 1 0 2028 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7045
timestamp 1682952543
transform 1 0 2060 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7162
timestamp 1682952543
transform 1 0 2060 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6993
timestamp 1682952543
transform 1 0 2092 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7033
timestamp 1682952543
transform 1 0 2084 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6949
timestamp 1682952543
transform 1 0 2076 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6950
timestamp 1682952543
transform 1 0 2092 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7046
timestamp 1682952543
transform 1 0 2084 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6954
timestamp 1682952543
transform 1 0 2124 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6955
timestamp 1682952543
transform 1 0 2172 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7047
timestamp 1682952543
transform 1 0 2116 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7130
timestamp 1682952543
transform 1 0 2116 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6979
timestamp 1682952543
transform 1 0 2132 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6980
timestamp 1682952543
transform 1 0 2196 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6942
timestamp 1682952543
transform 1 0 2268 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6956
timestamp 1682952543
transform 1 0 2316 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6981
timestamp 1682952543
transform 1 0 2268 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6994
timestamp 1682952543
transform 1 0 2228 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7034
timestamp 1682952543
transform 1 0 2156 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7035
timestamp 1682952543
transform 1 0 2212 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7075
timestamp 1682952543
transform 1 0 2132 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6951
timestamp 1682952543
transform 1 0 2156 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7048
timestamp 1682952543
transform 1 0 2132 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7131
timestamp 1682952543
transform 1 0 2164 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7132
timestamp 1682952543
transform 1 0 2196 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7163
timestamp 1682952543
transform 1 0 2148 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7164
timestamp 1682952543
transform 1 0 2180 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7036
timestamp 1682952543
transform 1 0 2268 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6957
timestamp 1682952543
transform 1 0 2396 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6995
timestamp 1682952543
transform 1 0 2372 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7037
timestamp 1682952543
transform 1 0 2340 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7038
timestamp 1682952543
transform 1 0 2364 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6952
timestamp 1682952543
transform 1 0 2228 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6953
timestamp 1682952543
transform 1 0 2268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6954
timestamp 1682952543
transform 1 0 2324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6955
timestamp 1682952543
transform 1 0 2364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6956
timestamp 1682952543
transform 1 0 2420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7049
timestamp 1682952543
transform 1 0 2244 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7133
timestamp 1682952543
transform 1 0 2228 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7050
timestamp 1682952543
transform 1 0 2340 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7165
timestamp 1682952543
transform 1 0 2372 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6958
timestamp 1682952543
transform 1 0 2444 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6996
timestamp 1682952543
transform 1 0 2436 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6957
timestamp 1682952543
transform 1 0 2436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6958
timestamp 1682952543
transform 1 0 2460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7051
timestamp 1682952543
transform 1 0 2428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7052
timestamp 1682952543
transform 1 0 2452 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7134
timestamp 1682952543
transform 1 0 2436 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7166
timestamp 1682952543
transform 1 0 2428 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_6899
timestamp 1682952543
transform 1 0 2476 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_7167
timestamp 1682952543
transform 1 0 2444 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7168
timestamp 1682952543
transform 1 0 2468 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_6959
timestamp 1682952543
transform 1 0 2484 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6959
timestamp 1682952543
transform 1 0 2524 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7053
timestamp 1682952543
transform 1 0 2516 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6997
timestamp 1682952543
transform 1 0 2596 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6960
timestamp 1682952543
transform 1 0 2556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7054
timestamp 1682952543
transform 1 0 2532 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7135
timestamp 1682952543
transform 1 0 2532 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7136
timestamp 1682952543
transform 1 0 2580 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7169
timestamp 1682952543
transform 1 0 2532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7170
timestamp 1682952543
transform 1 0 2572 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6960
timestamp 1682952543
transform 1 0 2692 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6982
timestamp 1682952543
transform 1 0 2652 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6998
timestamp 1682952543
transform 1 0 2644 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6961
timestamp 1682952543
transform 1 0 2628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6962
timestamp 1682952543
transform 1 0 2700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7055
timestamp 1682952543
transform 1 0 2652 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7137
timestamp 1682952543
transform 1 0 2700 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6999
timestamp 1682952543
transform 1 0 2788 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7039
timestamp 1682952543
transform 1 0 2780 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7040
timestamp 1682952543
transform 1 0 2804 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6963
timestamp 1682952543
transform 1 0 2780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6964
timestamp 1682952543
transform 1 0 2788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6965
timestamp 1682952543
transform 1 0 2804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7056
timestamp 1682952543
transform 1 0 2780 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7057
timestamp 1682952543
transform 1 0 2796 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7058
timestamp 1682952543
transform 1 0 2812 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7059
timestamp 1682952543
transform 1 0 2820 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7138
timestamp 1682952543
transform 1 0 2796 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7139
timestamp 1682952543
transform 1 0 2812 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_6966
timestamp 1682952543
transform 1 0 2844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7060
timestamp 1682952543
transform 1 0 2844 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7041
timestamp 1682952543
transform 1 0 2884 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6967
timestamp 1682952543
transform 1 0 2860 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7076
timestamp 1682952543
transform 1 0 2868 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6968
timestamp 1682952543
transform 1 0 2876 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6969
timestamp 1682952543
transform 1 0 2892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7061
timestamp 1682952543
transform 1 0 2868 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7062
timestamp 1682952543
transform 1 0 2884 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7063
timestamp 1682952543
transform 1 0 2892 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7096
timestamp 1682952543
transform 1 0 2908 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6943
timestamp 1682952543
transform 1 0 3012 0 1 1265
box -3 -3 3 3
use M2_M1  M2_M1_6970
timestamp 1682952543
transform 1 0 2964 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7077
timestamp 1682952543
transform 1 0 2972 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_7078
timestamp 1682952543
transform 1 0 3004 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6971
timestamp 1682952543
transform 1 0 3020 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7064
timestamp 1682952543
transform 1 0 2940 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7097
timestamp 1682952543
transform 1 0 3012 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6961
timestamp 1682952543
transform 1 0 3116 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6983
timestamp 1682952543
transform 1 0 3148 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_6972
timestamp 1682952543
transform 1 0 3068 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6973
timestamp 1682952543
transform 1 0 3124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7065
timestamp 1682952543
transform 1 0 3148 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7140
timestamp 1682952543
transform 1 0 3116 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7171
timestamp 1682952543
transform 1 0 3116 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7000
timestamp 1682952543
transform 1 0 3164 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6974
timestamp 1682952543
transform 1 0 3164 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7172
timestamp 1682952543
transform 1 0 3172 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7001
timestamp 1682952543
transform 1 0 3196 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7042
timestamp 1682952543
transform 1 0 3212 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6975
timestamp 1682952543
transform 1 0 3212 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7066
timestamp 1682952543
transform 1 0 3188 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7067
timestamp 1682952543
transform 1 0 3204 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7098
timestamp 1682952543
transform 1 0 3212 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7068
timestamp 1682952543
transform 1 0 3220 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7141
timestamp 1682952543
transform 1 0 3188 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7173
timestamp 1682952543
transform 1 0 3220 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6944
timestamp 1682952543
transform 1 0 3236 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_7142
timestamp 1682952543
transform 1 0 3236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6945
timestamp 1682952543
transform 1 0 3268 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6962
timestamp 1682952543
transform 1 0 3300 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7079
timestamp 1682952543
transform 1 0 3260 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6976
timestamp 1682952543
transform 1 0 3284 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7080
timestamp 1682952543
transform 1 0 3308 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7069
timestamp 1682952543
transform 1 0 3260 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7099
timestamp 1682952543
transform 1 0 3284 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7143
timestamp 1682952543
transform 1 0 3276 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7002
timestamp 1682952543
transform 1 0 3372 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7043
timestamp 1682952543
transform 1 0 3356 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6977
timestamp 1682952543
transform 1 0 3356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6978
timestamp 1682952543
transform 1 0 3364 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6963
timestamp 1682952543
transform 1 0 3420 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7044
timestamp 1682952543
transform 1 0 3404 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6979
timestamp 1682952543
transform 1 0 3372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6980
timestamp 1682952543
transform 1 0 3404 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6984
timestamp 1682952543
transform 1 0 3428 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_6981
timestamp 1682952543
transform 1 0 3452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7070
timestamp 1682952543
transform 1 0 3372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7071
timestamp 1682952543
transform 1 0 3380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7072
timestamp 1682952543
transform 1 0 3396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7073
timestamp 1682952543
transform 1 0 3412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7074
timestamp 1682952543
transform 1 0 3428 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7144
timestamp 1682952543
transform 1 0 3396 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7174
timestamp 1682952543
transform 1 0 3404 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7145
timestamp 1682952543
transform 1 0 3452 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6964
timestamp 1682952543
transform 1 0 3516 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7003
timestamp 1682952543
transform 1 0 3548 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7045
timestamp 1682952543
transform 1 0 3540 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_7046
timestamp 1682952543
transform 1 0 3572 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6982
timestamp 1682952543
transform 1 0 3540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6983
timestamp 1682952543
transform 1 0 3548 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6984
timestamp 1682952543
transform 1 0 3572 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7047
timestamp 1682952543
transform 1 0 3588 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6985
timestamp 1682952543
transform 1 0 3588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7075
timestamp 1682952543
transform 1 0 3548 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7076
timestamp 1682952543
transform 1 0 3564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7077
timestamp 1682952543
transform 1 0 3580 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7175
timestamp 1682952543
transform 1 0 3580 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7004
timestamp 1682952543
transform 1 0 3644 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6986
timestamp 1682952543
transform 1 0 3644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7078
timestamp 1682952543
transform 1 0 3636 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7048
timestamp 1682952543
transform 1 0 3684 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6987
timestamp 1682952543
transform 1 0 3684 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7079
timestamp 1682952543
transform 1 0 3660 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7080
timestamp 1682952543
transform 1 0 3676 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7100
timestamp 1682952543
transform 1 0 3684 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7049
timestamp 1682952543
transform 1 0 3700 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6988
timestamp 1682952543
transform 1 0 3700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7081
timestamp 1682952543
transform 1 0 3692 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7101
timestamp 1682952543
transform 1 0 3700 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7176
timestamp 1682952543
transform 1 0 3692 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7005
timestamp 1682952543
transform 1 0 3748 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_7050
timestamp 1682952543
transform 1 0 3732 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6989
timestamp 1682952543
transform 1 0 3732 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6990
timestamp 1682952543
transform 1 0 3748 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6946
timestamp 1682952543
transform 1 0 3804 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_7006
timestamp 1682952543
transform 1 0 3844 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6991
timestamp 1682952543
transform 1 0 3796 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7082
timestamp 1682952543
transform 1 0 3716 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7083
timestamp 1682952543
transform 1 0 3724 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7084
timestamp 1682952543
transform 1 0 3740 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7085
timestamp 1682952543
transform 1 0 3756 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7086
timestamp 1682952543
transform 1 0 3772 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7146
timestamp 1682952543
transform 1 0 3740 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7177
timestamp 1682952543
transform 1 0 3724 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7147
timestamp 1682952543
transform 1 0 3796 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6965
timestamp 1682952543
transform 1 0 3892 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7051
timestamp 1682952543
transform 1 0 3868 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6947
timestamp 1682952543
transform 1 0 3980 0 1 1265
box -3 -3 3 3
use M3_M2  M3_M2_6966
timestamp 1682952543
transform 1 0 3980 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7007
timestamp 1682952543
transform 1 0 3972 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6992
timestamp 1682952543
transform 1 0 3868 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7081
timestamp 1682952543
transform 1 0 3884 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_7082
timestamp 1682952543
transform 1 0 3924 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_6993
timestamp 1682952543
transform 1 0 3932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7087
timestamp 1682952543
transform 1 0 3884 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7148
timestamp 1682952543
transform 1 0 3932 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7052
timestamp 1682952543
transform 1 0 3980 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6994
timestamp 1682952543
transform 1 0 3980 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_7102
timestamp 1682952543
transform 1 0 3980 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_7178
timestamp 1682952543
transform 1 0 3868 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7179
timestamp 1682952543
transform 1 0 3916 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7180
timestamp 1682952543
transform 1 0 3964 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_7008
timestamp 1682952543
transform 1 0 3996 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_6995
timestamp 1682952543
transform 1 0 3996 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6967
timestamp 1682952543
transform 1 0 4012 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_7053
timestamp 1682952543
transform 1 0 4028 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_6996
timestamp 1682952543
transform 1 0 4028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7088
timestamp 1682952543
transform 1 0 4004 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7103
timestamp 1682952543
transform 1 0 4012 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7089
timestamp 1682952543
transform 1 0 4020 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7090
timestamp 1682952543
transform 1 0 4036 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_7149
timestamp 1682952543
transform 1 0 4020 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_7181
timestamp 1682952543
transform 1 0 4036 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6968
timestamp 1682952543
transform 1 0 4076 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_6997
timestamp 1682952543
transform 1 0 4100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_6998
timestamp 1682952543
transform 1 0 4148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7091
timestamp 1682952543
transform 1 0 4068 0 1 1205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_58
timestamp 1682952543
transform 1 0 48 0 1 1170
box -10 -3 10 3
use FILL  FILL_3080
timestamp 1682952543
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1682952543
transform 1 0 80 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_481
timestamp 1682952543
transform 1 0 88 0 1 1170
box -9 -3 26 105
use FILL  FILL_3082
timestamp 1682952543
transform 1 0 104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1682952543
transform 1 0 112 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_288
timestamp 1682952543
transform -1 0 160 0 1 1170
box -8 -3 46 105
use FILL  FILL_3084
timestamp 1682952543
transform 1 0 160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3085
timestamp 1682952543
transform 1 0 168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1682952543
transform 1 0 176 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_482
timestamp 1682952543
transform 1 0 184 0 1 1170
box -9 -3 26 105
use FILL  FILL_3087
timestamp 1682952543
transform 1 0 200 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_289
timestamp 1682952543
transform 1 0 208 0 1 1170
box -8 -3 46 105
use FILL  FILL_3088
timestamp 1682952543
transform 1 0 248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1682952543
transform 1 0 256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1682952543
transform 1 0 264 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_483
timestamp 1682952543
transform 1 0 272 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_423
timestamp 1682952543
transform 1 0 288 0 1 1170
box -8 -3 104 105
use FILL  FILL_3091
timestamp 1682952543
transform 1 0 384 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_484
timestamp 1682952543
transform 1 0 392 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_424
timestamp 1682952543
transform 1 0 408 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_7182
timestamp 1682952543
transform 1 0 516 0 1 1175
box -3 -3 3 3
use FILL  FILL_3092
timestamp 1682952543
transform 1 0 504 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7183
timestamp 1682952543
transform 1 0 548 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_305
timestamp 1682952543
transform 1 0 512 0 1 1170
box -8 -3 46 105
use FILL  FILL_3093
timestamp 1682952543
transform 1 0 552 0 1 1170
box -8 -3 16 105
use FILL  FILL_3098
timestamp 1682952543
transform 1 0 560 0 1 1170
box -8 -3 16 105
use FILL  FILL_3100
timestamp 1682952543
transform 1 0 568 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_487
timestamp 1682952543
transform 1 0 576 0 1 1170
box -9 -3 26 105
use FILL  FILL_3102
timestamp 1682952543
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1682952543
transform 1 0 600 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7184
timestamp 1682952543
transform 1 0 636 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_7185
timestamp 1682952543
transform 1 0 660 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_429
timestamp 1682952543
transform 1 0 608 0 1 1170
box -8 -3 104 105
use FILL  FILL_3104
timestamp 1682952543
transform 1 0 704 0 1 1170
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1682952543
transform 1 0 712 0 1 1170
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1682952543
transform 1 0 720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1682952543
transform 1 0 728 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_488
timestamp 1682952543
transform 1 0 736 0 1 1170
box -9 -3 26 105
use FILL  FILL_3108
timestamp 1682952543
transform 1 0 752 0 1 1170
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1682952543
transform 1 0 760 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_430
timestamp 1682952543
transform 1 0 768 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_489
timestamp 1682952543
transform -1 0 880 0 1 1170
box -9 -3 26 105
use FILL  FILL_3110
timestamp 1682952543
transform 1 0 880 0 1 1170
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1682952543
transform 1 0 888 0 1 1170
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1682952543
transform 1 0 896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1682952543
transform 1 0 904 0 1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_86
timestamp 1682952543
transform 1 0 912 0 1 1170
box -8 -3 32 105
use FILL  FILL_3114
timestamp 1682952543
transform 1 0 936 0 1 1170
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1682952543
transform 1 0 944 0 1 1170
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1682952543
transform 1 0 952 0 1 1170
box -8 -3 16 105
use FILL  FILL_3117
timestamp 1682952543
transform 1 0 960 0 1 1170
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1682952543
transform 1 0 968 0 1 1170
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1682952543
transform 1 0 976 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_122
timestamp 1682952543
transform 1 0 984 0 1 1170
box -8 -3 34 105
use FILL  FILL_3120
timestamp 1682952543
transform 1 0 1016 0 1 1170
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1682952543
transform 1 0 1024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1682952543
transform 1 0 1032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1682952543
transform 1 0 1040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3126
timestamp 1682952543
transform 1 0 1048 0 1 1170
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1682952543
transform 1 0 1056 0 1 1170
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1682952543
transform 1 0 1064 0 1 1170
box -8 -3 16 105
use BUFX2  BUFX2_96
timestamp 1682952543
transform -1 0 1096 0 1 1170
box -5 -3 28 105
use FILL  FILL_3129
timestamp 1682952543
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_123
timestamp 1682952543
transform -1 0 1136 0 1 1170
box -8 -3 34 105
use FILL  FILL_3130
timestamp 1682952543
transform 1 0 1136 0 1 1170
box -8 -3 16 105
use FILL  FILL_3131
timestamp 1682952543
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1682952543
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1682952543
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3134
timestamp 1682952543
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_490
timestamp 1682952543
transform 1 0 1176 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_7186
timestamp 1682952543
transform 1 0 1228 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_307
timestamp 1682952543
transform -1 0 1232 0 1 1170
box -8 -3 46 105
use FILL  FILL_3135
timestamp 1682952543
transform 1 0 1232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1682952543
transform 1 0 1240 0 1 1170
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1682952543
transform 1 0 1248 0 1 1170
box -8 -3 16 105
use FILL  FILL_3141
timestamp 1682952543
transform 1 0 1256 0 1 1170
box -8 -3 16 105
use FILL  FILL_3142
timestamp 1682952543
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1682952543
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1682952543
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_308
timestamp 1682952543
transform -1 0 1328 0 1 1170
box -8 -3 46 105
use FILL  FILL_3145
timestamp 1682952543
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1682952543
transform 1 0 1336 0 1 1170
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1682952543
transform 1 0 1344 0 1 1170
box -8 -3 16 105
use FILL  FILL_3150
timestamp 1682952543
transform 1 0 1352 0 1 1170
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1682952543
transform 1 0 1360 0 1 1170
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1682952543
transform 1 0 1368 0 1 1170
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1682952543
transform 1 0 1376 0 1 1170
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1682952543
transform 1 0 1384 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_309
timestamp 1682952543
transform -1 0 1432 0 1 1170
box -8 -3 46 105
use FILL  FILL_3156
timestamp 1682952543
transform 1 0 1432 0 1 1170
box -8 -3 16 105
use FILL  FILL_3157
timestamp 1682952543
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use FILL  FILL_3158
timestamp 1682952543
transform 1 0 1448 0 1 1170
box -8 -3 16 105
use FILL  FILL_3159
timestamp 1682952543
transform 1 0 1456 0 1 1170
box -8 -3 16 105
use FILL  FILL_3160
timestamp 1682952543
transform 1 0 1464 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7187
timestamp 1682952543
transform 1 0 1492 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_492
timestamp 1682952543
transform 1 0 1472 0 1 1170
box -9 -3 26 105
use FILL  FILL_3161
timestamp 1682952543
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1682952543
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_493
timestamp 1682952543
transform -1 0 1520 0 1 1170
box -9 -3 26 105
use FILL  FILL_3163
timestamp 1682952543
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1682952543
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_3165
timestamp 1682952543
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1682952543
transform 1 0 1544 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_494
timestamp 1682952543
transform -1 0 1568 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_437
timestamp 1682952543
transform 1 0 1568 0 1 1170
box -8 -3 104 105
use FILL  FILL_3167
timestamp 1682952543
transform 1 0 1664 0 1 1170
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1682952543
transform 1 0 1672 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_310
timestamp 1682952543
transform 1 0 1680 0 1 1170
box -8 -3 46 105
use FILL  FILL_3169
timestamp 1682952543
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1682952543
transform 1 0 1728 0 1 1170
box -8 -3 16 105
use FILL  FILL_3171
timestamp 1682952543
transform 1 0 1736 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7188
timestamp 1682952543
transform 1 0 1780 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_311
timestamp 1682952543
transform -1 0 1784 0 1 1170
box -8 -3 46 105
use FILL  FILL_3172
timestamp 1682952543
transform 1 0 1784 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_438
timestamp 1682952543
transform -1 0 1888 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_439
timestamp 1682952543
transform 1 0 1888 0 1 1170
box -8 -3 104 105
use FILL  FILL_3173
timestamp 1682952543
transform 1 0 1984 0 1 1170
box -8 -3 16 105
use FILL  FILL_3174
timestamp 1682952543
transform 1 0 1992 0 1 1170
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1682952543
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7189
timestamp 1682952543
transform 1 0 2020 0 1 1175
box -3 -3 3 3
use FILL  FILL_3176
timestamp 1682952543
transform 1 0 2008 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_495
timestamp 1682952543
transform -1 0 2032 0 1 1170
box -9 -3 26 105
use FILL  FILL_3177
timestamp 1682952543
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1682952543
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3196
timestamp 1682952543
transform 1 0 2048 0 1 1170
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1682952543
transform 1 0 2056 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_313
timestamp 1682952543
transform 1 0 2064 0 1 1170
box -8 -3 46 105
use FILL  FILL_3198
timestamp 1682952543
transform 1 0 2104 0 1 1170
box -8 -3 16 105
use FILL  FILL_3203
timestamp 1682952543
transform 1 0 2112 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_444
timestamp 1682952543
transform 1 0 2120 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_501
timestamp 1682952543
transform 1 0 2216 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_445
timestamp 1682952543
transform 1 0 2232 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_446
timestamp 1682952543
transform 1 0 2328 0 1 1170
box -8 -3 104 105
use FILL  FILL_3204
timestamp 1682952543
transform 1 0 2424 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_314
timestamp 1682952543
transform 1 0 2432 0 1 1170
box -8 -3 46 105
use FILL  FILL_3205
timestamp 1682952543
transform 1 0 2472 0 1 1170
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1682952543
transform 1 0 2480 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_502
timestamp 1682952543
transform -1 0 2504 0 1 1170
box -9 -3 26 105
use FILL  FILL_3207
timestamp 1682952543
transform 1 0 2504 0 1 1170
box -8 -3 16 105
use FILL  FILL_3208
timestamp 1682952543
transform 1 0 2512 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_447
timestamp 1682952543
transform 1 0 2520 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_503
timestamp 1682952543
transform 1 0 2616 0 1 1170
box -9 -3 26 105
use FILL  FILL_3209
timestamp 1682952543
transform 1 0 2632 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_448
timestamp 1682952543
transform 1 0 2640 0 1 1170
box -8 -3 104 105
use FILL  FILL_3210
timestamp 1682952543
transform 1 0 2736 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_507
timestamp 1682952543
transform 1 0 2744 0 1 1170
box -9 -3 26 105
use FILL  FILL_3227
timestamp 1682952543
transform 1 0 2760 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7190
timestamp 1682952543
transform 1 0 2780 0 1 1175
box -3 -3 3 3
use FILL  FILL_3228
timestamp 1682952543
transform 1 0 2768 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_316
timestamp 1682952543
transform 1 0 2776 0 1 1170
box -8 -3 46 105
use FILL  FILL_3229
timestamp 1682952543
transform 1 0 2816 0 1 1170
box -8 -3 16 105
use FILL  FILL_3230
timestamp 1682952543
transform 1 0 2824 0 1 1170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1682952543
transform 1 0 2832 0 1 1170
box -8 -3 16 105
use FILL  FILL_3232
timestamp 1682952543
transform 1 0 2840 0 1 1170
box -8 -3 16 105
use FILL  FILL_3233
timestamp 1682952543
transform 1 0 2848 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_292
timestamp 1682952543
transform 1 0 2856 0 1 1170
box -8 -3 46 105
use FILL  FILL_3234
timestamp 1682952543
transform 1 0 2896 0 1 1170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1682952543
transform 1 0 2904 0 1 1170
box -8 -3 16 105
use FILL  FILL_3236
timestamp 1682952543
transform 1 0 2912 0 1 1170
box -8 -3 16 105
use FILL  FILL_3237
timestamp 1682952543
transform 1 0 2920 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_452
timestamp 1682952543
transform 1 0 2928 0 1 1170
box -8 -3 104 105
use FILL  FILL_3238
timestamp 1682952543
transform 1 0 3024 0 1 1170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1682952543
transform 1 0 3032 0 1 1170
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1682952543
transform 1 0 3040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1682952543
transform 1 0 3048 0 1 1170
box -8 -3 16 105
use FILL  FILL_3256
timestamp 1682952543
transform 1 0 3056 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7191
timestamp 1682952543
transform 1 0 3124 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_7192
timestamp 1682952543
transform 1 0 3156 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_453
timestamp 1682952543
transform -1 0 3160 0 1 1170
box -8 -3 104 105
use FILL  FILL_3257
timestamp 1682952543
transform 1 0 3160 0 1 1170
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1682952543
transform 1 0 3168 0 1 1170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1682952543
transform 1 0 3176 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7193
timestamp 1682952543
transform 1 0 3228 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_317
timestamp 1682952543
transform 1 0 3184 0 1 1170
box -8 -3 46 105
use FILL  FILL_3260
timestamp 1682952543
transform 1 0 3224 0 1 1170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1682952543
transform 1 0 3232 0 1 1170
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1682952543
transform 1 0 3240 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7194
timestamp 1682952543
transform 1 0 3340 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_454
timestamp 1682952543
transform 1 0 3248 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_7195
timestamp 1682952543
transform 1 0 3364 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_510
timestamp 1682952543
transform 1 0 3344 0 1 1170
box -9 -3 26 105
use INVX2  INVX2_511
timestamp 1682952543
transform -1 0 3376 0 1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_318
timestamp 1682952543
transform 1 0 3376 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_7196
timestamp 1682952543
transform 1 0 3428 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_455
timestamp 1682952543
transform 1 0 3416 0 1 1170
box -8 -3 104 105
use FILL  FILL_3263
timestamp 1682952543
transform 1 0 3512 0 1 1170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1682952543
transform 1 0 3520 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_515
timestamp 1682952543
transform 1 0 3528 0 1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_320
timestamp 1682952543
transform 1 0 3544 0 1 1170
box -8 -3 46 105
use FILL  FILL_3282
timestamp 1682952543
transform 1 0 3584 0 1 1170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1682952543
transform 1 0 3592 0 1 1170
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1682952543
transform 1 0 3600 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_516
timestamp 1682952543
transform -1 0 3624 0 1 1170
box -9 -3 26 105
use FILL  FILL_3285
timestamp 1682952543
transform 1 0 3624 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7197
timestamp 1682952543
transform 1 0 3644 0 1 1175
box -3 -3 3 3
use FILL  FILL_3286
timestamp 1682952543
transform 1 0 3632 0 1 1170
box -8 -3 16 105
use FILL  FILL_3287
timestamp 1682952543
transform 1 0 3640 0 1 1170
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1682952543
transform 1 0 3648 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_321
timestamp 1682952543
transform 1 0 3656 0 1 1170
box -8 -3 46 105
use FILL  FILL_3289
timestamp 1682952543
transform 1 0 3696 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_517
timestamp 1682952543
transform -1 0 3720 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_7198
timestamp 1682952543
transform 1 0 3748 0 1 1175
box -3 -3 3 3
use M3_M2  M3_M2_7199
timestamp 1682952543
transform 1 0 3772 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_322
timestamp 1682952543
transform -1 0 3760 0 1 1170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_457
timestamp 1682952543
transform 1 0 3760 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_7200
timestamp 1682952543
transform 1 0 3884 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_518
timestamp 1682952543
transform 1 0 3856 0 1 1170
box -9 -3 26 105
use M3_M2  M3_M2_7201
timestamp 1682952543
transform 1 0 3900 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_458
timestamp 1682952543
transform 1 0 3872 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_519
timestamp 1682952543
transform 1 0 3968 0 1 1170
box -9 -3 26 105
use FILL  FILL_3290
timestamp 1682952543
transform 1 0 3984 0 1 1170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1682952543
transform 1 0 3992 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_323
timestamp 1682952543
transform 1 0 4000 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_7202
timestamp 1682952543
transform 1 0 4052 0 1 1175
box -3 -3 3 3
use FILL  FILL_3301
timestamp 1682952543
transform 1 0 4040 0 1 1170
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1682952543
transform 1 0 4048 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_462
timestamp 1682952543
transform 1 0 4056 0 1 1170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_59
timestamp 1682952543
transform 1 0 4177 0 1 1170
box -10 -3 10 3
use M3_M2  M3_M2_7203
timestamp 1682952543
transform 1 0 132 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7231
timestamp 1682952543
transform 1 0 84 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7252
timestamp 1682952543
transform 1 0 100 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7096
timestamp 1682952543
transform 1 0 84 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7204
timestamp 1682952543
transform 1 0 180 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7253
timestamp 1682952543
transform 1 0 180 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7097
timestamp 1682952543
transform 1 0 180 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7232
timestamp 1682952543
transform 1 0 364 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7254
timestamp 1682952543
transform 1 0 276 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7255
timestamp 1682952543
transform 1 0 388 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7098
timestamp 1682952543
transform 1 0 276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7099
timestamp 1682952543
transform 1 0 364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7100
timestamp 1682952543
transform 1 0 388 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7178
timestamp 1682952543
transform 1 0 116 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7179
timestamp 1682952543
transform 1 0 164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7180
timestamp 1682952543
transform 1 0 212 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7181
timestamp 1682952543
transform 1 0 260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7182
timestamp 1682952543
transform 1 0 324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7183
timestamp 1682952543
transform 1 0 356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7184
timestamp 1682952543
transform 1 0 364 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7321
timestamp 1682952543
transform 1 0 116 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7305
timestamp 1682952543
transform 1 0 388 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7185
timestamp 1682952543
transform 1 0 436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7186
timestamp 1682952543
transform 1 0 468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7187
timestamp 1682952543
transform 1 0 476 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7322
timestamp 1682952543
transform 1 0 324 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7323
timestamp 1682952543
transform 1 0 364 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7324
timestamp 1682952543
transform 1 0 436 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7325
timestamp 1682952543
transform 1 0 476 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7358
timestamp 1682952543
transform 1 0 468 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7383
timestamp 1682952543
transform 1 0 468 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7404
timestamp 1682952543
transform 1 0 476 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7188
timestamp 1682952543
transform 1 0 492 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7326
timestamp 1682952543
transform 1 0 500 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7384
timestamp 1682952543
transform 1 0 492 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7101
timestamp 1682952543
transform 1 0 516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7102
timestamp 1682952543
transform 1 0 524 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7205
timestamp 1682952543
transform 1 0 556 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7233
timestamp 1682952543
transform 1 0 556 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7189
timestamp 1682952543
transform 1 0 532 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7190
timestamp 1682952543
transform 1 0 548 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7359
timestamp 1682952543
transform 1 0 524 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7405
timestamp 1682952543
transform 1 0 540 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7103
timestamp 1682952543
transform 1 0 564 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7104
timestamp 1682952543
transform 1 0 572 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7327
timestamp 1682952543
transform 1 0 564 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7360
timestamp 1682952543
transform 1 0 572 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7234
timestamp 1682952543
transform 1 0 596 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7256
timestamp 1682952543
transform 1 0 596 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7105
timestamp 1682952543
transform 1 0 596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7106
timestamp 1682952543
transform 1 0 612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7191
timestamp 1682952543
transform 1 0 588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7192
timestamp 1682952543
transform 1 0 604 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7385
timestamp 1682952543
transform 1 0 588 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7406
timestamp 1682952543
transform 1 0 580 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7206
timestamp 1682952543
transform 1 0 628 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7193
timestamp 1682952543
transform 1 0 620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7282
timestamp 1682952543
transform 1 0 644 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7235
timestamp 1682952543
transform 1 0 716 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7107
timestamp 1682952543
transform 1 0 652 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7108
timestamp 1682952543
transform 1 0 668 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7194
timestamp 1682952543
transform 1 0 644 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7328
timestamp 1682952543
transform 1 0 620 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7306
timestamp 1682952543
transform 1 0 668 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_7236
timestamp 1682952543
transform 1 0 820 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7109
timestamp 1682952543
transform 1 0 836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7195
timestamp 1682952543
transform 1 0 708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7196
timestamp 1682952543
transform 1 0 748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7197
timestamp 1682952543
transform 1 0 756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7198
timestamp 1682952543
transform 1 0 804 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7407
timestamp 1682952543
transform 1 0 684 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7408
timestamp 1682952543
transform 1 0 708 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7307
timestamp 1682952543
transform 1 0 836 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_7237
timestamp 1682952543
transform 1 0 876 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7238
timestamp 1682952543
transform 1 0 892 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7110
timestamp 1682952543
transform 1 0 860 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7283
timestamp 1682952543
transform 1 0 900 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7308
timestamp 1682952543
transform 1 0 860 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7111
timestamp 1682952543
transform 1 0 1028 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7199
timestamp 1682952543
transform 1 0 900 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7200
timestamp 1682952543
transform 1 0 940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7201
timestamp 1682952543
transform 1 0 948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7202
timestamp 1682952543
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7361
timestamp 1682952543
transform 1 0 852 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7362
timestamp 1682952543
transform 1 0 892 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7093
timestamp 1682952543
transform 1 0 1052 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_7257
timestamp 1682952543
transform 1 0 1060 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7258
timestamp 1682952543
transform 1 0 1084 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7112
timestamp 1682952543
transform 1 0 1076 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7203
timestamp 1682952543
transform 1 0 1084 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7409
timestamp 1682952543
transform 1 0 1076 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7259
timestamp 1682952543
transform 1 0 1188 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7260
timestamp 1682952543
transform 1 0 1204 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7113
timestamp 1682952543
transform 1 0 1100 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7284
timestamp 1682952543
transform 1 0 1180 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7114
timestamp 1682952543
transform 1 0 1188 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7204
timestamp 1682952543
transform 1 0 1124 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7205
timestamp 1682952543
transform 1 0 1180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7115
timestamp 1682952543
transform 1 0 1212 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7309
timestamp 1682952543
transform 1 0 1196 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7206
timestamp 1682952543
transform 1 0 1204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7207
timestamp 1682952543
transform 1 0 1220 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7329
timestamp 1682952543
transform 1 0 1180 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7293
timestamp 1682952543
transform 1 0 1188 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_7410
timestamp 1682952543
transform 1 0 1116 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7411
timestamp 1682952543
transform 1 0 1132 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7330
timestamp 1682952543
transform 1 0 1212 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7207
timestamp 1682952543
transform 1 0 1284 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7208
timestamp 1682952543
transform 1 0 1324 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7239
timestamp 1682952543
transform 1 0 1332 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7285
timestamp 1682952543
transform 1 0 1292 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7116
timestamp 1682952543
transform 1 0 1332 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7208
timestamp 1682952543
transform 1 0 1308 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7331
timestamp 1682952543
transform 1 0 1260 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7332
timestamp 1682952543
transform 1 0 1308 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7240
timestamp 1682952543
transform 1 0 1372 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7241
timestamp 1682952543
transform 1 0 1444 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7117
timestamp 1682952543
transform 1 0 1372 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7209
timestamp 1682952543
transform 1 0 1412 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7210
timestamp 1682952543
transform 1 0 1468 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7211
timestamp 1682952543
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7242
timestamp 1682952543
transform 1 0 1492 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7118
timestamp 1682952543
transform 1 0 1492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7212
timestamp 1682952543
transform 1 0 1500 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7386
timestamp 1682952543
transform 1 0 1500 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7209
timestamp 1682952543
transform 1 0 1532 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7119
timestamp 1682952543
transform 1 0 1516 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7120
timestamp 1682952543
transform 1 0 1532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7213
timestamp 1682952543
transform 1 0 1540 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7286
timestamp 1682952543
transform 1 0 1564 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7287
timestamp 1682952543
transform 1 0 1604 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7121
timestamp 1682952543
transform 1 0 1644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7214
timestamp 1682952543
transform 1 0 1564 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7215
timestamp 1682952543
transform 1 0 1620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7387
timestamp 1682952543
transform 1 0 1564 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7122
timestamp 1682952543
transform 1 0 1668 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7288
timestamp 1682952543
transform 1 0 1716 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7216
timestamp 1682952543
transform 1 0 1716 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7388
timestamp 1682952543
transform 1 0 1684 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7389
timestamp 1682952543
transform 1 0 1748 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7289
timestamp 1682952543
transform 1 0 1764 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7123
timestamp 1682952543
transform 1 0 1772 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7217
timestamp 1682952543
transform 1 0 1764 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7261
timestamp 1682952543
transform 1 0 1796 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7124
timestamp 1682952543
transform 1 0 1788 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7218
timestamp 1682952543
transform 1 0 1780 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7219
timestamp 1682952543
transform 1 0 1796 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7310
timestamp 1682952543
transform 1 0 1804 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_7412
timestamp 1682952543
transform 1 0 1804 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7210
timestamp 1682952543
transform 1 0 1820 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7094
timestamp 1682952543
transform 1 0 1820 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7125
timestamp 1682952543
transform 1 0 1844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7294
timestamp 1682952543
transform 1 0 1836 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_7333
timestamp 1682952543
transform 1 0 1844 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7126
timestamp 1682952543
transform 1 0 1860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7220
timestamp 1682952543
transform 1 0 1860 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7334
timestamp 1682952543
transform 1 0 1860 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7211
timestamp 1682952543
transform 1 0 1900 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7363
timestamp 1682952543
transform 1 0 1908 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7212
timestamp 1682952543
transform 1 0 1932 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7127
timestamp 1682952543
transform 1 0 1924 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7290
timestamp 1682952543
transform 1 0 1972 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7291
timestamp 1682952543
transform 1 0 1996 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7221
timestamp 1682952543
transform 1 0 1972 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7311
timestamp 1682952543
transform 1 0 2004 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_7335
timestamp 1682952543
transform 1 0 1988 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7413
timestamp 1682952543
transform 1 0 2012 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7222
timestamp 1682952543
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7128
timestamp 1682952543
transform 1 0 2052 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7336
timestamp 1682952543
transform 1 0 2044 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7223
timestamp 1682952543
transform 1 0 2060 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7390
timestamp 1682952543
transform 1 0 2052 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7224
timestamp 1682952543
transform 1 0 2076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7129
timestamp 1682952543
transform 1 0 2108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7130
timestamp 1682952543
transform 1 0 2116 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7364
timestamp 1682952543
transform 1 0 2116 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7213
timestamp 1682952543
transform 1 0 2132 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7131
timestamp 1682952543
transform 1 0 2132 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7225
timestamp 1682952543
transform 1 0 2148 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7292
timestamp 1682952543
transform 1 0 2164 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7132
timestamp 1682952543
transform 1 0 2172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7226
timestamp 1682952543
transform 1 0 2164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7227
timestamp 1682952543
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7337
timestamp 1682952543
transform 1 0 2164 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7365
timestamp 1682952543
transform 1 0 2156 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7095
timestamp 1682952543
transform 1 0 2196 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7133
timestamp 1682952543
transform 1 0 2196 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7338
timestamp 1682952543
transform 1 0 2196 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7366
timestamp 1682952543
transform 1 0 2188 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7391
timestamp 1682952543
transform 1 0 2172 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7414
timestamp 1682952543
transform 1 0 2180 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7214
timestamp 1682952543
transform 1 0 2244 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7293
timestamp 1682952543
transform 1 0 2236 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7134
timestamp 1682952543
transform 1 0 2244 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7262
timestamp 1682952543
transform 1 0 2276 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7135
timestamp 1682952543
transform 1 0 2276 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7136
timestamp 1682952543
transform 1 0 2292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7137
timestamp 1682952543
transform 1 0 2300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7228
timestamp 1682952543
transform 1 0 2260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7229
timestamp 1682952543
transform 1 0 2268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7230
timestamp 1682952543
transform 1 0 2284 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7339
timestamp 1682952543
transform 1 0 2292 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7392
timestamp 1682952543
transform 1 0 2268 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7215
timestamp 1682952543
transform 1 0 2340 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7138
timestamp 1682952543
transform 1 0 2412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7231
timestamp 1682952543
transform 1 0 2316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7232
timestamp 1682952543
transform 1 0 2324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7233
timestamp 1682952543
transform 1 0 2332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7234
timestamp 1682952543
transform 1 0 2364 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7340
timestamp 1682952543
transform 1 0 2324 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7341
timestamp 1682952543
transform 1 0 2364 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7367
timestamp 1682952543
transform 1 0 2332 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7393
timestamp 1682952543
transform 1 0 2316 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7394
timestamp 1682952543
transform 1 0 2412 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7216
timestamp 1682952543
transform 1 0 2436 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7139
timestamp 1682952543
transform 1 0 2436 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7140
timestamp 1682952543
transform 1 0 2524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7235
timestamp 1682952543
transform 1 0 2460 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7236
timestamp 1682952543
transform 1 0 2516 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7342
timestamp 1682952543
transform 1 0 2436 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7343
timestamp 1682952543
transform 1 0 2484 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7344
timestamp 1682952543
transform 1 0 2516 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7415
timestamp 1682952543
transform 1 0 2436 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7416
timestamp 1682952543
transform 1 0 2468 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7417
timestamp 1682952543
transform 1 0 2508 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7263
timestamp 1682952543
transform 1 0 2596 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7141
timestamp 1682952543
transform 1 0 2628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7142
timestamp 1682952543
transform 1 0 2644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7237
timestamp 1682952543
transform 1 0 2540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7238
timestamp 1682952543
transform 1 0 2548 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7239
timestamp 1682952543
transform 1 0 2580 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7345
timestamp 1682952543
transform 1 0 2540 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7312
timestamp 1682952543
transform 1 0 2628 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_7346
timestamp 1682952543
transform 1 0 2580 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7264
timestamp 1682952543
transform 1 0 2668 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7240
timestamp 1682952543
transform 1 0 2652 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7313
timestamp 1682952543
transform 1 0 2660 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7143
timestamp 1682952543
transform 1 0 2676 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7241
timestamp 1682952543
transform 1 0 2668 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7368
timestamp 1682952543
transform 1 0 2636 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7418
timestamp 1682952543
transform 1 0 2556 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7369
timestamp 1682952543
transform 1 0 2668 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7314
timestamp 1682952543
transform 1 0 2708 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7242
timestamp 1682952543
transform 1 0 2716 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7370
timestamp 1682952543
transform 1 0 2724 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7395
timestamp 1682952543
transform 1 0 2724 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7295
timestamp 1682952543
transform 1 0 2740 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7243
timestamp 1682952543
transform 1 0 2764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7244
timestamp 1682952543
transform 1 0 2788 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7347
timestamp 1682952543
transform 1 0 2788 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7303
timestamp 1682952543
transform 1 0 2788 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_7396
timestamp 1682952543
transform 1 0 2780 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7265
timestamp 1682952543
transform 1 0 2820 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7144
timestamp 1682952543
transform 1 0 2820 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7266
timestamp 1682952543
transform 1 0 2852 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7145
timestamp 1682952543
transform 1 0 2852 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7294
timestamp 1682952543
transform 1 0 2860 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7245
timestamp 1682952543
transform 1 0 2820 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7246
timestamp 1682952543
transform 1 0 2836 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7247
timestamp 1682952543
transform 1 0 2852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7248
timestamp 1682952543
transform 1 0 2860 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7249
timestamp 1682952543
transform 1 0 2868 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7296
timestamp 1682952543
transform 1 0 2812 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_7371
timestamp 1682952543
transform 1 0 2812 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7397
timestamp 1682952543
transform 1 0 2812 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7372
timestamp 1682952543
transform 1 0 2836 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7373
timestamp 1682952543
transform 1 0 2852 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7398
timestamp 1682952543
transform 1 0 2836 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7399
timestamp 1682952543
transform 1 0 2860 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7374
timestamp 1682952543
transform 1 0 2876 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7250
timestamp 1682952543
transform 1 0 2916 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7297
timestamp 1682952543
transform 1 0 2900 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7304
timestamp 1682952543
transform 1 0 2908 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_7400
timestamp 1682952543
transform 1 0 2916 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7251
timestamp 1682952543
transform 1 0 2932 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7315
timestamp 1682952543
transform 1 0 2948 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7298
timestamp 1682952543
transform 1 0 2948 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_7419
timestamp 1682952543
transform 1 0 2940 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7217
timestamp 1682952543
transform 1 0 2980 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7146
timestamp 1682952543
transform 1 0 2964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7147
timestamp 1682952543
transform 1 0 2980 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7252
timestamp 1682952543
transform 1 0 2972 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7348
timestamp 1682952543
transform 1 0 2972 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7218
timestamp 1682952543
transform 1 0 2996 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7253
timestamp 1682952543
transform 1 0 2996 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7254
timestamp 1682952543
transform 1 0 3004 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7420
timestamp 1682952543
transform 1 0 2996 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7267
timestamp 1682952543
transform 1 0 3028 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7148
timestamp 1682952543
transform 1 0 3020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7255
timestamp 1682952543
transform 1 0 3028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7149
timestamp 1682952543
transform 1 0 3052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7150
timestamp 1682952543
transform 1 0 3068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7256
timestamp 1682952543
transform 1 0 3076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7151
timestamp 1682952543
transform 1 0 3116 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7257
timestamp 1682952543
transform 1 0 3132 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7219
timestamp 1682952543
transform 1 0 3172 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7152
timestamp 1682952543
transform 1 0 3156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7153
timestamp 1682952543
transform 1 0 3172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7258
timestamp 1682952543
transform 1 0 3148 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7259
timestamp 1682952543
transform 1 0 3164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7260
timestamp 1682952543
transform 1 0 3172 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7220
timestamp 1682952543
transform 1 0 3196 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7268
timestamp 1682952543
transform 1 0 3188 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7299
timestamp 1682952543
transform 1 0 3180 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_7295
timestamp 1682952543
transform 1 0 3196 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7261
timestamp 1682952543
transform 1 0 3204 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7262
timestamp 1682952543
transform 1 0 3220 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7349
timestamp 1682952543
transform 1 0 3204 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7300
timestamp 1682952543
transform 1 0 3212 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7305
timestamp 1682952543
transform 1 0 3196 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_7375
timestamp 1682952543
transform 1 0 3212 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7243
timestamp 1682952543
transform 1 0 3260 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7269
timestamp 1682952543
transform 1 0 3244 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7154
timestamp 1682952543
transform 1 0 3244 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7296
timestamp 1682952543
transform 1 0 3260 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7263
timestamp 1682952543
transform 1 0 3228 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7264
timestamp 1682952543
transform 1 0 3236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7265
timestamp 1682952543
transform 1 0 3252 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7350
timestamp 1682952543
transform 1 0 3252 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7421
timestamp 1682952543
transform 1 0 3244 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_7270
timestamp 1682952543
transform 1 0 3300 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7155
timestamp 1682952543
transform 1 0 3292 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7156
timestamp 1682952543
transform 1 0 3300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7266
timestamp 1682952543
transform 1 0 3284 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7401
timestamp 1682952543
transform 1 0 3276 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7297
timestamp 1682952543
transform 1 0 3316 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7271
timestamp 1682952543
transform 1 0 3332 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7157
timestamp 1682952543
transform 1 0 3324 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7267
timestamp 1682952543
transform 1 0 3316 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7298
timestamp 1682952543
transform 1 0 3348 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7158
timestamp 1682952543
transform 1 0 3356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7159
timestamp 1682952543
transform 1 0 3364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7268
timestamp 1682952543
transform 1 0 3332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7269
timestamp 1682952543
transform 1 0 3348 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7270
timestamp 1682952543
transform 1 0 3364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7271
timestamp 1682952543
transform 1 0 3372 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7351
timestamp 1682952543
transform 1 0 3340 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7376
timestamp 1682952543
transform 1 0 3348 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7377
timestamp 1682952543
transform 1 0 3364 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7272
timestamp 1682952543
transform 1 0 3436 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7160
timestamp 1682952543
transform 1 0 3460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7272
timestamp 1682952543
transform 1 0 3412 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7352
timestamp 1682952543
transform 1 0 3412 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7402
timestamp 1682952543
transform 1 0 3460 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7273
timestamp 1682952543
transform 1 0 3476 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7221
timestamp 1682952543
transform 1 0 3500 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7244
timestamp 1682952543
transform 1 0 3516 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7161
timestamp 1682952543
transform 1 0 3476 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7299
timestamp 1682952543
transform 1 0 3484 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7300
timestamp 1682952543
transform 1 0 3500 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7273
timestamp 1682952543
transform 1 0 3484 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7316
timestamp 1682952543
transform 1 0 3492 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7274
timestamp 1682952543
transform 1 0 3500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7275
timestamp 1682952543
transform 1 0 3516 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7301
timestamp 1682952543
transform 1 0 3524 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_7378
timestamp 1682952543
transform 1 0 3516 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7222
timestamp 1682952543
transform 1 0 3548 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7223
timestamp 1682952543
transform 1 0 3564 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7224
timestamp 1682952543
transform 1 0 3588 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7225
timestamp 1682952543
transform 1 0 3604 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7162
timestamp 1682952543
transform 1 0 3540 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7317
timestamp 1682952543
transform 1 0 3540 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7302
timestamp 1682952543
transform 1 0 3540 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_7245
timestamp 1682952543
transform 1 0 3580 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7274
timestamp 1682952543
transform 1 0 3556 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7163
timestamp 1682952543
transform 1 0 3556 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7276
timestamp 1682952543
transform 1 0 3588 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7318
timestamp 1682952543
transform 1 0 3596 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_7226
timestamp 1682952543
transform 1 0 3708 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7246
timestamp 1682952543
transform 1 0 3668 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7247
timestamp 1682952543
transform 1 0 3692 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7164
timestamp 1682952543
transform 1 0 3652 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7227
timestamp 1682952543
transform 1 0 3756 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7228
timestamp 1682952543
transform 1 0 3788 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7248
timestamp 1682952543
transform 1 0 3836 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7275
timestamp 1682952543
transform 1 0 3772 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7276
timestamp 1682952543
transform 1 0 3796 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7277
timestamp 1682952543
transform 1 0 3852 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7278
timestamp 1682952543
transform 1 0 3868 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7165
timestamp 1682952543
transform 1 0 3748 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7166
timestamp 1682952543
transform 1 0 3836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7167
timestamp 1682952543
transform 1 0 3852 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7301
timestamp 1682952543
transform 1 0 3860 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7168
timestamp 1682952543
transform 1 0 3868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7169
timestamp 1682952543
transform 1 0 3876 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7277
timestamp 1682952543
transform 1 0 3636 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7278
timestamp 1682952543
transform 1 0 3676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7279
timestamp 1682952543
transform 1 0 3732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7280
timestamp 1682952543
transform 1 0 3796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7281
timestamp 1682952543
transform 1 0 3836 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7282
timestamp 1682952543
transform 1 0 3844 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7283
timestamp 1682952543
transform 1 0 3860 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7353
timestamp 1682952543
transform 1 0 3556 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7403
timestamp 1682952543
transform 1 0 3636 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_7354
timestamp 1682952543
transform 1 0 3836 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7302
timestamp 1682952543
transform 1 0 3884 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7284
timestamp 1682952543
transform 1 0 3884 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7355
timestamp 1682952543
transform 1 0 3876 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7379
timestamp 1682952543
transform 1 0 3876 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7279
timestamp 1682952543
transform 1 0 3916 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_7380
timestamp 1682952543
transform 1 0 3908 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7170
timestamp 1682952543
transform 1 0 3916 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7249
timestamp 1682952543
transform 1 0 3940 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7229
timestamp 1682952543
transform 1 0 4012 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7250
timestamp 1682952543
transform 1 0 4004 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7171
timestamp 1682952543
transform 1 0 3964 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7303
timestamp 1682952543
transform 1 0 3972 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7280
timestamp 1682952543
transform 1 0 4020 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7172
timestamp 1682952543
transform 1 0 3980 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7173
timestamp 1682952543
transform 1 0 3996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7174
timestamp 1682952543
transform 1 0 4004 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_7304
timestamp 1682952543
transform 1 0 4012 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_7230
timestamp 1682952543
transform 1 0 4108 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_7251
timestamp 1682952543
transform 1 0 4092 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_7281
timestamp 1682952543
transform 1 0 4076 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7175
timestamp 1682952543
transform 1 0 4020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7176
timestamp 1682952543
transform 1 0 4036 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7177
timestamp 1682952543
transform 1 0 4052 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7285
timestamp 1682952543
transform 1 0 3956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7286
timestamp 1682952543
transform 1 0 3972 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7287
timestamp 1682952543
transform 1 0 3980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7288
timestamp 1682952543
transform 1 0 3988 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7381
timestamp 1682952543
transform 1 0 3948 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_7319
timestamp 1682952543
transform 1 0 3996 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7289
timestamp 1682952543
transform 1 0 4012 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7290
timestamp 1682952543
transform 1 0 4028 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7356
timestamp 1682952543
transform 1 0 3988 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7357
timestamp 1682952543
transform 1 0 4028 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_7382
timestamp 1682952543
transform 1 0 4028 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7291
timestamp 1682952543
transform 1 0 4076 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_7320
timestamp 1682952543
transform 1 0 4124 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7292
timestamp 1682952543
transform 1 0 4132 0 1 1125
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_60
timestamp 1682952543
transform 1 0 24 0 1 1070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_425
timestamp 1682952543
transform 1 0 72 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_426
timestamp 1682952543
transform 1 0 168 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_427
timestamp 1682952543
transform 1 0 264 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_485
timestamp 1682952543
transform 1 0 360 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_428
timestamp 1682952543
transform 1 0 376 0 -1 1170
box -8 -3 104 105
use FILL  FILL_3094
timestamp 1682952543
transform 1 0 472 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_486
timestamp 1682952543
transform -1 0 496 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3095
timestamp 1682952543
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1682952543
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_290
timestamp 1682952543
transform -1 0 552 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3097
timestamp 1682952543
transform 1 0 552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1682952543
transform 1 0 560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1682952543
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7422
timestamp 1682952543
transform 1 0 604 0 1 1075
box -3 -3 3 3
use OAI22X1  OAI22X1_306
timestamp 1682952543
transform 1 0 576 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3124
timestamp 1682952543
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use AND2X2  AND2X2_51
timestamp 1682952543
transform -1 0 656 0 -1 1170
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_431
timestamp 1682952543
transform 1 0 656 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_432
timestamp 1682952543
transform -1 0 848 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_433
timestamp 1682952543
transform 1 0 848 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_434
timestamp 1682952543
transform -1 0 1040 0 -1 1170
box -8 -3 104 105
use FILL  FILL_3125
timestamp 1682952543
transform 1 0 1040 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_87
timestamp 1682952543
transform 1 0 1048 0 -1 1170
box -8 -3 32 105
use FILL  FILL_3136
timestamp 1682952543
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1682952543
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_435
timestamp 1682952543
transform 1 0 1088 0 -1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_124
timestamp 1682952543
transform -1 0 1216 0 -1 1170
box -8 -3 34 105
use INVX2  INVX2_491
timestamp 1682952543
transform -1 0 1232 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3138
timestamp 1682952543
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1682952543
transform 1 0 1240 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_436
timestamp 1682952543
transform -1 0 1344 0 -1 1170
box -8 -3 104 105
use FILL  FILL_3149
timestamp 1682952543
transform 1 0 1344 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3151
timestamp 1682952543
transform 1 0 1352 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_440
timestamp 1682952543
transform 1 0 1360 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_496
timestamp 1682952543
transform 1 0 1456 0 -1 1170
box -9 -3 26 105
use BUFX2  BUFX2_97
timestamp 1682952543
transform 1 0 1472 0 -1 1170
box -5 -3 28 105
use FILL  FILL_3178
timestamp 1682952543
transform 1 0 1496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1682952543
transform 1 0 1504 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7423
timestamp 1682952543
transform 1 0 1540 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_7424
timestamp 1682952543
transform 1 0 1556 0 1 1075
box -3 -3 3 3
use OAI22X1  OAI22X1_312
timestamp 1682952543
transform 1 0 1512 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3180
timestamp 1682952543
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_441
timestamp 1682952543
transform -1 0 1656 0 -1 1170
box -8 -3 104 105
use M3_M2  M3_M2_7425
timestamp 1682952543
transform 1 0 1708 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_7426
timestamp 1682952543
transform 1 0 1756 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_442
timestamp 1682952543
transform 1 0 1656 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_497
timestamp 1682952543
transform 1 0 1752 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_498
timestamp 1682952543
transform 1 0 1768 0 -1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_125
timestamp 1682952543
transform 1 0 1784 0 -1 1170
box -8 -3 34 105
use FILL  FILL_3181
timestamp 1682952543
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1682952543
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3183
timestamp 1682952543
transform 1 0 1832 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_88
timestamp 1682952543
transform 1 0 1840 0 -1 1170
box -8 -3 32 105
use FILL  FILL_3184
timestamp 1682952543
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1682952543
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3186
timestamp 1682952543
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1682952543
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1682952543
transform 1 0 1896 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1682952543
transform 1 0 1904 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_443
timestamp 1682952543
transform 1 0 1912 0 -1 1170
box -8 -3 104 105
use FILL  FILL_3190
timestamp 1682952543
transform 1 0 2008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1682952543
transform 1 0 2016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1682952543
transform 1 0 2024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1682952543
transform 1 0 2032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1682952543
transform 1 0 2040 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_499
timestamp 1682952543
transform 1 0 2048 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3199
timestamp 1682952543
transform 1 0 2064 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_500
timestamp 1682952543
transform -1 0 2088 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3200
timestamp 1682952543
transform 1 0 2088 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1682952543
transform 1 0 2096 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1682952543
transform 1 0 2104 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_504
timestamp 1682952543
transform 1 0 2112 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3211
timestamp 1682952543
transform 1 0 2128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1682952543
transform 1 0 2136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3213
timestamp 1682952543
transform 1 0 2144 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_315
timestamp 1682952543
transform -1 0 2192 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3214
timestamp 1682952543
transform 1 0 2192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1682952543
transform 1 0 2200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1682952543
transform 1 0 2208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3217
timestamp 1682952543
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_89
timestamp 1682952543
transform 1 0 2224 0 -1 1170
box -8 -3 32 105
use FILL  FILL_3218
timestamp 1682952543
transform 1 0 2248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1682952543
transform 1 0 2256 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7427
timestamp 1682952543
transform 1 0 2308 0 1 1075
box -3 -3 3 3
use AOI22X1  AOI22X1_291
timestamp 1682952543
transform 1 0 2264 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3220
timestamp 1682952543
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_505
timestamp 1682952543
transform 1 0 2312 0 -1 1170
box -9 -3 26 105
use M3_M2  M3_M2_7428
timestamp 1682952543
transform 1 0 2388 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_7429
timestamp 1682952543
transform 1 0 2404 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_449
timestamp 1682952543
transform -1 0 2424 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_450
timestamp 1682952543
transform 1 0 2424 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_506
timestamp 1682952543
transform 1 0 2520 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3221
timestamp 1682952543
transform 1 0 2536 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_451
timestamp 1682952543
transform -1 0 2640 0 -1 1170
box -8 -3 104 105
use M3_M2  M3_M2_7430
timestamp 1682952543
transform 1 0 2676 0 1 1075
box -3 -3 3 3
use AND2X2  AND2X2_52
timestamp 1682952543
transform 1 0 2640 0 -1 1170
box -8 -3 40 105
use FILL  FILL_3222
timestamp 1682952543
transform 1 0 2672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1682952543
transform 1 0 2680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1682952543
transform 1 0 2688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1682952543
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7431
timestamp 1682952543
transform 1 0 2732 0 1 1075
box -3 -3 3 3
use AND2X2  AND2X2_53
timestamp 1682952543
transform 1 0 2704 0 -1 1170
box -8 -3 40 105
use FILL  FILL_3226
timestamp 1682952543
transform 1 0 2736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1682952543
transform 1 0 2744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1682952543
transform 1 0 2752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1682952543
transform 1 0 2760 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_62
timestamp 1682952543
transform -1 0 2800 0 -1 1170
box -8 -3 40 105
use M3_M2  M3_M2_7432
timestamp 1682952543
transform 1 0 2812 0 1 1075
box -3 -3 3 3
use FILL  FILL_3242
timestamp 1682952543
transform 1 0 2800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1682952543
transform 1 0 2808 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_293
timestamp 1682952543
transform -1 0 2856 0 -1 1170
box -8 -3 46 105
use INVX2  INVX2_508
timestamp 1682952543
transform -1 0 2872 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3244
timestamp 1682952543
transform 1 0 2872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3245
timestamp 1682952543
transform 1 0 2880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1682952543
transform 1 0 2888 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_63
timestamp 1682952543
transform -1 0 2928 0 -1 1170
box -8 -3 40 105
use FILL  FILL_3247
timestamp 1682952543
transform 1 0 2928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1682952543
transform 1 0 2936 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3249
timestamp 1682952543
transform 1 0 2944 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7433
timestamp 1682952543
transform 1 0 2996 0 1 1075
box -3 -3 3 3
use AOI22X1  AOI22X1_294
timestamp 1682952543
transform 1 0 2952 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3250
timestamp 1682952543
transform 1 0 2992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1682952543
transform 1 0 3000 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_509
timestamp 1682952543
transform -1 0 3024 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3252
timestamp 1682952543
transform 1 0 3024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3265
timestamp 1682952543
transform 1 0 3032 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_512
timestamp 1682952543
transform -1 0 3056 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3266
timestamp 1682952543
transform 1 0 3056 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1682952543
transform 1 0 3064 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1682952543
transform 1 0 3072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3269
timestamp 1682952543
transform 1 0 3080 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_513
timestamp 1682952543
transform 1 0 3088 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3270
timestamp 1682952543
transform 1 0 3104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1682952543
transform 1 0 3112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3272
timestamp 1682952543
transform 1 0 3120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1682952543
transform 1 0 3128 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_319
timestamp 1682952543
transform -1 0 3176 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3274
timestamp 1682952543
transform 1 0 3176 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_64
timestamp 1682952543
transform -1 0 3216 0 -1 1170
box -8 -3 40 105
use INVX2  INVX2_514
timestamp 1682952543
transform 1 0 3216 0 -1 1170
box -9 -3 26 105
use AOI22X1  AOI22X1_295
timestamp 1682952543
transform -1 0 3272 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3275
timestamp 1682952543
transform 1 0 3272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1682952543
transform 1 0 3280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1682952543
transform 1 0 3288 0 -1 1170
box -8 -3 16 105
use BUFX2  BUFX2_98
timestamp 1682952543
transform -1 0 3320 0 -1 1170
box -5 -3 28 105
use FILL  FILL_3278
timestamp 1682952543
transform 1 0 3320 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_296
timestamp 1682952543
transform 1 0 3328 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3279
timestamp 1682952543
transform 1 0 3368 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_456
timestamp 1682952543
transform -1 0 3472 0 -1 1170
box -8 -3 104 105
use FILL  FILL_3280
timestamp 1682952543
transform 1 0 3472 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_297
timestamp 1682952543
transform 1 0 3480 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3281
timestamp 1682952543
transform 1 0 3520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3292
timestamp 1682952543
transform 1 0 3528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1682952543
transform 1 0 3536 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_459
timestamp 1682952543
transform 1 0 3544 0 -1 1170
box -8 -3 104 105
use M3_M2  M3_M2_7434
timestamp 1682952543
transform 1 0 3668 0 1 1075
box -3 -3 3 3
use M3_M2  M3_M2_7435
timestamp 1682952543
transform 1 0 3692 0 1 1075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_460
timestamp 1682952543
transform 1 0 3640 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_461
timestamp 1682952543
transform 1 0 3736 0 -1 1170
box -8 -3 104 105
use OAI22X1  OAI22X1_324
timestamp 1682952543
transform 1 0 3832 0 -1 1170
box -8 -3 46 105
use FILL  FILL_3294
timestamp 1682952543
transform 1 0 3872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1682952543
transform 1 0 3880 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_520
timestamp 1682952543
transform 1 0 3888 0 -1 1170
box -9 -3 26 105
use FILL  FILL_3296
timestamp 1682952543
transform 1 0 3904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3297
timestamp 1682952543
transform 1 0 3912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1682952543
transform 1 0 3920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1682952543
transform 1 0 3928 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1682952543
transform 1 0 3936 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_7436
timestamp 1682952543
transform 1 0 3956 0 1 1075
box -3 -3 3 3
use OAI22X1  OAI22X1_325
timestamp 1682952543
transform -1 0 3984 0 -1 1170
box -8 -3 46 105
use M3_M2  M3_M2_7437
timestamp 1682952543
transform 1 0 3996 0 1 1075
box -3 -3 3 3
use INVX2  INVX2_521
timestamp 1682952543
transform -1 0 4000 0 -1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_326
timestamp 1682952543
transform 1 0 4000 0 -1 1170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_463
timestamp 1682952543
transform 1 0 4040 0 -1 1170
box -8 -3 104 105
use FILL  FILL_3303
timestamp 1682952543
transform 1 0 4136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1682952543
transform 1 0 4144 0 -1 1170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_61
timestamp 1682952543
transform 1 0 4201 0 1 1070
box -10 -3 10 3
use M3_M2  M3_M2_7500
timestamp 1682952543
transform 1 0 124 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7501
timestamp 1682952543
transform 1 0 172 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7502
timestamp 1682952543
transform 1 0 188 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7312
timestamp 1682952543
transform 1 0 124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7313
timestamp 1682952543
transform 1 0 164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7314
timestamp 1682952543
transform 1 0 172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7315
timestamp 1682952543
transform 1 0 188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7316
timestamp 1682952543
transform 1 0 204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7449
timestamp 1682952543
transform 1 0 84 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7568
timestamp 1682952543
transform 1 0 172 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7450
timestamp 1682952543
transform 1 0 180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7451
timestamp 1682952543
transform 1 0 196 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7604
timestamp 1682952543
transform 1 0 164 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7569
timestamp 1682952543
transform 1 0 204 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7438
timestamp 1682952543
transform 1 0 324 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7461
timestamp 1682952543
transform 1 0 332 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7503
timestamp 1682952543
transform 1 0 324 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7534
timestamp 1682952543
transform 1 0 236 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7317
timestamp 1682952543
transform 1 0 260 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7535
timestamp 1682952543
transform 1 0 276 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7318
timestamp 1682952543
transform 1 0 316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7319
timestamp 1682952543
transform 1 0 324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7320
timestamp 1682952543
transform 1 0 340 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7321
timestamp 1682952543
transform 1 0 356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7322
timestamp 1682952543
transform 1 0 364 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7323
timestamp 1682952543
transform 1 0 372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7324
timestamp 1682952543
transform 1 0 388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7452
timestamp 1682952543
transform 1 0 212 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7453
timestamp 1682952543
transform 1 0 220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7454
timestamp 1682952543
transform 1 0 236 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7455
timestamp 1682952543
transform 1 0 324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7456
timestamp 1682952543
transform 1 0 348 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7605
timestamp 1682952543
transform 1 0 212 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7536
timestamp 1682952543
transform 1 0 404 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7462
timestamp 1682952543
transform 1 0 452 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7504
timestamp 1682952543
transform 1 0 484 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7505
timestamp 1682952543
transform 1 0 524 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7475
timestamp 1682952543
transform 1 0 548 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7325
timestamp 1682952543
transform 1 0 420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7326
timestamp 1682952543
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7327
timestamp 1682952543
transform 1 0 516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7328
timestamp 1682952543
transform 1 0 524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7329
timestamp 1682952543
transform 1 0 532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7457
timestamp 1682952543
transform 1 0 380 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7570
timestamp 1682952543
transform 1 0 388 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7458
timestamp 1682952543
transform 1 0 396 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7459
timestamp 1682952543
transform 1 0 404 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7606
timestamp 1682952543
transform 1 0 396 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7460
timestamp 1682952543
transform 1 0 436 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7537
timestamp 1682952543
transform 1 0 548 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7330
timestamp 1682952543
transform 1 0 556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7331
timestamp 1682952543
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7538
timestamp 1682952543
transform 1 0 604 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7446
timestamp 1682952543
transform 1 0 652 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7463
timestamp 1682952543
transform 1 0 636 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7476
timestamp 1682952543
transform 1 0 644 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7332
timestamp 1682952543
transform 1 0 620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7333
timestamp 1682952543
transform 1 0 636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7334
timestamp 1682952543
transform 1 0 652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7461
timestamp 1682952543
transform 1 0 540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7462
timestamp 1682952543
transform 1 0 548 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7463
timestamp 1682952543
transform 1 0 564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7464
timestamp 1682952543
transform 1 0 580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7465
timestamp 1682952543
transform 1 0 588 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7466
timestamp 1682952543
transform 1 0 604 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7467
timestamp 1682952543
transform 1 0 612 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7607
timestamp 1682952543
transform 1 0 452 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7608
timestamp 1682952543
transform 1 0 476 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7609
timestamp 1682952543
transform 1 0 516 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7610
timestamp 1682952543
transform 1 0 564 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7611
timestamp 1682952543
transform 1 0 612 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7571
timestamp 1682952543
transform 1 0 652 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7612
timestamp 1682952543
transform 1 0 644 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7557
timestamp 1682952543
transform 1 0 652 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7468
timestamp 1682952543
transform 1 0 668 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7477
timestamp 1682952543
transform 1 0 708 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7307
timestamp 1682952543
transform 1 0 692 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_7539
timestamp 1682952543
transform 1 0 692 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7439
timestamp 1682952543
transform 1 0 732 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7447
timestamp 1682952543
transform 1 0 740 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7506
timestamp 1682952543
transform 1 0 732 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7335
timestamp 1682952543
transform 1 0 724 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7572
timestamp 1682952543
transform 1 0 724 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7507
timestamp 1682952543
transform 1 0 756 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7508
timestamp 1682952543
transform 1 0 772 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7336
timestamp 1682952543
transform 1 0 740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7337
timestamp 1682952543
transform 1 0 756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7469
timestamp 1682952543
transform 1 0 732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7470
timestamp 1682952543
transform 1 0 748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7471
timestamp 1682952543
transform 1 0 772 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7613
timestamp 1682952543
transform 1 0 756 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7614
timestamp 1682952543
transform 1 0 772 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7558
timestamp 1682952543
transform 1 0 780 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_7639
timestamp 1682952543
transform 1 0 748 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7640
timestamp 1682952543
transform 1 0 764 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7478
timestamp 1682952543
transform 1 0 788 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7338
timestamp 1682952543
transform 1 0 788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7339
timestamp 1682952543
transform 1 0 804 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7573
timestamp 1682952543
transform 1 0 804 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7472
timestamp 1682952543
transform 1 0 820 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7641
timestamp 1682952543
transform 1 0 820 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7340
timestamp 1682952543
transform 1 0 844 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7479
timestamp 1682952543
transform 1 0 892 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7509
timestamp 1682952543
transform 1 0 876 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7341
timestamp 1682952543
transform 1 0 860 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7342
timestamp 1682952543
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7343
timestamp 1682952543
transform 1 0 892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7344
timestamp 1682952543
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7473
timestamp 1682952543
transform 1 0 868 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7615
timestamp 1682952543
transform 1 0 876 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7510
timestamp 1682952543
transform 1 0 908 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7574
timestamp 1682952543
transform 1 0 900 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7474
timestamp 1682952543
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7559
timestamp 1682952543
transform 1 0 908 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_7642
timestamp 1682952543
transform 1 0 908 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7475
timestamp 1682952543
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7616
timestamp 1682952543
transform 1 0 932 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7643
timestamp 1682952543
transform 1 0 940 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7511
timestamp 1682952543
transform 1 0 964 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7575
timestamp 1682952543
transform 1 0 956 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7512
timestamp 1682952543
transform 1 0 980 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7540
timestamp 1682952543
transform 1 0 980 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7476
timestamp 1682952543
transform 1 0 980 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7345
timestamp 1682952543
transform 1 0 996 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7480
timestamp 1682952543
transform 1 0 1036 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7308
timestamp 1682952543
transform 1 0 1012 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_7481
timestamp 1682952543
transform 1 0 1076 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7513
timestamp 1682952543
transform 1 0 1060 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7346
timestamp 1682952543
transform 1 0 1028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7347
timestamp 1682952543
transform 1 0 1036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7348
timestamp 1682952543
transform 1 0 1060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7349
timestamp 1682952543
transform 1 0 1076 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7477
timestamp 1682952543
transform 1 0 1036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7478
timestamp 1682952543
transform 1 0 1052 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7576
timestamp 1682952543
transform 1 0 1060 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7479
timestamp 1682952543
transform 1 0 1068 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7514
timestamp 1682952543
transform 1 0 1108 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7480
timestamp 1682952543
transform 1 0 1108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7309
timestamp 1682952543
transform 1 0 1132 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7350
timestamp 1682952543
transform 1 0 1124 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7577
timestamp 1682952543
transform 1 0 1172 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7440
timestamp 1682952543
transform 1 0 1204 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7515
timestamp 1682952543
transform 1 0 1204 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7351
timestamp 1682952543
transform 1 0 1196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7352
timestamp 1682952543
transform 1 0 1204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7481
timestamp 1682952543
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7482
timestamp 1682952543
transform 1 0 1220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7306
timestamp 1682952543
transform 1 0 1244 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_7353
timestamp 1682952543
transform 1 0 1236 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7617
timestamp 1682952543
transform 1 0 1236 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7448
timestamp 1682952543
transform 1 0 1268 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7483
timestamp 1682952543
transform 1 0 1260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7484
timestamp 1682952543
transform 1 0 1268 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7354
timestamp 1682952543
transform 1 0 1276 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7441
timestamp 1682952543
transform 1 0 1316 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_7355
timestamp 1682952543
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7644
timestamp 1682952543
transform 1 0 1340 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7449
timestamp 1682952543
transform 1 0 1356 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7356
timestamp 1682952543
transform 1 0 1356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7357
timestamp 1682952543
transform 1 0 1396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7358
timestamp 1682952543
transform 1 0 1452 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7485
timestamp 1682952543
transform 1 0 1372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7486
timestamp 1682952543
transform 1 0 1460 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7645
timestamp 1682952543
transform 1 0 1372 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7646
timestamp 1682952543
transform 1 0 1460 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7359
timestamp 1682952543
transform 1 0 1476 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7541
timestamp 1682952543
transform 1 0 1508 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7360
timestamp 1682952543
transform 1 0 1516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7487
timestamp 1682952543
transform 1 0 1500 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7578
timestamp 1682952543
transform 1 0 1508 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7542
timestamp 1682952543
transform 1 0 1532 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7488
timestamp 1682952543
transform 1 0 1524 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7560
timestamp 1682952543
transform 1 0 1524 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_7482
timestamp 1682952543
transform 1 0 1556 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7483
timestamp 1682952543
transform 1 0 1580 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7361
timestamp 1682952543
transform 1 0 1548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7362
timestamp 1682952543
transform 1 0 1564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7363
timestamp 1682952543
transform 1 0 1580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7561
timestamp 1682952543
transform 1 0 1540 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7489
timestamp 1682952543
transform 1 0 1556 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7579
timestamp 1682952543
transform 1 0 1564 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7490
timestamp 1682952543
transform 1 0 1572 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7464
timestamp 1682952543
transform 1 0 1628 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7364
timestamp 1682952543
transform 1 0 1620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7365
timestamp 1682952543
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7465
timestamp 1682952543
transform 1 0 1692 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7484
timestamp 1682952543
transform 1 0 1676 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7543
timestamp 1682952543
transform 1 0 1668 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7485
timestamp 1682952543
transform 1 0 1716 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7366
timestamp 1682952543
transform 1 0 1676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7367
timestamp 1682952543
transform 1 0 1692 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7368
timestamp 1682952543
transform 1 0 1708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7369
timestamp 1682952543
transform 1 0 1716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7491
timestamp 1682952543
transform 1 0 1652 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7580
timestamp 1682952543
transform 1 0 1660 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7492
timestamp 1682952543
transform 1 0 1668 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7493
timestamp 1682952543
transform 1 0 1684 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7581
timestamp 1682952543
transform 1 0 1692 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7544
timestamp 1682952543
transform 1 0 1724 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7370
timestamp 1682952543
transform 1 0 1732 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7545
timestamp 1682952543
transform 1 0 1740 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7466
timestamp 1682952543
transform 1 0 1764 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7486
timestamp 1682952543
transform 1 0 1780 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7371
timestamp 1682952543
transform 1 0 1748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7372
timestamp 1682952543
transform 1 0 1756 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7546
timestamp 1682952543
transform 1 0 1764 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7373
timestamp 1682952543
transform 1 0 1772 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7547
timestamp 1682952543
transform 1 0 1780 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7487
timestamp 1682952543
transform 1 0 1828 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7374
timestamp 1682952543
transform 1 0 1788 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7375
timestamp 1682952543
transform 1 0 1796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7376
timestamp 1682952543
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7494
timestamp 1682952543
transform 1 0 1700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7495
timestamp 1682952543
transform 1 0 1708 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7496
timestamp 1682952543
transform 1 0 1740 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7647
timestamp 1682952543
transform 1 0 1700 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7582
timestamp 1682952543
transform 1 0 1748 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7548
timestamp 1682952543
transform 1 0 1844 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7497
timestamp 1682952543
transform 1 0 1756 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7498
timestamp 1682952543
transform 1 0 1764 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7499
timestamp 1682952543
transform 1 0 1788 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7500
timestamp 1682952543
transform 1 0 1876 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7648
timestamp 1682952543
transform 1 0 1740 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7649
timestamp 1682952543
transform 1 0 1764 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7650
timestamp 1682952543
transform 1 0 1796 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7377
timestamp 1682952543
transform 1 0 1916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7378
timestamp 1682952543
transform 1 0 1924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7310
timestamp 1682952543
transform 1 0 1956 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7501
timestamp 1682952543
transform 1 0 1948 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7502
timestamp 1682952543
transform 1 0 1988 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7488
timestamp 1682952543
transform 1 0 2052 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7489
timestamp 1682952543
transform 1 0 2092 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7442
timestamp 1682952543
transform 1 0 2148 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7467
timestamp 1682952543
transform 1 0 2116 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7516
timestamp 1682952543
transform 1 0 2108 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7490
timestamp 1682952543
transform 1 0 2140 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7379
timestamp 1682952543
transform 1 0 2052 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7380
timestamp 1682952543
transform 1 0 2084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7381
timestamp 1682952543
transform 1 0 2092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7382
timestamp 1682952543
transform 1 0 2108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7383
timestamp 1682952543
transform 1 0 2124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7384
timestamp 1682952543
transform 1 0 2140 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7503
timestamp 1682952543
transform 1 0 2004 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7583
timestamp 1682952543
transform 1 0 2044 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7504
timestamp 1682952543
transform 1 0 2108 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7505
timestamp 1682952543
transform 1 0 2116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7506
timestamp 1682952543
transform 1 0 2132 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7618
timestamp 1682952543
transform 1 0 2092 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7651
timestamp 1682952543
transform 1 0 2004 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7652
timestamp 1682952543
transform 1 0 2084 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7584
timestamp 1682952543
transform 1 0 2148 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7443
timestamp 1682952543
transform 1 0 2180 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7517
timestamp 1682952543
transform 1 0 2172 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7385
timestamp 1682952543
transform 1 0 2164 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7386
timestamp 1682952543
transform 1 0 2172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7387
timestamp 1682952543
transform 1 0 2188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7507
timestamp 1682952543
transform 1 0 2156 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7653
timestamp 1682952543
transform 1 0 2132 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7549
timestamp 1682952543
transform 1 0 2196 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7388
timestamp 1682952543
transform 1 0 2204 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7389
timestamp 1682952543
transform 1 0 2212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7508
timestamp 1682952543
transform 1 0 2172 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7654
timestamp 1682952543
transform 1 0 2164 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7655
timestamp 1682952543
transform 1 0 2188 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7656
timestamp 1682952543
transform 1 0 2204 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7619
timestamp 1682952543
transform 1 0 2228 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7444
timestamp 1682952543
transform 1 0 2244 0 1 1065
box -3 -3 3 3
use M2_M1  M2_M1_7509
timestamp 1682952543
transform 1 0 2244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7390
timestamp 1682952543
transform 1 0 2268 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7311
timestamp 1682952543
transform 1 0 2276 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7391
timestamp 1682952543
transform 1 0 2284 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7585
timestamp 1682952543
transform 1 0 2284 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7392
timestamp 1682952543
transform 1 0 2308 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7657
timestamp 1682952543
transform 1 0 2292 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7510
timestamp 1682952543
transform 1 0 2316 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7550
timestamp 1682952543
transform 1 0 2348 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7393
timestamp 1682952543
transform 1 0 2356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7511
timestamp 1682952543
transform 1 0 2348 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7394
timestamp 1682952543
transform 1 0 2380 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7518
timestamp 1682952543
transform 1 0 2412 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7395
timestamp 1682952543
transform 1 0 2404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7396
timestamp 1682952543
transform 1 0 2412 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7397
timestamp 1682952543
transform 1 0 2428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7398
timestamp 1682952543
transform 1 0 2444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7512
timestamp 1682952543
transform 1 0 2388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7513
timestamp 1682952543
transform 1 0 2396 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7658
timestamp 1682952543
transform 1 0 2380 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7586
timestamp 1682952543
transform 1 0 2404 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7514
timestamp 1682952543
transform 1 0 2412 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7587
timestamp 1682952543
transform 1 0 2428 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7620
timestamp 1682952543
transform 1 0 2444 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7659
timestamp 1682952543
transform 1 0 2436 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7519
timestamp 1682952543
transform 1 0 2460 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7450
timestamp 1682952543
transform 1 0 2484 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7468
timestamp 1682952543
transform 1 0 2500 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7520
timestamp 1682952543
transform 1 0 2484 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7551
timestamp 1682952543
transform 1 0 2476 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7491
timestamp 1682952543
transform 1 0 2540 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7399
timestamp 1682952543
transform 1 0 2484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7400
timestamp 1682952543
transform 1 0 2500 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7401
timestamp 1682952543
transform 1 0 2508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7402
timestamp 1682952543
transform 1 0 2524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7403
timestamp 1682952543
transform 1 0 2540 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7404
timestamp 1682952543
transform 1 0 2548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7515
timestamp 1682952543
transform 1 0 2468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7516
timestamp 1682952543
transform 1 0 2476 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7660
timestamp 1682952543
transform 1 0 2460 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7588
timestamp 1682952543
transform 1 0 2508 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7517
timestamp 1682952543
transform 1 0 2516 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7621
timestamp 1682952543
transform 1 0 2500 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7622
timestamp 1682952543
transform 1 0 2516 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7405
timestamp 1682952543
transform 1 0 2572 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7518
timestamp 1682952543
transform 1 0 2580 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7661
timestamp 1682952543
transform 1 0 2580 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7406
timestamp 1682952543
transform 1 0 2604 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7492
timestamp 1682952543
transform 1 0 2620 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7552
timestamp 1682952543
transform 1 0 2620 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7493
timestamp 1682952543
transform 1 0 2644 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7494
timestamp 1682952543
transform 1 0 2660 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7407
timestamp 1682952543
transform 1 0 2628 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7408
timestamp 1682952543
transform 1 0 2644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7409
timestamp 1682952543
transform 1 0 2652 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7519
timestamp 1682952543
transform 1 0 2612 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7520
timestamp 1682952543
transform 1 0 2620 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7589
timestamp 1682952543
transform 1 0 2652 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7451
timestamp 1682952543
transform 1 0 2676 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7623
timestamp 1682952543
transform 1 0 2668 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7452
timestamp 1682952543
transform 1 0 2692 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7562
timestamp 1682952543
transform 1 0 2700 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_7662
timestamp 1682952543
transform 1 0 2700 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7469
timestamp 1682952543
transform 1 0 2724 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7521
timestamp 1682952543
transform 1 0 2716 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7553
timestamp 1682952543
transform 1 0 2732 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7453
timestamp 1682952543
transform 1 0 2764 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7521
timestamp 1682952543
transform 1 0 2756 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7410
timestamp 1682952543
transform 1 0 2740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7522
timestamp 1682952543
transform 1 0 2732 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7522
timestamp 1682952543
transform 1 0 2780 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7411
timestamp 1682952543
transform 1 0 2764 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7554
timestamp 1682952543
transform 1 0 2772 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7412
timestamp 1682952543
transform 1 0 2780 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7413
timestamp 1682952543
transform 1 0 2796 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7414
timestamp 1682952543
transform 1 0 2804 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7523
timestamp 1682952543
transform 1 0 2772 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7624
timestamp 1682952543
transform 1 0 2780 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7663
timestamp 1682952543
transform 1 0 2796 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7523
timestamp 1682952543
transform 1 0 2820 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7415
timestamp 1682952543
transform 1 0 2836 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7555
timestamp 1682952543
transform 1 0 2844 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7524
timestamp 1682952543
transform 1 0 2812 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7525
timestamp 1682952543
transform 1 0 2828 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7590
timestamp 1682952543
transform 1 0 2836 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7526
timestamp 1682952543
transform 1 0 2844 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7625
timestamp 1682952543
transform 1 0 2820 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7664
timestamp 1682952543
transform 1 0 2844 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7556
timestamp 1682952543
transform 1 0 2860 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7470
timestamp 1682952543
transform 1 0 2876 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7524
timestamp 1682952543
transform 1 0 2908 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7557
timestamp 1682952543
transform 1 0 2876 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7416
timestamp 1682952543
transform 1 0 2924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7527
timestamp 1682952543
transform 1 0 2876 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7591
timestamp 1682952543
transform 1 0 2900 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7592
timestamp 1682952543
transform 1 0 2924 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7626
timestamp 1682952543
transform 1 0 2892 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7495
timestamp 1682952543
transform 1 0 2972 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7665
timestamp 1682952543
transform 1 0 2876 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7666
timestamp 1682952543
transform 1 0 2916 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7667
timestamp 1682952543
transform 1 0 2964 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7417
timestamp 1682952543
transform 1 0 2980 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7593
timestamp 1682952543
transform 1 0 2988 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7454
timestamp 1682952543
transform 1 0 3036 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7525
timestamp 1682952543
transform 1 0 3020 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7526
timestamp 1682952543
transform 1 0 3076 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7418
timestamp 1682952543
transform 1 0 3012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7419
timestamp 1682952543
transform 1 0 3028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7420
timestamp 1682952543
transform 1 0 3044 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7421
timestamp 1682952543
transform 1 0 3076 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7528
timestamp 1682952543
transform 1 0 2996 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7529
timestamp 1682952543
transform 1 0 3004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7530
timestamp 1682952543
transform 1 0 3020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7531
timestamp 1682952543
transform 1 0 3036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7532
timestamp 1682952543
transform 1 0 3124 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7627
timestamp 1682952543
transform 1 0 3012 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7668
timestamp 1682952543
transform 1 0 3020 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7628
timestamp 1682952543
transform 1 0 3084 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7445
timestamp 1682952543
transform 1 0 3196 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7558
timestamp 1682952543
transform 1 0 3148 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7422
timestamp 1682952543
transform 1 0 3196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7423
timestamp 1682952543
transform 1 0 3228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7424
timestamp 1682952543
transform 1 0 3236 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7425
timestamp 1682952543
transform 1 0 3244 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7533
timestamp 1682952543
transform 1 0 3148 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7594
timestamp 1682952543
transform 1 0 3196 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7595
timestamp 1682952543
transform 1 0 3236 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7534
timestamp 1682952543
transform 1 0 3244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7426
timestamp 1682952543
transform 1 0 3276 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7596
timestamp 1682952543
transform 1 0 3260 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7597
timestamp 1682952543
transform 1 0 3276 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7427
timestamp 1682952543
transform 1 0 3308 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7471
timestamp 1682952543
transform 1 0 3356 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7496
timestamp 1682952543
transform 1 0 3332 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7559
timestamp 1682952543
transform 1 0 3324 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7428
timestamp 1682952543
transform 1 0 3332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7429
timestamp 1682952543
transform 1 0 3348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7535
timestamp 1682952543
transform 1 0 3316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7536
timestamp 1682952543
transform 1 0 3324 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7629
timestamp 1682952543
transform 1 0 3316 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7669
timestamp 1682952543
transform 1 0 3308 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7598
timestamp 1682952543
transform 1 0 3332 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7537
timestamp 1682952543
transform 1 0 3340 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7599
timestamp 1682952543
transform 1 0 3348 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7455
timestamp 1682952543
transform 1 0 3380 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7527
timestamp 1682952543
transform 1 0 3396 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7560
timestamp 1682952543
transform 1 0 3364 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7430
timestamp 1682952543
transform 1 0 3380 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7561
timestamp 1682952543
transform 1 0 3388 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7431
timestamp 1682952543
transform 1 0 3396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7538
timestamp 1682952543
transform 1 0 3356 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7539
timestamp 1682952543
transform 1 0 3372 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7540
timestamp 1682952543
transform 1 0 3388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7432
timestamp 1682952543
transform 1 0 3412 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7541
timestamp 1682952543
transform 1 0 3420 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7670
timestamp 1682952543
transform 1 0 3412 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7528
timestamp 1682952543
transform 1 0 3476 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7433
timestamp 1682952543
transform 1 0 3460 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7562
timestamp 1682952543
transform 1 0 3468 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7600
timestamp 1682952543
transform 1 0 3460 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7542
timestamp 1682952543
transform 1 0 3508 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7630
timestamp 1682952543
transform 1 0 3428 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7631
timestamp 1682952543
transform 1 0 3508 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7671
timestamp 1682952543
transform 1 0 3436 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7529
timestamp 1682952543
transform 1 0 3524 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7434
timestamp 1682952543
transform 1 0 3524 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7601
timestamp 1682952543
transform 1 0 3532 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7497
timestamp 1682952543
transform 1 0 3548 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7435
timestamp 1682952543
transform 1 0 3548 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7632
timestamp 1682952543
transform 1 0 3548 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7456
timestamp 1682952543
transform 1 0 3572 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7530
timestamp 1682952543
transform 1 0 3596 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7436
timestamp 1682952543
transform 1 0 3596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7543
timestamp 1682952543
transform 1 0 3564 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7544
timestamp 1682952543
transform 1 0 3572 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7545
timestamp 1682952543
transform 1 0 3588 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7672
timestamp 1682952543
transform 1 0 3564 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7602
timestamp 1682952543
transform 1 0 3596 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7633
timestamp 1682952543
transform 1 0 3588 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7673
timestamp 1682952543
transform 1 0 3588 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7472
timestamp 1682952543
transform 1 0 3612 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7563
timestamp 1682952543
transform 1 0 3612 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7546
timestamp 1682952543
transform 1 0 3612 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7457
timestamp 1682952543
transform 1 0 3628 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7458
timestamp 1682952543
transform 1 0 3676 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7473
timestamp 1682952543
transform 1 0 3636 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_7498
timestamp 1682952543
transform 1 0 3716 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7499
timestamp 1682952543
transform 1 0 3764 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_7531
timestamp 1682952543
transform 1 0 3732 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7437
timestamp 1682952543
transform 1 0 3660 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7564
timestamp 1682952543
transform 1 0 3724 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7547
timestamp 1682952543
transform 1 0 3636 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7634
timestamp 1682952543
transform 1 0 3660 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7674
timestamp 1682952543
transform 1 0 3628 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7675
timestamp 1682952543
transform 1 0 3668 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7676
timestamp 1682952543
transform 1 0 3684 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7438
timestamp 1682952543
transform 1 0 3732 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7565
timestamp 1682952543
transform 1 0 3740 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7439
timestamp 1682952543
transform 1 0 3748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7440
timestamp 1682952543
transform 1 0 3764 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7603
timestamp 1682952543
transform 1 0 3732 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7459
timestamp 1682952543
transform 1 0 3788 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7460
timestamp 1682952543
transform 1 0 3860 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_7474
timestamp 1682952543
transform 1 0 3788 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7441
timestamp 1682952543
transform 1 0 3812 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7548
timestamp 1682952543
transform 1 0 3740 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7549
timestamp 1682952543
transform 1 0 3756 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7550
timestamp 1682952543
transform 1 0 3772 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7551
timestamp 1682952543
transform 1 0 3788 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7635
timestamp 1682952543
transform 1 0 3756 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7677
timestamp 1682952543
transform 1 0 3756 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7636
timestamp 1682952543
transform 1 0 3812 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7442
timestamp 1682952543
transform 1 0 3884 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7443
timestamp 1682952543
transform 1 0 3948 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7566
timestamp 1682952543
transform 1 0 3964 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7552
timestamp 1682952543
transform 1 0 3900 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7532
timestamp 1682952543
transform 1 0 4028 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7444
timestamp 1682952543
transform 1 0 3996 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7567
timestamp 1682952543
transform 1 0 4004 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7445
timestamp 1682952543
transform 1 0 4012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7446
timestamp 1682952543
transform 1 0 4028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7447
timestamp 1682952543
transform 1 0 4076 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7553
timestamp 1682952543
transform 1 0 4004 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7554
timestamp 1682952543
transform 1 0 4020 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7555
timestamp 1682952543
transform 1 0 4036 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7556
timestamp 1682952543
transform 1 0 4052 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7637
timestamp 1682952543
transform 1 0 4020 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7638
timestamp 1682952543
transform 1 0 4076 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7533
timestamp 1682952543
transform 1 0 4148 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7448
timestamp 1682952543
transform 1 0 4148 0 1 1015
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_62
timestamp 1682952543
transform 1 0 48 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_7678
timestamp 1682952543
transform 1 0 108 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7679
timestamp 1682952543
transform 1 0 148 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_464
timestamp 1682952543
transform 1 0 72 0 1 970
box -8 -3 104 105
use INVX2  INVX2_522
timestamp 1682952543
transform -1 0 184 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_298
timestamp 1682952543
transform 1 0 184 0 1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_466
timestamp 1682952543
transform 1 0 224 0 1 970
box -8 -3 104 105
use AOI22X1  AOI22X1_299
timestamp 1682952543
transform 1 0 320 0 1 970
box -8 -3 46 105
use OAI22X1  OAI22X1_327
timestamp 1682952543
transform 1 0 360 0 1 970
box -8 -3 46 105
use BUFX2  BUFX2_99
timestamp 1682952543
transform -1 0 424 0 1 970
box -5 -3 28 105
use M3_M2  M3_M2_7680
timestamp 1682952543
transform 1 0 436 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_467
timestamp 1682952543
transform 1 0 424 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_7681
timestamp 1682952543
transform 1 0 532 0 1 975
box -3 -3 3 3
use INVX2  INVX2_523
timestamp 1682952543
transform -1 0 536 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_300
timestamp 1682952543
transform 1 0 536 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_301
timestamp 1682952543
transform -1 0 616 0 1 970
box -8 -3 46 105
use AND2X2  AND2X2_54
timestamp 1682952543
transform -1 0 648 0 1 970
box -8 -3 40 105
use NOR2X1  NOR2X1_90
timestamp 1682952543
transform 1 0 648 0 1 970
box -8 -3 32 105
use FILL  FILL_3305
timestamp 1682952543
transform 1 0 672 0 1 970
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1682952543
transform 1 0 680 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_126
timestamp 1682952543
transform -1 0 720 0 1 970
box -8 -3 34 105
use FILL  FILL_3307
timestamp 1682952543
transform 1 0 720 0 1 970
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1682952543
transform 1 0 728 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_305
timestamp 1682952543
transform 1 0 736 0 1 970
box -8 -3 46 105
use FILL  FILL_3333
timestamp 1682952543
transform 1 0 776 0 1 970
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1682952543
transform 1 0 784 0 1 970
box -8 -3 16 105
use FILL  FILL_3339
timestamp 1682952543
transform 1 0 792 0 1 970
box -8 -3 16 105
use INVX2  INVX2_529
timestamp 1682952543
transform 1 0 800 0 1 970
box -9 -3 26 105
use FILL  FILL_3340
timestamp 1682952543
transform 1 0 816 0 1 970
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1682952543
transform 1 0 824 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7682
timestamp 1682952543
transform 1 0 844 0 1 975
box -3 -3 3 3
use FILL  FILL_3344
timestamp 1682952543
transform 1 0 832 0 1 970
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1682952543
transform 1 0 840 0 1 970
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1682952543
transform 1 0 848 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7683
timestamp 1682952543
transform 1 0 868 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_306
timestamp 1682952543
transform 1 0 856 0 1 970
box -8 -3 46 105
use FILL  FILL_3350
timestamp 1682952543
transform 1 0 896 0 1 970
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1682952543
transform 1 0 904 0 1 970
box -8 -3 16 105
use INVX2  INVX2_530
timestamp 1682952543
transform 1 0 912 0 1 970
box -9 -3 26 105
use FILL  FILL_3354
timestamp 1682952543
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1682952543
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1682952543
transform 1 0 944 0 1 970
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1682952543
transform 1 0 952 0 1 970
box -8 -3 16 105
use INVX2  INVX2_531
timestamp 1682952543
transform 1 0 960 0 1 970
box -9 -3 26 105
use FILL  FILL_3358
timestamp 1682952543
transform 1 0 976 0 1 970
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1682952543
transform 1 0 984 0 1 970
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1682952543
transform 1 0 992 0 1 970
box -8 -3 16 105
use FILL  FILL_3361
timestamp 1682952543
transform 1 0 1000 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_127
timestamp 1682952543
transform -1 0 1040 0 1 970
box -8 -3 34 105
use M3_M2  M3_M2_7684
timestamp 1682952543
transform 1 0 1068 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_308
timestamp 1682952543
transform -1 0 1080 0 1 970
box -8 -3 46 105
use FILL  FILL_3362
timestamp 1682952543
transform 1 0 1080 0 1 970
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1682952543
transform 1 0 1088 0 1 970
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1682952543
transform 1 0 1096 0 1 970
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1682952543
transform 1 0 1104 0 1 970
box -8 -3 16 105
use INVX2  INVX2_533
timestamp 1682952543
transform 1 0 1112 0 1 970
box -9 -3 26 105
use FILL  FILL_3378
timestamp 1682952543
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1682952543
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1682952543
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1682952543
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1682952543
transform 1 0 1160 0 1 970
box -8 -3 16 105
use FILL  FILL_3386
timestamp 1682952543
transform 1 0 1168 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_130
timestamp 1682952543
transform -1 0 1208 0 1 970
box -8 -3 34 105
use FILL  FILL_3387
timestamp 1682952543
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1682952543
transform 1 0 1216 0 1 970
box -8 -3 16 105
use INVX2  INVX2_534
timestamp 1682952543
transform 1 0 1224 0 1 970
box -9 -3 26 105
use FILL  FILL_3389
timestamp 1682952543
transform 1 0 1240 0 1 970
box -8 -3 16 105
use INVX2  INVX2_535
timestamp 1682952543
transform -1 0 1264 0 1 970
box -9 -3 26 105
use M3_M2  M3_M2_7685
timestamp 1682952543
transform 1 0 1276 0 1 975
box -3 -3 3 3
use FILL  FILL_3390
timestamp 1682952543
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1682952543
transform 1 0 1272 0 1 970
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1682952543
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1682952543
transform 1 0 1288 0 1 970
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1682952543
transform 1 0 1296 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_55
timestamp 1682952543
transform 1 0 1304 0 1 970
box -8 -3 40 105
use M3_M2  M3_M2_7686
timestamp 1682952543
transform 1 0 1348 0 1 975
box -3 -3 3 3
use FILL  FILL_3395
timestamp 1682952543
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_3396
timestamp 1682952543
transform 1 0 1344 0 1 970
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1682952543
transform 1 0 1352 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_470
timestamp 1682952543
transform 1 0 1360 0 1 970
box -8 -3 104 105
use BUFX2  BUFX2_100
timestamp 1682952543
transform -1 0 1480 0 1 970
box -5 -3 28 105
use FILL  FILL_3404
timestamp 1682952543
transform 1 0 1480 0 1 970
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1682952543
transform 1 0 1488 0 1 970
box -8 -3 16 105
use INVX2  INVX2_537
timestamp 1682952543
transform 1 0 1496 0 1 970
box -9 -3 26 105
use FILL  FILL_3406
timestamp 1682952543
transform 1 0 1512 0 1 970
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1682952543
transform 1 0 1520 0 1 970
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1682952543
transform 1 0 1528 0 1 970
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1682952543
transform 1 0 1536 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_309
timestamp 1682952543
transform -1 0 1584 0 1 970
box -8 -3 46 105
use FILL  FILL_3410
timestamp 1682952543
transform 1 0 1584 0 1 970
box -8 -3 16 105
use FILL  FILL_3411
timestamp 1682952543
transform 1 0 1592 0 1 970
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1682952543
transform 1 0 1600 0 1 970
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1682952543
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1682952543
transform 1 0 1616 0 1 970
box -8 -3 16 105
use INVX2  INVX2_538
timestamp 1682952543
transform -1 0 1640 0 1 970
box -9 -3 26 105
use FILL  FILL_3415
timestamp 1682952543
transform 1 0 1640 0 1 970
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1682952543
transform 1 0 1648 0 1 970
box -8 -3 16 105
use INVX2  INVX2_539
timestamp 1682952543
transform -1 0 1672 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_310
timestamp 1682952543
transform -1 0 1712 0 1 970
box -8 -3 46 105
use AOI22X1  AOI22X1_311
timestamp 1682952543
transform -1 0 1752 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_7687
timestamp 1682952543
transform 1 0 1772 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7688
timestamp 1682952543
transform 1 0 1788 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_312
timestamp 1682952543
transform 1 0 1752 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_7689
timestamp 1682952543
transform 1 0 1812 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_471
timestamp 1682952543
transform -1 0 1888 0 1 970
box -8 -3 104 105
use FILL  FILL_3417
timestamp 1682952543
transform 1 0 1888 0 1 970
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1682952543
transform 1 0 1896 0 1 970
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1682952543
transform 1 0 1904 0 1 970
box -8 -3 16 105
use INVX2  INVX2_540
timestamp 1682952543
transform -1 0 1928 0 1 970
box -9 -3 26 105
use FILL  FILL_3420
timestamp 1682952543
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_3421
timestamp 1682952543
transform 1 0 1936 0 1 970
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1682952543
transform 1 0 1944 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_64
timestamp 1682952543
transform -1 0 1976 0 1 970
box -8 -3 32 105
use M3_M2  M3_M2_7690
timestamp 1682952543
transform 1 0 1988 0 1 975
box -3 -3 3 3
use FILL  FILL_3423
timestamp 1682952543
transform 1 0 1976 0 1 970
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1682952543
transform 1 0 1984 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7691
timestamp 1682952543
transform 1 0 2076 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_472
timestamp 1682952543
transform 1 0 1992 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_7692
timestamp 1682952543
transform 1 0 2100 0 1 975
box -3 -3 3 3
use INVX2  INVX2_541
timestamp 1682952543
transform -1 0 2104 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_313
timestamp 1682952543
transform 1 0 2104 0 1 970
box -8 -3 46 105
use INVX2  INVX2_542
timestamp 1682952543
transform -1 0 2160 0 1 970
box -9 -3 26 105
use FILL  FILL_3425
timestamp 1682952543
transform 1 0 2160 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_314
timestamp 1682952543
transform 1 0 2168 0 1 970
box -8 -3 46 105
use FILL  FILL_3426
timestamp 1682952543
transform 1 0 2208 0 1 970
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1682952543
transform 1 0 2216 0 1 970
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1682952543
transform 1 0 2224 0 1 970
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1682952543
transform 1 0 2232 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7693
timestamp 1682952543
transform 1 0 2268 0 1 975
box -3 -3 3 3
use OAI21X1  OAI21X1_131
timestamp 1682952543
transform 1 0 2240 0 1 970
box -8 -3 34 105
use FILL  FILL_3430
timestamp 1682952543
transform 1 0 2272 0 1 970
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1682952543
transform 1 0 2280 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7694
timestamp 1682952543
transform 1 0 2308 0 1 975
box -3 -3 3 3
use AND2X2  AND2X2_56
timestamp 1682952543
transform -1 0 2320 0 1 970
box -8 -3 40 105
use FILL  FILL_3432
timestamp 1682952543
transform 1 0 2320 0 1 970
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1682952543
transform 1 0 2328 0 1 970
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1682952543
transform 1 0 2336 0 1 970
box -8 -3 16 105
use FILL  FILL_3435
timestamp 1682952543
transform 1 0 2344 0 1 970
box -8 -3 16 105
use FILL  FILL_3436
timestamp 1682952543
transform 1 0 2352 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_57
timestamp 1682952543
transform -1 0 2392 0 1 970
box -8 -3 40 105
use M3_M2  M3_M2_7695
timestamp 1682952543
transform 1 0 2404 0 1 975
box -3 -3 3 3
use INVX2  INVX2_543
timestamp 1682952543
transform 1 0 2392 0 1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_315
timestamp 1682952543
transform 1 0 2408 0 1 970
box -8 -3 46 105
use FILL  FILL_3437
timestamp 1682952543
transform 1 0 2448 0 1 970
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1682952543
transform 1 0 2456 0 1 970
box -8 -3 16 105
use FILL  FILL_3439
timestamp 1682952543
transform 1 0 2464 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_58
timestamp 1682952543
transform 1 0 2472 0 1 970
box -8 -3 40 105
use AOI22X1  AOI22X1_318
timestamp 1682952543
transform 1 0 2504 0 1 970
box -8 -3 46 105
use FILL  FILL_3463
timestamp 1682952543
transform 1 0 2544 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7696
timestamp 1682952543
transform 1 0 2564 0 1 975
box -3 -3 3 3
use FILL  FILL_3468
timestamp 1682952543
transform 1 0 2552 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_335
timestamp 1682952543
transform -1 0 2600 0 1 970
box -8 -3 46 105
use FILL  FILL_3469
timestamp 1682952543
transform 1 0 2600 0 1 970
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1682952543
transform 1 0 2608 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7697
timestamp 1682952543
transform 1 0 2628 0 1 975
box -3 -3 3 3
use AND2X2  AND2X2_59
timestamp 1682952543
transform 1 0 2616 0 1 970
box -8 -3 40 105
use FILL  FILL_3474
timestamp 1682952543
transform 1 0 2648 0 1 970
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1682952543
transform 1 0 2656 0 1 970
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1682952543
transform 1 0 2664 0 1 970
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1682952543
transform 1 0 2672 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7698
timestamp 1682952543
transform 1 0 2708 0 1 975
box -3 -3 3 3
use NOR2X1  NOR2X1_94
timestamp 1682952543
transform -1 0 2704 0 1 970
box -8 -3 32 105
use FILL  FILL_3478
timestamp 1682952543
transform 1 0 2704 0 1 970
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1682952543
transform 1 0 2712 0 1 970
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1682952543
transform 1 0 2720 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7699
timestamp 1682952543
transform 1 0 2740 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7700
timestamp 1682952543
transform 1 0 2764 0 1 975
box -3 -3 3 3
use AND2X2  AND2X2_60
timestamp 1682952543
transform 1 0 2728 0 1 970
box -8 -3 40 105
use FILL  FILL_3481
timestamp 1682952543
transform 1 0 2760 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_61
timestamp 1682952543
transform 1 0 2768 0 1 970
box -8 -3 40 105
use FILL  FILL_3482
timestamp 1682952543
transform 1 0 2800 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7701
timestamp 1682952543
transform 1 0 2836 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_336
timestamp 1682952543
transform 1 0 2808 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_7702
timestamp 1682952543
transform 1 0 2860 0 1 975
box -3 -3 3 3
use FILL  FILL_3483
timestamp 1682952543
transform 1 0 2848 0 1 970
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1682952543
transform 1 0 2856 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_480
timestamp 1682952543
transform 1 0 2864 0 1 970
box -8 -3 104 105
use INVX2  INVX2_550
timestamp 1682952543
transform 1 0 2960 0 1 970
box -9 -3 26 105
use FILL  FILL_3489
timestamp 1682952543
transform 1 0 2976 0 1 970
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1682952543
transform 1 0 2984 0 1 970
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1682952543
transform 1 0 2992 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_338
timestamp 1682952543
transform 1 0 3000 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_7703
timestamp 1682952543
transform 1 0 3084 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_481
timestamp 1682952543
transform -1 0 3136 0 1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_482
timestamp 1682952543
transform 1 0 3136 0 1 970
box -8 -3 104 105
use FILL  FILL_3492
timestamp 1682952543
transform 1 0 3232 0 1 970
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1682952543
transform 1 0 3240 0 1 970
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1682952543
transform 1 0 3248 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_321
timestamp 1682952543
transform -1 0 3296 0 1 970
box -8 -3 46 105
use FILL  FILL_3495
timestamp 1682952543
transform 1 0 3296 0 1 970
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1682952543
transform 1 0 3304 0 1 970
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1682952543
transform 1 0 3312 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7704
timestamp 1682952543
transform 1 0 3340 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_339
timestamp 1682952543
transform 1 0 3320 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_7705
timestamp 1682952543
transform 1 0 3380 0 1 975
box -3 -3 3 3
use FILL  FILL_3498
timestamp 1682952543
transform 1 0 3360 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_340
timestamp 1682952543
transform 1 0 3368 0 1 970
box -8 -3 46 105
use FILL  FILL_3499
timestamp 1682952543
transform 1 0 3408 0 1 970
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1682952543
transform 1 0 3416 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7706
timestamp 1682952543
transform 1 0 3436 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_483
timestamp 1682952543
transform -1 0 3520 0 1 970
box -8 -3 104 105
use FILL  FILL_3501
timestamp 1682952543
transform 1 0 3520 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7707
timestamp 1682952543
transform 1 0 3540 0 1 975
box -3 -3 3 3
use FILL  FILL_3502
timestamp 1682952543
transform 1 0 3528 0 1 970
box -8 -3 16 105
use INVX2  INVX2_551
timestamp 1682952543
transform -1 0 3552 0 1 970
box -9 -3 26 105
use FILL  FILL_3503
timestamp 1682952543
transform 1 0 3552 0 1 970
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1682952543
transform 1 0 3560 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7708
timestamp 1682952543
transform 1 0 3580 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_341
timestamp 1682952543
transform 1 0 3568 0 1 970
box -8 -3 46 105
use FILL  FILL_3505
timestamp 1682952543
transform 1 0 3608 0 1 970
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1682952543
transform 1 0 3616 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_484
timestamp 1682952543
transform 1 0 3624 0 1 970
box -8 -3 104 105
use INVX2  INVX2_552
timestamp 1682952543
transform 1 0 3720 0 1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_342
timestamp 1682952543
transform -1 0 3776 0 1 970
box -8 -3 46 105
use M3_M2  M3_M2_7709
timestamp 1682952543
transform 1 0 3796 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7710
timestamp 1682952543
transform 1 0 3820 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_485
timestamp 1682952543
transform 1 0 3776 0 1 970
box -8 -3 104 105
use INVX2  INVX2_553
timestamp 1682952543
transform 1 0 3872 0 1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_486
timestamp 1682952543
transform 1 0 3888 0 1 970
box -8 -3 104 105
use INVX2  INVX2_554
timestamp 1682952543
transform 1 0 3984 0 1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_343
timestamp 1682952543
transform 1 0 4000 0 1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_490
timestamp 1682952543
transform 1 0 4040 0 1 970
box -8 -3 104 105
use INVX2  INVX2_563
timestamp 1682952543
transform 1 0 4136 0 1 970
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_63
timestamp 1682952543
transform 1 0 4177 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_7761
timestamp 1682952543
transform 1 0 84 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7762
timestamp 1682952543
transform 1 0 108 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7739
timestamp 1682952543
transform 1 0 212 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7763
timestamp 1682952543
transform 1 0 188 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7566
timestamp 1682952543
transform 1 0 84 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7792
timestamp 1682952543
transform 1 0 164 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7567
timestamp 1682952543
transform 1 0 180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7568
timestamp 1682952543
transform 1 0 188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7569
timestamp 1682952543
transform 1 0 196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7685
timestamp 1682952543
transform 1 0 132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7686
timestamp 1682952543
transform 1 0 164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7687
timestamp 1682952543
transform 1 0 172 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7858
timestamp 1682952543
transform 1 0 132 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7793
timestamp 1682952543
transform 1 0 204 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7570
timestamp 1682952543
transform 1 0 212 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7571
timestamp 1682952543
transform 1 0 220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7688
timestamp 1682952543
transform 1 0 204 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7824
timestamp 1682952543
transform 1 0 212 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7689
timestamp 1682952543
transform 1 0 220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7690
timestamp 1682952543
transform 1 0 228 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7572
timestamp 1682952543
transform 1 0 236 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7825
timestamp 1682952543
transform 1 0 236 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7859
timestamp 1682952543
transform 1 0 228 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7573
timestamp 1682952543
transform 1 0 252 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7826
timestamp 1682952543
transform 1 0 252 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7574
timestamp 1682952543
transform 1 0 268 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7691
timestamp 1682952543
transform 1 0 260 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7764
timestamp 1682952543
transform 1 0 292 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7794
timestamp 1682952543
transform 1 0 284 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7765
timestamp 1682952543
transform 1 0 324 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7575
timestamp 1682952543
transform 1 0 292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7576
timestamp 1682952543
transform 1 0 316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7692
timestamp 1682952543
transform 1 0 284 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7827
timestamp 1682952543
transform 1 0 292 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7693
timestamp 1682952543
transform 1 0 300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7694
timestamp 1682952543
transform 1 0 316 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7828
timestamp 1682952543
transform 1 0 332 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7711
timestamp 1682952543
transform 1 0 356 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7740
timestamp 1682952543
transform 1 0 372 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7795
timestamp 1682952543
transform 1 0 348 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7577
timestamp 1682952543
transform 1 0 356 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7796
timestamp 1682952543
transform 1 0 364 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7578
timestamp 1682952543
transform 1 0 372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7695
timestamp 1682952543
transform 1 0 340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7696
timestamp 1682952543
transform 1 0 348 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7829
timestamp 1682952543
transform 1 0 356 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7697
timestamp 1682952543
transform 1 0 364 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7830
timestamp 1682952543
transform 1 0 372 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7860
timestamp 1682952543
transform 1 0 340 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7911
timestamp 1682952543
transform 1 0 356 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7698
timestamp 1682952543
transform 1 0 388 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7861
timestamp 1682952543
transform 1 0 396 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7831
timestamp 1682952543
transform 1 0 412 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7898
timestamp 1682952543
transform 1 0 412 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7912
timestamp 1682952543
transform 1 0 404 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7699
timestamp 1682952543
transform 1 0 428 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7862
timestamp 1682952543
transform 1 0 428 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7863
timestamp 1682952543
transform 1 0 452 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7913
timestamp 1682952543
transform 1 0 452 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7741
timestamp 1682952543
transform 1 0 508 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7766
timestamp 1682952543
transform 1 0 500 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7579
timestamp 1682952543
transform 1 0 476 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7580
timestamp 1682952543
transform 1 0 484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7581
timestamp 1682952543
transform 1 0 500 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7700
timestamp 1682952543
transform 1 0 468 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7832
timestamp 1682952543
transform 1 0 484 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7701
timestamp 1682952543
transform 1 0 492 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7742
timestamp 1682952543
transform 1 0 540 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7743
timestamp 1682952543
transform 1 0 556 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7582
timestamp 1682952543
transform 1 0 532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7702
timestamp 1682952543
transform 1 0 524 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7833
timestamp 1682952543
transform 1 0 532 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7767
timestamp 1682952543
transform 1 0 572 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7583
timestamp 1682952543
transform 1 0 556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7584
timestamp 1682952543
transform 1 0 572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7703
timestamp 1682952543
transform 1 0 540 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7864
timestamp 1682952543
transform 1 0 524 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7834
timestamp 1682952543
transform 1 0 556 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7704
timestamp 1682952543
transform 1 0 564 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7865
timestamp 1682952543
transform 1 0 564 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7797
timestamp 1682952543
transform 1 0 588 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7835
timestamp 1682952543
transform 1 0 580 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7585
timestamp 1682952543
transform 1 0 596 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7768
timestamp 1682952543
transform 1 0 612 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7705
timestamp 1682952543
transform 1 0 620 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7866
timestamp 1682952543
transform 1 0 620 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7586
timestamp 1682952543
transform 1 0 636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7706
timestamp 1682952543
transform 1 0 660 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7867
timestamp 1682952543
transform 1 0 660 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7914
timestamp 1682952543
transform 1 0 636 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7712
timestamp 1682952543
transform 1 0 724 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7563
timestamp 1682952543
transform 1 0 724 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7798
timestamp 1682952543
transform 1 0 724 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7707
timestamp 1682952543
transform 1 0 724 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7744
timestamp 1682952543
transform 1 0 764 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7564
timestamp 1682952543
transform 1 0 764 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_7587
timestamp 1682952543
transform 1 0 796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7708
timestamp 1682952543
transform 1 0 796 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7931
timestamp 1682952543
transform 1 0 796 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7588
timestamp 1682952543
transform 1 0 812 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7769
timestamp 1682952543
transform 1 0 852 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7589
timestamp 1682952543
transform 1 0 868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7709
timestamp 1682952543
transform 1 0 852 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7710
timestamp 1682952543
transform 1 0 860 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7711
timestamp 1682952543
transform 1 0 876 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7712
timestamp 1682952543
transform 1 0 892 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7915
timestamp 1682952543
transform 1 0 860 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7932
timestamp 1682952543
transform 1 0 876 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7590
timestamp 1682952543
transform 1 0 908 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7770
timestamp 1682952543
transform 1 0 956 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7591
timestamp 1682952543
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7713
timestamp 1682952543
transform 1 0 932 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7714
timestamp 1682952543
transform 1 0 940 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7868
timestamp 1682952543
transform 1 0 924 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7933
timestamp 1682952543
transform 1 0 924 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7869
timestamp 1682952543
transform 1 0 940 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7810
timestamp 1682952543
transform 1 0 956 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7565
timestamp 1682952543
transform 1 0 964 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7916
timestamp 1682952543
transform 1 0 972 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7592
timestamp 1682952543
transform 1 0 988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7715
timestamp 1682952543
transform 1 0 996 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7593
timestamp 1682952543
transform 1 0 1012 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7771
timestamp 1682952543
transform 1 0 1020 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7799
timestamp 1682952543
transform 1 0 1036 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7716
timestamp 1682952543
transform 1 0 1036 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7811
timestamp 1682952543
transform 1 0 1020 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7594
timestamp 1682952543
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7836
timestamp 1682952543
transform 1 0 1068 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7713
timestamp 1682952543
transform 1 0 1076 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7595
timestamp 1682952543
transform 1 0 1076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7717
timestamp 1682952543
transform 1 0 1092 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7772
timestamp 1682952543
transform 1 0 1124 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7800
timestamp 1682952543
transform 1 0 1132 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7718
timestamp 1682952543
transform 1 0 1124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7719
timestamp 1682952543
transform 1 0 1132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7812
timestamp 1682952543
transform 1 0 1148 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7934
timestamp 1682952543
transform 1 0 1164 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7917
timestamp 1682952543
transform 1 0 1180 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7714
timestamp 1682952543
transform 1 0 1196 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7715
timestamp 1682952543
transform 1 0 1220 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7596
timestamp 1682952543
transform 1 0 1196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7597
timestamp 1682952543
transform 1 0 1204 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7870
timestamp 1682952543
transform 1 0 1196 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7801
timestamp 1682952543
transform 1 0 1212 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7598
timestamp 1682952543
transform 1 0 1220 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7802
timestamp 1682952543
transform 1 0 1228 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7599
timestamp 1682952543
transform 1 0 1236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7720
timestamp 1682952543
transform 1 0 1212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7721
timestamp 1682952543
transform 1 0 1228 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7722
timestamp 1682952543
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7871
timestamp 1682952543
transform 1 0 1236 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7837
timestamp 1682952543
transform 1 0 1252 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7773
timestamp 1682952543
transform 1 0 1292 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7803
timestamp 1682952543
transform 1 0 1292 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7600
timestamp 1682952543
transform 1 0 1340 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7723
timestamp 1682952543
transform 1 0 1292 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7918
timestamp 1682952543
transform 1 0 1340 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7601
timestamp 1682952543
transform 1 0 1356 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7716
timestamp 1682952543
transform 1 0 1380 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7602
timestamp 1682952543
transform 1 0 1388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7724
timestamp 1682952543
transform 1 0 1380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7725
timestamp 1682952543
transform 1 0 1396 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7717
timestamp 1682952543
transform 1 0 1412 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7726
timestamp 1682952543
transform 1 0 1412 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7745
timestamp 1682952543
transform 1 0 1436 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7603
timestamp 1682952543
transform 1 0 1428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7604
timestamp 1682952543
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7919
timestamp 1682952543
transform 1 0 1444 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7718
timestamp 1682952543
transform 1 0 1468 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7746
timestamp 1682952543
transform 1 0 1460 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7719
timestamp 1682952543
transform 1 0 1492 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7605
timestamp 1682952543
transform 1 0 1484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7727
timestamp 1682952543
transform 1 0 1516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7728
timestamp 1682952543
transform 1 0 1564 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7720
timestamp 1682952543
transform 1 0 1588 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7721
timestamp 1682952543
transform 1 0 1644 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7747
timestamp 1682952543
transform 1 0 1604 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7748
timestamp 1682952543
transform 1 0 1652 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7606
timestamp 1682952543
transform 1 0 1588 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7729
timestamp 1682952543
transform 1 0 1636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7607
timestamp 1682952543
transform 1 0 1676 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7749
timestamp 1682952543
transform 1 0 1708 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7730
timestamp 1682952543
transform 1 0 1708 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7750
timestamp 1682952543
transform 1 0 1756 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7804
timestamp 1682952543
transform 1 0 1732 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7608
timestamp 1682952543
transform 1 0 1740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7609
timestamp 1682952543
transform 1 0 1756 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7731
timestamp 1682952543
transform 1 0 1732 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7732
timestamp 1682952543
transform 1 0 1748 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7899
timestamp 1682952543
transform 1 0 1748 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7751
timestamp 1682952543
transform 1 0 1772 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7900
timestamp 1682952543
transform 1 0 1764 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7610
timestamp 1682952543
transform 1 0 1780 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7872
timestamp 1682952543
transform 1 0 1780 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7611
timestamp 1682952543
transform 1 0 1796 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7805
timestamp 1682952543
transform 1 0 1804 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7733
timestamp 1682952543
transform 1 0 1804 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7734
timestamp 1682952543
transform 1 0 1812 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7901
timestamp 1682952543
transform 1 0 1804 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7838
timestamp 1682952543
transform 1 0 1820 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7735
timestamp 1682952543
transform 1 0 1828 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7736
timestamp 1682952543
transform 1 0 1844 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7873
timestamp 1682952543
transform 1 0 1828 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7902
timestamp 1682952543
transform 1 0 1820 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7903
timestamp 1682952543
transform 1 0 1844 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7935
timestamp 1682952543
transform 1 0 1836 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7612
timestamp 1682952543
transform 1 0 1860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7613
timestamp 1682952543
transform 1 0 1876 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7806
timestamp 1682952543
transform 1 0 1948 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7839
timestamp 1682952543
transform 1 0 1908 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7737
timestamp 1682952543
transform 1 0 1916 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7840
timestamp 1682952543
transform 1 0 1940 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7722
timestamp 1682952543
transform 1 0 2004 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7614
timestamp 1682952543
transform 1 0 1972 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7807
timestamp 1682952543
transform 1 0 1980 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7615
timestamp 1682952543
transform 1 0 1988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7616
timestamp 1682952543
transform 1 0 1996 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7752
timestamp 1682952543
transform 1 0 2044 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7753
timestamp 1682952543
transform 1 0 2068 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7617
timestamp 1682952543
transform 1 0 2028 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7618
timestamp 1682952543
transform 1 0 2036 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7808
timestamp 1682952543
transform 1 0 2044 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7619
timestamp 1682952543
transform 1 0 2052 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7620
timestamp 1682952543
transform 1 0 2068 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7621
timestamp 1682952543
transform 1 0 2076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7738
timestamp 1682952543
transform 1 0 1956 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7739
timestamp 1682952543
transform 1 0 1964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7740
timestamp 1682952543
transform 1 0 1980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7741
timestamp 1682952543
transform 1 0 1996 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7742
timestamp 1682952543
transform 1 0 2012 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7874
timestamp 1682952543
transform 1 0 1924 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7875
timestamp 1682952543
transform 1 0 1948 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7876
timestamp 1682952543
transform 1 0 1988 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7877
timestamp 1682952543
transform 1 0 2004 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7904
timestamp 1682952543
transform 1 0 1964 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7936
timestamp 1682952543
transform 1 0 1932 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7841
timestamp 1682952543
transform 1 0 2028 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7743
timestamp 1682952543
transform 1 0 2044 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7744
timestamp 1682952543
transform 1 0 2060 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7842
timestamp 1682952543
transform 1 0 2068 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7813
timestamp 1682952543
transform 1 0 2028 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7937
timestamp 1682952543
transform 1 0 2012 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7878
timestamp 1682952543
transform 1 0 2044 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7622
timestamp 1682952543
transform 1 0 2100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7745
timestamp 1682952543
transform 1 0 2092 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7746
timestamp 1682952543
transform 1 0 2100 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7879
timestamp 1682952543
transform 1 0 2100 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7754
timestamp 1682952543
transform 1 0 2116 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7905
timestamp 1682952543
transform 1 0 2108 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7723
timestamp 1682952543
transform 1 0 2172 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7623
timestamp 1682952543
transform 1 0 2132 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7624
timestamp 1682952543
transform 1 0 2148 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7625
timestamp 1682952543
transform 1 0 2164 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7626
timestamp 1682952543
transform 1 0 2252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7747
timestamp 1682952543
transform 1 0 2124 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7748
timestamp 1682952543
transform 1 0 2140 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7843
timestamp 1682952543
transform 1 0 2148 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7844
timestamp 1682952543
transform 1 0 2164 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7724
timestamp 1682952543
transform 1 0 2356 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7774
timestamp 1682952543
transform 1 0 2332 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7725
timestamp 1682952543
transform 1 0 2412 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7775
timestamp 1682952543
transform 1 0 2404 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7627
timestamp 1682952543
transform 1 0 2276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7628
timestamp 1682952543
transform 1 0 2292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7749
timestamp 1682952543
transform 1 0 2188 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7750
timestamp 1682952543
transform 1 0 2244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7751
timestamp 1682952543
transform 1 0 2260 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7880
timestamp 1682952543
transform 1 0 2140 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7881
timestamp 1682952543
transform 1 0 2252 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7809
timestamp 1682952543
transform 1 0 2340 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7810
timestamp 1682952543
transform 1 0 2372 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7629
timestamp 1682952543
transform 1 0 2388 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7845
timestamp 1682952543
transform 1 0 2292 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7752
timestamp 1682952543
transform 1 0 2324 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7753
timestamp 1682952543
transform 1 0 2372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7814
timestamp 1682952543
transform 1 0 2276 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7906
timestamp 1682952543
transform 1 0 2260 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7938
timestamp 1682952543
transform 1 0 2212 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7939
timestamp 1682952543
transform 1 0 2252 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7907
timestamp 1682952543
transform 1 0 2356 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7940
timestamp 1682952543
transform 1 0 2300 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7846
timestamp 1682952543
transform 1 0 2388 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7726
timestamp 1682952543
transform 1 0 2500 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7754
timestamp 1682952543
transform 1 0 2436 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7755
timestamp 1682952543
transform 1 0 2468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7756
timestamp 1682952543
transform 1 0 2484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7630
timestamp 1682952543
transform 1 0 2508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7757
timestamp 1682952543
transform 1 0 2516 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7815
timestamp 1682952543
transform 1 0 2508 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7941
timestamp 1682952543
transform 1 0 2540 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7811
timestamp 1682952543
transform 1 0 2548 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7727
timestamp 1682952543
transform 1 0 2588 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7728
timestamp 1682952543
transform 1 0 2604 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7631
timestamp 1682952543
transform 1 0 2564 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7812
timestamp 1682952543
transform 1 0 2572 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7632
timestamp 1682952543
transform 1 0 2580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7633
timestamp 1682952543
transform 1 0 2596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7634
timestamp 1682952543
transform 1 0 2604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7758
timestamp 1682952543
transform 1 0 2572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7759
timestamp 1682952543
transform 1 0 2588 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7882
timestamp 1682952543
transform 1 0 2564 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7847
timestamp 1682952543
transform 1 0 2596 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7883
timestamp 1682952543
transform 1 0 2588 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7942
timestamp 1682952543
transform 1 0 2572 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7729
timestamp 1682952543
transform 1 0 2620 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7848
timestamp 1682952543
transform 1 0 2612 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7730
timestamp 1682952543
transform 1 0 2700 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7755
timestamp 1682952543
transform 1 0 2668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7756
timestamp 1682952543
transform 1 0 2716 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7776
timestamp 1682952543
transform 1 0 2708 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7777
timestamp 1682952543
transform 1 0 2732 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7731
timestamp 1682952543
transform 1 0 2788 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7778
timestamp 1682952543
transform 1 0 2772 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7813
timestamp 1682952543
transform 1 0 2684 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7814
timestamp 1682952543
transform 1 0 2708 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7635
timestamp 1682952543
transform 1 0 2732 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7815
timestamp 1682952543
transform 1 0 2748 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7636
timestamp 1682952543
transform 1 0 2756 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7816
timestamp 1682952543
transform 1 0 2764 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7779
timestamp 1682952543
transform 1 0 2804 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7637
timestamp 1682952543
transform 1 0 2780 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7638
timestamp 1682952543
transform 1 0 2788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7639
timestamp 1682952543
transform 1 0 2804 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7760
timestamp 1682952543
transform 1 0 2636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7761
timestamp 1682952543
transform 1 0 2644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7762
timestamp 1682952543
transform 1 0 2652 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7849
timestamp 1682952543
transform 1 0 2660 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7763
timestamp 1682952543
transform 1 0 2684 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7850
timestamp 1682952543
transform 1 0 2732 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7764
timestamp 1682952543
transform 1 0 2748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7765
timestamp 1682952543
transform 1 0 2764 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7766
timestamp 1682952543
transform 1 0 2780 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7884
timestamp 1682952543
transform 1 0 2644 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7885
timestamp 1682952543
transform 1 0 2684 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7920
timestamp 1682952543
transform 1 0 2668 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7921
timestamp 1682952543
transform 1 0 2684 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7922
timestamp 1682952543
transform 1 0 2708 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7943
timestamp 1682952543
transform 1 0 2636 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7944
timestamp 1682952543
transform 1 0 2660 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7945
timestamp 1682952543
transform 1 0 2748 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7851
timestamp 1682952543
transform 1 0 2788 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7780
timestamp 1682952543
transform 1 0 2828 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7640
timestamp 1682952543
transform 1 0 2828 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7767
timestamp 1682952543
transform 1 0 2796 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7768
timestamp 1682952543
transform 1 0 2812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7769
timestamp 1682952543
transform 1 0 2820 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7886
timestamp 1682952543
transform 1 0 2796 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7887
timestamp 1682952543
transform 1 0 2820 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7923
timestamp 1682952543
transform 1 0 2812 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7946
timestamp 1682952543
transform 1 0 2812 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7852
timestamp 1682952543
transform 1 0 2844 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7770
timestamp 1682952543
transform 1 0 2852 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7947
timestamp 1682952543
transform 1 0 2836 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7641
timestamp 1682952543
transform 1 0 2860 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7781
timestamp 1682952543
transform 1 0 2924 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7642
timestamp 1682952543
transform 1 0 2948 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7771
timestamp 1682952543
transform 1 0 2900 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7924
timestamp 1682952543
transform 1 0 2868 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7643
timestamp 1682952543
transform 1 0 2972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7644
timestamp 1682952543
transform 1 0 2988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7645
timestamp 1682952543
transform 1 0 3004 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7646
timestamp 1682952543
transform 1 0 3012 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7772
timestamp 1682952543
transform 1 0 2980 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7773
timestamp 1682952543
transform 1 0 2996 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7732
timestamp 1682952543
transform 1 0 3028 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7774
timestamp 1682952543
transform 1 0 3020 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7733
timestamp 1682952543
transform 1 0 3044 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7782
timestamp 1682952543
transform 1 0 3076 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7647
timestamp 1682952543
transform 1 0 3036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7648
timestamp 1682952543
transform 1 0 3044 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7817
timestamp 1682952543
transform 1 0 3052 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7649
timestamp 1682952543
transform 1 0 3060 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7818
timestamp 1682952543
transform 1 0 3068 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7650
timestamp 1682952543
transform 1 0 3076 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7775
timestamp 1682952543
transform 1 0 3052 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7776
timestamp 1682952543
transform 1 0 3068 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7888
timestamp 1682952543
transform 1 0 3052 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7777
timestamp 1682952543
transform 1 0 3084 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7783
timestamp 1682952543
transform 1 0 3180 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7651
timestamp 1682952543
transform 1 0 3108 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7819
timestamp 1682952543
transform 1 0 3132 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7778
timestamp 1682952543
transform 1 0 3132 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7853
timestamp 1682952543
transform 1 0 3196 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7652
timestamp 1682952543
transform 1 0 3220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7779
timestamp 1682952543
transform 1 0 3204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7780
timestamp 1682952543
transform 1 0 3212 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7948
timestamp 1682952543
transform 1 0 3116 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7949
timestamp 1682952543
transform 1 0 3188 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7820
timestamp 1682952543
transform 1 0 3228 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7653
timestamp 1682952543
transform 1 0 3236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7654
timestamp 1682952543
transform 1 0 3252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7655
timestamp 1682952543
transform 1 0 3260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7781
timestamp 1682952543
transform 1 0 3244 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7784
timestamp 1682952543
transform 1 0 3308 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7656
timestamp 1682952543
transform 1 0 3276 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7657
timestamp 1682952543
transform 1 0 3292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7658
timestamp 1682952543
transform 1 0 3308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7782
timestamp 1682952543
transform 1 0 3268 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7783
timestamp 1682952543
transform 1 0 3276 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7784
timestamp 1682952543
transform 1 0 3300 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7785
timestamp 1682952543
transform 1 0 3316 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7925
timestamp 1682952543
transform 1 0 3284 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7926
timestamp 1682952543
transform 1 0 3308 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7734
timestamp 1682952543
transform 1 0 3324 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7785
timestamp 1682952543
transform 1 0 3324 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7735
timestamp 1682952543
transform 1 0 3372 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7786
timestamp 1682952543
transform 1 0 3364 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7659
timestamp 1682952543
transform 1 0 3324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7660
timestamp 1682952543
transform 1 0 3332 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7661
timestamp 1682952543
transform 1 0 3348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7662
timestamp 1682952543
transform 1 0 3364 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7821
timestamp 1682952543
transform 1 0 3372 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7786
timestamp 1682952543
transform 1 0 3340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7787
timestamp 1682952543
transform 1 0 3356 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7788
timestamp 1682952543
transform 1 0 3372 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7822
timestamp 1682952543
transform 1 0 3388 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7736
timestamp 1682952543
transform 1 0 3404 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7737
timestamp 1682952543
transform 1 0 3436 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7787
timestamp 1682952543
transform 1 0 3420 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7663
timestamp 1682952543
transform 1 0 3396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7664
timestamp 1682952543
transform 1 0 3404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7665
timestamp 1682952543
transform 1 0 3420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7666
timestamp 1682952543
transform 1 0 3436 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7854
timestamp 1682952543
transform 1 0 3396 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7789
timestamp 1682952543
transform 1 0 3404 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7855
timestamp 1682952543
transform 1 0 3412 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7790
timestamp 1682952543
transform 1 0 3428 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7950
timestamp 1682952543
transform 1 0 3420 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7791
timestamp 1682952543
transform 1 0 3444 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7927
timestamp 1682952543
transform 1 0 3468 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7951
timestamp 1682952543
transform 1 0 3476 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7667
timestamp 1682952543
transform 1 0 3492 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7889
timestamp 1682952543
transform 1 0 3492 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7928
timestamp 1682952543
transform 1 0 3492 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7668
timestamp 1682952543
transform 1 0 3508 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7823
timestamp 1682952543
transform 1 0 3532 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7792
timestamp 1682952543
transform 1 0 3532 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7793
timestamp 1682952543
transform 1 0 3588 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7890
timestamp 1682952543
transform 1 0 3532 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7816
timestamp 1682952543
transform 1 0 3596 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7757
timestamp 1682952543
transform 1 0 3612 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7669
timestamp 1682952543
transform 1 0 3636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7817
timestamp 1682952543
transform 1 0 3628 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7891
timestamp 1682952543
transform 1 0 3636 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7819
timestamp 1682952543
transform 1 0 3612 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_7820
timestamp 1682952543
transform 1 0 3628 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_7952
timestamp 1682952543
transform 1 0 3604 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7929
timestamp 1682952543
transform 1 0 3628 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7953
timestamp 1682952543
transform 1 0 3636 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7758
timestamp 1682952543
transform 1 0 3668 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7788
timestamp 1682952543
transform 1 0 3660 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7789
timestamp 1682952543
transform 1 0 3684 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7670
timestamp 1682952543
transform 1 0 3660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7671
timestamp 1682952543
transform 1 0 3668 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7672
timestamp 1682952543
transform 1 0 3684 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7794
timestamp 1682952543
transform 1 0 3660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7795
timestamp 1682952543
transform 1 0 3676 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7892
timestamp 1682952543
transform 1 0 3676 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7954
timestamp 1682952543
transform 1 0 3660 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7673
timestamp 1682952543
transform 1 0 3708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7796
timestamp 1682952543
transform 1 0 3700 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7908
timestamp 1682952543
transform 1 0 3700 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7955
timestamp 1682952543
transform 1 0 3692 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7759
timestamp 1682952543
transform 1 0 3724 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7674
timestamp 1682952543
transform 1 0 3740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7797
timestamp 1682952543
transform 1 0 3716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7798
timestamp 1682952543
transform 1 0 3732 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7675
timestamp 1682952543
transform 1 0 3772 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7799
timestamp 1682952543
transform 1 0 3764 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7818
timestamp 1682952543
transform 1 0 3772 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7956
timestamp 1682952543
transform 1 0 3772 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7738
timestamp 1682952543
transform 1 0 3820 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7790
timestamp 1682952543
transform 1 0 3820 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7676
timestamp 1682952543
transform 1 0 3788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7677
timestamp 1682952543
transform 1 0 3804 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7678
timestamp 1682952543
transform 1 0 3820 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7679
timestamp 1682952543
transform 1 0 3828 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7856
timestamp 1682952543
transform 1 0 3788 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7800
timestamp 1682952543
transform 1 0 3812 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7909
timestamp 1682952543
transform 1 0 3812 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7801
timestamp 1682952543
transform 1 0 3836 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7893
timestamp 1682952543
transform 1 0 3828 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7910
timestamp 1682952543
transform 1 0 3836 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7760
timestamp 1682952543
transform 1 0 3884 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7802
timestamp 1682952543
transform 1 0 3868 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7803
timestamp 1682952543
transform 1 0 3884 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7804
timestamp 1682952543
transform 1 0 3892 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7930
timestamp 1682952543
transform 1 0 3868 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7894
timestamp 1682952543
transform 1 0 3892 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7680
timestamp 1682952543
transform 1 0 3916 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7895
timestamp 1682952543
transform 1 0 3916 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7791
timestamp 1682952543
transform 1 0 3932 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7681
timestamp 1682952543
transform 1 0 3980 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7805
timestamp 1682952543
transform 1 0 3972 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7857
timestamp 1682952543
transform 1 0 3980 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7682
timestamp 1682952543
transform 1 0 4004 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7683
timestamp 1682952543
transform 1 0 4020 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7684
timestamp 1682952543
transform 1 0 4036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7806
timestamp 1682952543
transform 1 0 4004 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7807
timestamp 1682952543
transform 1 0 4028 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7896
timestamp 1682952543
transform 1 0 4028 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7808
timestamp 1682952543
transform 1 0 4044 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7897
timestamp 1682952543
transform 1 0 4044 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7809
timestamp 1682952543
transform 1 0 4124 0 1 925
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_64
timestamp 1682952543
transform 1 0 24 0 1 870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_465
timestamp 1682952543
transform 1 0 72 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_524
timestamp 1682952543
transform -1 0 184 0 -1 970
box -9 -3 26 105
use AOI22X1  AOI22X1_302
timestamp 1682952543
transform 1 0 184 0 -1 970
box -8 -3 46 105
use INVX2  INVX2_525
timestamp 1682952543
transform -1 0 240 0 -1 970
box -9 -3 26 105
use FILL  FILL_3308
timestamp 1682952543
transform 1 0 240 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_526
timestamp 1682952543
transform 1 0 248 0 -1 970
box -9 -3 26 105
use FILL  FILL_3309
timestamp 1682952543
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1682952543
transform 1 0 272 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_303
timestamp 1682952543
transform 1 0 280 0 -1 970
box -8 -3 46 105
use FILL  FILL_3311
timestamp 1682952543
transform 1 0 320 0 -1 970
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1682952543
transform 1 0 328 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_328
timestamp 1682952543
transform 1 0 336 0 -1 970
box -8 -3 46 105
use FILL  FILL_3313
timestamp 1682952543
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_3314
timestamp 1682952543
transform 1 0 384 0 -1 970
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1682952543
transform 1 0 392 0 -1 970
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1682952543
transform 1 0 400 0 -1 970
box -8 -3 16 105
use FILL  FILL_3317
timestamp 1682952543
transform 1 0 408 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_527
timestamp 1682952543
transform -1 0 432 0 -1 970
box -9 -3 26 105
use FILL  FILL_3318
timestamp 1682952543
transform 1 0 432 0 -1 970
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1682952543
transform 1 0 440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1682952543
transform 1 0 448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1682952543
transform 1 0 456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1682952543
transform 1 0 464 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_304
timestamp 1682952543
transform -1 0 512 0 -1 970
box -8 -3 46 105
use FILL  FILL_3323
timestamp 1682952543
transform 1 0 512 0 -1 970
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1682952543
transform 1 0 520 0 -1 970
box -8 -3 16 105
use FILL  FILL_3325
timestamp 1682952543
transform 1 0 528 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_329
timestamp 1682952543
transform 1 0 536 0 -1 970
box -8 -3 46 105
use FILL  FILL_3326
timestamp 1682952543
transform 1 0 576 0 -1 970
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1682952543
transform 1 0 584 0 -1 970
box -8 -3 16 105
use FILL  FILL_3328
timestamp 1682952543
transform 1 0 592 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_528
timestamp 1682952543
transform 1 0 600 0 -1 970
box -9 -3 26 105
use FILL  FILL_3329
timestamp 1682952543
transform 1 0 616 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_468
timestamp 1682952543
transform 1 0 624 0 -1 970
box -8 -3 104 105
use FILL  FILL_3330
timestamp 1682952543
transform 1 0 720 0 -1 970
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1682952543
transform 1 0 728 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_91
timestamp 1682952543
transform 1 0 736 0 -1 970
box -8 -3 32 105
use FILL  FILL_3334
timestamp 1682952543
transform 1 0 760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1682952543
transform 1 0 768 0 -1 970
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1682952543
transform 1 0 776 0 -1 970
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1682952543
transform 1 0 784 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7957
timestamp 1682952543
transform 1 0 820 0 1 875
box -3 -3 3 3
use NOR2X1  NOR2X1_92
timestamp 1682952543
transform 1 0 792 0 -1 970
box -8 -3 32 105
use FILL  FILL_3341
timestamp 1682952543
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1682952543
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3345
timestamp 1682952543
transform 1 0 832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1682952543
transform 1 0 840 0 -1 970
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1682952543
transform 1 0 848 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_307
timestamp 1682952543
transform 1 0 856 0 -1 970
box -8 -3 46 105
use FILL  FILL_3351
timestamp 1682952543
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3353
timestamp 1682952543
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1682952543
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1682952543
transform 1 0 920 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7958
timestamp 1682952543
transform 1 0 948 0 1 875
box -3 -3 3 3
use OAI21X1  OAI21X1_128
timestamp 1682952543
transform 1 0 928 0 -1 970
box -8 -3 34 105
use M3_M2  M3_M2_7959
timestamp 1682952543
transform 1 0 972 0 1 875
box -3 -3 3 3
use FILL  FILL_3367
timestamp 1682952543
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3368
timestamp 1682952543
transform 1 0 968 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_93
timestamp 1682952543
transform 1 0 976 0 -1 970
box -8 -3 32 105
use FILL  FILL_3369
timestamp 1682952543
transform 1 0 1000 0 -1 970
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1682952543
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_129
timestamp 1682952543
transform -1 0 1048 0 -1 970
box -8 -3 34 105
use FILL  FILL_3371
timestamp 1682952543
transform 1 0 1048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1682952543
transform 1 0 1056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1682952543
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_3374
timestamp 1682952543
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_532
timestamp 1682952543
transform 1 0 1080 0 -1 970
box -9 -3 26 105
use FILL  FILL_3375
timestamp 1682952543
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1682952543
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_63
timestamp 1682952543
transform 1 0 1112 0 -1 970
box -8 -3 32 105
use FILL  FILL_3380
timestamp 1682952543
transform 1 0 1136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1682952543
transform 1 0 1144 0 -1 970
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1682952543
transform 1 0 1152 0 -1 970
box -8 -3 16 105
use FILL  FILL_3398
timestamp 1682952543
transform 1 0 1160 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_536
timestamp 1682952543
transform -1 0 1184 0 -1 970
box -9 -3 26 105
use FILL  FILL_3399
timestamp 1682952543
transform 1 0 1184 0 -1 970
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1682952543
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_330
timestamp 1682952543
transform -1 0 1240 0 -1 970
box -8 -3 46 105
use FILL  FILL_3401
timestamp 1682952543
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7960
timestamp 1682952543
transform 1 0 1260 0 1 875
box -3 -3 3 3
use FILL  FILL_3402
timestamp 1682952543
transform 1 0 1248 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_469
timestamp 1682952543
transform -1 0 1352 0 -1 970
box -8 -3 104 105
use FILL  FILL_3403
timestamp 1682952543
transform 1 0 1352 0 -1 970
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1682952543
transform 1 0 1360 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_331
timestamp 1682952543
transform -1 0 1408 0 -1 970
box -8 -3 46 105
use FILL  FILL_3441
timestamp 1682952543
transform 1 0 1408 0 -1 970
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1682952543
transform 1 0 1416 0 -1 970
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1682952543
transform 1 0 1424 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_544
timestamp 1682952543
transform -1 0 1448 0 -1 970
box -9 -3 26 105
use FILL  FILL_3444
timestamp 1682952543
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1682952543
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1682952543
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_473
timestamp 1682952543
transform 1 0 1472 0 -1 970
box -8 -3 104 105
use FILL  FILL_3447
timestamp 1682952543
transform 1 0 1568 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_474
timestamp 1682952543
transform 1 0 1576 0 -1 970
box -8 -3 104 105
use FILL  FILL_3448
timestamp 1682952543
transform 1 0 1672 0 -1 970
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1682952543
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use FILL  FILL_3450
timestamp 1682952543
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1682952543
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1682952543
transform 1 0 1704 0 -1 970
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1682952543
transform 1 0 1712 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_332
timestamp 1682952543
transform 1 0 1720 0 -1 970
box -8 -3 46 105
use FILL  FILL_3454
timestamp 1682952543
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1682952543
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_545
timestamp 1682952543
transform 1 0 1776 0 -1 970
box -9 -3 26 105
use FILL  FILL_3456
timestamp 1682952543
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1682952543
transform 1 0 1800 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_316
timestamp 1682952543
transform 1 0 1808 0 -1 970
box -8 -3 46 105
use FILL  FILL_3458
timestamp 1682952543
transform 1 0 1848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1682952543
transform 1 0 1856 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_475
timestamp 1682952543
transform 1 0 1864 0 -1 970
box -8 -3 104 105
use AOI22X1  AOI22X1_317
timestamp 1682952543
transform -1 0 2000 0 -1 970
box -8 -3 46 105
use OAI21X1  OAI21X1_132
timestamp 1682952543
transform 1 0 2000 0 -1 970
box -8 -3 34 105
use OAI22X1  OAI22X1_333
timestamp 1682952543
transform 1 0 2032 0 -1 970
box -8 -3 46 105
use FILL  FILL_3460
timestamp 1682952543
transform 1 0 2072 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_546
timestamp 1682952543
transform 1 0 2080 0 -1 970
box -9 -3 26 105
use FILL  FILL_3461
timestamp 1682952543
transform 1 0 2096 0 -1 970
box -8 -3 16 105
use FILL  FILL_3462
timestamp 1682952543
transform 1 0 2104 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_334
timestamp 1682952543
transform 1 0 2112 0 -1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_476
timestamp 1682952543
transform 1 0 2152 0 -1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_133
timestamp 1682952543
transform 1 0 2248 0 -1 970
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_477
timestamp 1682952543
transform 1 0 2280 0 -1 970
box -8 -3 104 105
use M3_M2  M3_M2_7961
timestamp 1682952543
transform 1 0 2420 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_478
timestamp 1682952543
transform 1 0 2376 0 -1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_134
timestamp 1682952543
transform 1 0 2472 0 -1 970
box -8 -3 34 105
use FILL  FILL_3464
timestamp 1682952543
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1682952543
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_547
timestamp 1682952543
transform -1 0 2536 0 -1 970
box -9 -3 26 105
use FILL  FILL_3466
timestamp 1682952543
transform 1 0 2536 0 -1 970
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1682952543
transform 1 0 2544 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7962
timestamp 1682952543
transform 1 0 2564 0 1 875
box -3 -3 3 3
use FILL  FILL_3471
timestamp 1682952543
transform 1 0 2552 0 -1 970
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1682952543
transform 1 0 2560 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7963
timestamp 1682952543
transform 1 0 2580 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_319
timestamp 1682952543
transform 1 0 2568 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_7964
timestamp 1682952543
transform 1 0 2620 0 1 875
box -3 -3 3 3
use FILL  FILL_3473
timestamp 1682952543
transform 1 0 2608 0 -1 970
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1682952543
transform 1 0 2616 0 -1 970
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1682952543
transform 1 0 2624 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7965
timestamp 1682952543
transform 1 0 2652 0 1 875
box -3 -3 3 3
use INVX2  INVX2_548
timestamp 1682952543
transform 1 0 2632 0 -1 970
box -9 -3 26 105
use M3_M2  M3_M2_7966
timestamp 1682952543
transform 1 0 2668 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_479
timestamp 1682952543
transform -1 0 2744 0 -1 970
box -8 -3 104 105
use M3_M2  M3_M2_7967
timestamp 1682952543
transform 1 0 2780 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_320
timestamp 1682952543
transform 1 0 2744 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_7968
timestamp 1682952543
transform 1 0 2820 0 1 875
box -3 -3 3 3
use OAI22X1  OAI22X1_337
timestamp 1682952543
transform -1 0 2824 0 -1 970
box -8 -3 46 105
use FILL  FILL_3486
timestamp 1682952543
transform 1 0 2824 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_549
timestamp 1682952543
transform -1 0 2848 0 -1 970
box -9 -3 26 105
use FILL  FILL_3487
timestamp 1682952543
transform 1 0 2848 0 -1 970
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1682952543
transform 1 0 2856 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7969
timestamp 1682952543
transform 1 0 2908 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_487
timestamp 1682952543
transform -1 0 2960 0 -1 970
box -8 -3 104 105
use FILL  FILL_3508
timestamp 1682952543
transform 1 0 2960 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_344
timestamp 1682952543
transform -1 0 3008 0 -1 970
box -8 -3 46 105
use FILL  FILL_3509
timestamp 1682952543
transform 1 0 3008 0 -1 970
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1682952543
transform 1 0 3016 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_555
timestamp 1682952543
transform -1 0 3040 0 -1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_345
timestamp 1682952543
transform -1 0 3080 0 -1 970
box -8 -3 46 105
use FILL  FILL_3511
timestamp 1682952543
transform 1 0 3080 0 -1 970
box -8 -3 16 105
use FILL  FILL_3512
timestamp 1682952543
transform 1 0 3088 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_488
timestamp 1682952543
transform 1 0 3096 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_556
timestamp 1682952543
transform 1 0 3192 0 -1 970
box -9 -3 26 105
use FILL  FILL_3513
timestamp 1682952543
transform 1 0 3208 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_346
timestamp 1682952543
transform 1 0 3216 0 -1 970
box -8 -3 46 105
use M3_M2  M3_M2_7970
timestamp 1682952543
transform 1 0 3276 0 1 875
box -3 -3 3 3
use INVX2  INVX2_557
timestamp 1682952543
transform 1 0 3256 0 -1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_347
timestamp 1682952543
transform 1 0 3272 0 -1 970
box -8 -3 46 105
use INVX2  INVX2_558
timestamp 1682952543
transform -1 0 3328 0 -1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_348
timestamp 1682952543
transform 1 0 3328 0 -1 970
box -8 -3 46 105
use INVX2  INVX2_559
timestamp 1682952543
transform -1 0 3384 0 -1 970
box -9 -3 26 105
use FILL  FILL_3514
timestamp 1682952543
transform 1 0 3384 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7971
timestamp 1682952543
transform 1 0 3404 0 1 875
box -3 -3 3 3
use FILL  FILL_3515
timestamp 1682952543
transform 1 0 3392 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_349
timestamp 1682952543
transform 1 0 3400 0 -1 970
box -8 -3 46 105
use FILL  FILL_3516
timestamp 1682952543
transform 1 0 3440 0 -1 970
box -8 -3 16 105
use FILL  FILL_3517
timestamp 1682952543
transform 1 0 3448 0 -1 970
box -8 -3 16 105
use FILL  FILL_3518
timestamp 1682952543
transform 1 0 3456 0 -1 970
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1682952543
transform 1 0 3464 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_560
timestamp 1682952543
transform -1 0 3488 0 -1 970
box -9 -3 26 105
use FILL  FILL_3520
timestamp 1682952543
transform 1 0 3488 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7972
timestamp 1682952543
transform 1 0 3516 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_7973
timestamp 1682952543
transform 1 0 3556 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_489
timestamp 1682952543
transform 1 0 3496 0 -1 970
box -8 -3 104 105
use FILL  FILL_3521
timestamp 1682952543
transform 1 0 3592 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_65
timestamp 1682952543
transform -1 0 3632 0 -1 970
box -8 -3 40 105
use INVX2  INVX2_561
timestamp 1682952543
transform 1 0 3632 0 -1 970
box -9 -3 26 105
use FILL  FILL_3522
timestamp 1682952543
transform 1 0 3648 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7974
timestamp 1682952543
transform 1 0 3700 0 1 875
box -3 -3 3 3
use AOI22X1  AOI22X1_322
timestamp 1682952543
transform -1 0 3696 0 -1 970
box -8 -3 46 105
use FILL  FILL_3523
timestamp 1682952543
transform 1 0 3696 0 -1 970
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1682952543
transform 1 0 3704 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_323
timestamp 1682952543
transform 1 0 3712 0 -1 970
box -8 -3 46 105
use FILL  FILL_3525
timestamp 1682952543
transform 1 0 3752 0 -1 970
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1682952543
transform 1 0 3760 0 -1 970
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1682952543
transform 1 0 3768 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7975
timestamp 1682952543
transform 1 0 3788 0 1 875
box -3 -3 3 3
use FILL  FILL_3528
timestamp 1682952543
transform 1 0 3776 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_350
timestamp 1682952543
transform 1 0 3784 0 -1 970
box -8 -3 46 105
use FILL  FILL_3529
timestamp 1682952543
transform 1 0 3824 0 -1 970
box -8 -3 16 105
use FILL  FILL_3530
timestamp 1682952543
transform 1 0 3832 0 -1 970
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1682952543
transform 1 0 3840 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_324
timestamp 1682952543
transform 1 0 3848 0 -1 970
box -8 -3 46 105
use FILL  FILL_3532
timestamp 1682952543
transform 1 0 3888 0 -1 970
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1682952543
transform 1 0 3896 0 -1 970
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1682952543
transform 1 0 3904 0 -1 970
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1682952543
transform 1 0 3912 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_562
timestamp 1682952543
transform -1 0 3936 0 -1 970
box -9 -3 26 105
use FILL  FILL_3536
timestamp 1682952543
transform 1 0 3936 0 -1 970
box -8 -3 16 105
use FILL  FILL_3537
timestamp 1682952543
transform 1 0 3944 0 -1 970
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1682952543
transform 1 0 3952 0 -1 970
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1682952543
transform 1 0 3960 0 -1 970
box -8 -3 16 105
use FILL  FILL_3540
timestamp 1682952543
transform 1 0 3968 0 -1 970
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1682952543
transform 1 0 3976 0 -1 970
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1682952543
transform 1 0 3984 0 -1 970
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1682952543
transform 1 0 3992 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_351
timestamp 1682952543
transform 1 0 4000 0 -1 970
box -8 -3 46 105
use FILL  FILL_3544
timestamp 1682952543
transform 1 0 4040 0 -1 970
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1682952543
transform 1 0 4048 0 -1 970
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1682952543
transform 1 0 4056 0 -1 970
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1682952543
transform 1 0 4064 0 -1 970
box -8 -3 16 105
use FILL  FILL_3548
timestamp 1682952543
transform 1 0 4072 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_564
timestamp 1682952543
transform -1 0 4096 0 -1 970
box -9 -3 26 105
use FILL  FILL_3549
timestamp 1682952543
transform 1 0 4096 0 -1 970
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1682952543
transform 1 0 4104 0 -1 970
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1682952543
transform 1 0 4112 0 -1 970
box -8 -3 16 105
use FILL  FILL_3552
timestamp 1682952543
transform 1 0 4120 0 -1 970
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1682952543
transform 1 0 4128 0 -1 970
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1682952543
transform 1 0 4136 0 -1 970
box -8 -3 16 105
use FILL  FILL_3555
timestamp 1682952543
transform 1 0 4144 0 -1 970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_65
timestamp 1682952543
transform 1 0 4201 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_8035
timestamp 1682952543
transform 1 0 180 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8059
timestamp 1682952543
transform 1 0 132 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8060
timestamp 1682952543
transform 1 0 172 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8105
timestamp 1682952543
transform 1 0 84 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7837
timestamp 1682952543
transform 1 0 132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7838
timestamp 1682952543
transform 1 0 164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7839
timestamp 1682952543
transform 1 0 172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7840
timestamp 1682952543
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7961
timestamp 1682952543
transform 1 0 84 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8127
timestamp 1682952543
transform 1 0 164 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_7962
timestamp 1682952543
transform 1 0 180 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8128
timestamp 1682952543
transform 1 0 188 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_7963
timestamp 1682952543
transform 1 0 196 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8155
timestamp 1682952543
transform 1 0 204 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8036
timestamp 1682952543
transform 1 0 228 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7841
timestamp 1682952543
transform 1 0 220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7842
timestamp 1682952543
transform 1 0 228 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8037
timestamp 1682952543
transform 1 0 276 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7843
timestamp 1682952543
transform 1 0 260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7964
timestamp 1682952543
transform 1 0 252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7965
timestamp 1682952543
transform 1 0 276 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7995
timestamp 1682952543
transform 1 0 332 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_7844
timestamp 1682952543
transform 1 0 308 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7845
timestamp 1682952543
transform 1 0 316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7846
timestamp 1682952543
transform 1 0 332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7966
timestamp 1682952543
transform 1 0 324 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8129
timestamp 1682952543
transform 1 0 332 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7996
timestamp 1682952543
transform 1 0 364 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8061
timestamp 1682952543
transform 1 0 436 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8062
timestamp 1682952543
transform 1 0 484 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8063
timestamp 1682952543
transform 1 0 500 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8064
timestamp 1682952543
transform 1 0 540 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8106
timestamp 1682952543
transform 1 0 380 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7847
timestamp 1682952543
transform 1 0 388 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7848
timestamp 1682952543
transform 1 0 436 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7967
timestamp 1682952543
transform 1 0 340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7968
timestamp 1682952543
transform 1 0 356 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8107
timestamp 1682952543
transform 1 0 452 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7849
timestamp 1682952543
transform 1 0 500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7850
timestamp 1682952543
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7851
timestamp 1682952543
transform 1 0 540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7969
timestamp 1682952543
transform 1 0 452 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8156
timestamp 1682952543
transform 1 0 476 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8108
timestamp 1682952543
transform 1 0 548 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7852
timestamp 1682952543
transform 1 0 556 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8184
timestamp 1682952543
transform 1 0 524 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7997
timestamp 1682952543
transform 1 0 596 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8109
timestamp 1682952543
transform 1 0 572 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7853
timestamp 1682952543
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7854
timestamp 1682952543
transform 1 0 596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7970
timestamp 1682952543
transform 1 0 564 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7971
timestamp 1682952543
transform 1 0 572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7972
timestamp 1682952543
transform 1 0 588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8157
timestamp 1682952543
transform 1 0 588 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_7973
timestamp 1682952543
transform 1 0 604 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8065
timestamp 1682952543
transform 1 0 676 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8066
timestamp 1682952543
transform 1 0 716 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7855
timestamp 1682952543
transform 1 0 676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7856
timestamp 1682952543
transform 1 0 708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7857
timestamp 1682952543
transform 1 0 716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7974
timestamp 1682952543
transform 1 0 628 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8158
timestamp 1682952543
transform 1 0 628 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8159
timestamp 1682952543
transform 1 0 660 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8160
timestamp 1682952543
transform 1 0 708 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8038
timestamp 1682952543
transform 1 0 740 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7858
timestamp 1682952543
transform 1 0 740 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8110
timestamp 1682952543
transform 1 0 764 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7859
timestamp 1682952543
transform 1 0 772 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7860
timestamp 1682952543
transform 1 0 788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7975
timestamp 1682952543
transform 1 0 756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7976
timestamp 1682952543
transform 1 0 764 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7977
timestamp 1682952543
transform 1 0 780 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8161
timestamp 1682952543
transform 1 0 780 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8022
timestamp 1682952543
transform 1 0 820 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_7861
timestamp 1682952543
transform 1 0 804 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8111
timestamp 1682952543
transform 1 0 812 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7998
timestamp 1682952543
transform 1 0 852 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_7824
timestamp 1682952543
transform 1 0 852 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7862
timestamp 1682952543
transform 1 0 836 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8112
timestamp 1682952543
transform 1 0 852 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_8162
timestamp 1682952543
transform 1 0 852 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8067
timestamp 1682952543
transform 1 0 868 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7978
timestamp 1682952543
transform 1 0 868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8074
timestamp 1682952543
transform 1 0 868 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_8068
timestamp 1682952543
transform 1 0 892 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7863
timestamp 1682952543
transform 1 0 892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8075
timestamp 1682952543
transform 1 0 892 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_8185
timestamp 1682952543
transform 1 0 892 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_7979
timestamp 1682952543
transform 1 0 916 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7980
timestamp 1682952543
transform 1 0 924 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7981
timestamp 1682952543
transform 1 0 932 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7864
timestamp 1682952543
transform 1 0 948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7865
timestamp 1682952543
transform 1 0 972 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8163
timestamp 1682952543
transform 1 0 964 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8186
timestamp 1682952543
transform 1 0 964 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_7982
timestamp 1682952543
transform 1 0 996 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7825
timestamp 1682952543
transform 1 0 1012 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7826
timestamp 1682952543
transform 1 0 1020 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_8113
timestamp 1682952543
transform 1 0 1012 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7983
timestamp 1682952543
transform 1 0 1012 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8187
timestamp 1682952543
transform 1 0 1004 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_7866
timestamp 1682952543
transform 1 0 1036 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8069
timestamp 1682952543
transform 1 0 1060 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8070
timestamp 1682952543
transform 1 0 1100 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8071
timestamp 1682952543
transform 1 0 1156 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7867
timestamp 1682952543
transform 1 0 1100 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7984
timestamp 1682952543
transform 1 0 1076 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8130
timestamp 1682952543
transform 1 0 1084 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8114
timestamp 1682952543
transform 1 0 1116 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7868
timestamp 1682952543
transform 1 0 1156 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7999
timestamp 1682952543
transform 1 0 1228 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8072
timestamp 1682952543
transform 1 0 1212 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7869
timestamp 1682952543
transform 1 0 1204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7870
timestamp 1682952543
transform 1 0 1220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7985
timestamp 1682952543
transform 1 0 1092 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7986
timestamp 1682952543
transform 1 0 1180 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7987
timestamp 1682952543
transform 1 0 1196 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7988
timestamp 1682952543
transform 1 0 1212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7989
timestamp 1682952543
transform 1 0 1228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7990
timestamp 1682952543
transform 1 0 1236 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8164
timestamp 1682952543
transform 1 0 1220 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8188
timestamp 1682952543
transform 1 0 1196 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8189
timestamp 1682952543
transform 1 0 1236 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8000
timestamp 1682952543
transform 1 0 1268 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8073
timestamp 1682952543
transform 1 0 1252 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8074
timestamp 1682952543
transform 1 0 1276 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7871
timestamp 1682952543
transform 1 0 1252 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8115
timestamp 1682952543
transform 1 0 1260 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7872
timestamp 1682952543
transform 1 0 1268 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7873
timestamp 1682952543
transform 1 0 1276 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7991
timestamp 1682952543
transform 1 0 1260 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8165
timestamp 1682952543
transform 1 0 1268 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_7992
timestamp 1682952543
transform 1 0 1284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7874
timestamp 1682952543
transform 1 0 1300 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8131
timestamp 1682952543
transform 1 0 1300 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_7993
timestamp 1682952543
transform 1 0 1316 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8023
timestamp 1682952543
transform 1 0 1348 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_7994
timestamp 1682952543
transform 1 0 1332 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_7995
timestamp 1682952543
transform 1 0 1340 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8190
timestamp 1682952543
transform 1 0 1340 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8001
timestamp 1682952543
transform 1 0 1388 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_7875
timestamp 1682952543
transform 1 0 1364 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7876
timestamp 1682952543
transform 1 0 1380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7996
timestamp 1682952543
transform 1 0 1356 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8132
timestamp 1682952543
transform 1 0 1364 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_7997
timestamp 1682952543
transform 1 0 1372 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8166
timestamp 1682952543
transform 1 0 1380 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_7877
timestamp 1682952543
transform 1 0 1396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7998
timestamp 1682952543
transform 1 0 1404 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7976
timestamp 1682952543
transform 1 0 1452 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8002
timestamp 1682952543
transform 1 0 1436 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8024
timestamp 1682952543
transform 1 0 1420 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_8075
timestamp 1682952543
transform 1 0 1468 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8076
timestamp 1682952543
transform 1 0 1508 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7878
timestamp 1682952543
transform 1 0 1468 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8116
timestamp 1682952543
transform 1 0 1492 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7879
timestamp 1682952543
transform 1 0 1500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7880
timestamp 1682952543
transform 1 0 1508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7999
timestamp 1682952543
transform 1 0 1420 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8167
timestamp 1682952543
transform 1 0 1436 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8168
timestamp 1682952543
transform 1 0 1484 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8039
timestamp 1682952543
transform 1 0 1580 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7881
timestamp 1682952543
transform 1 0 1540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7882
timestamp 1682952543
transform 1 0 1548 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8117
timestamp 1682952543
transform 1 0 1556 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7883
timestamp 1682952543
transform 1 0 1564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7884
timestamp 1682952543
transform 1 0 1580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8000
timestamp 1682952543
transform 1 0 1548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8001
timestamp 1682952543
transform 1 0 1556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8002
timestamp 1682952543
transform 1 0 1572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8003
timestamp 1682952543
transform 1 0 1588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7977
timestamp 1682952543
transform 1 0 1692 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8003
timestamp 1682952543
transform 1 0 1612 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8004
timestamp 1682952543
transform 1 0 1668 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8077
timestamp 1682952543
transform 1 0 1684 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8078
timestamp 1682952543
transform 1 0 1716 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7885
timestamp 1682952543
transform 1 0 1636 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8118
timestamp 1682952543
transform 1 0 1676 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7827
timestamp 1682952543
transform 1 0 1732 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7886
timestamp 1682952543
transform 1 0 1684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7887
timestamp 1682952543
transform 1 0 1692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7888
timestamp 1682952543
transform 1 0 1708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7889
timestamp 1682952543
transform 1 0 1724 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8004
timestamp 1682952543
transform 1 0 1604 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8133
timestamp 1682952543
transform 1 0 1644 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8005
timestamp 1682952543
transform 1 0 1692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8006
timestamp 1682952543
transform 1 0 1700 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8134
timestamp 1682952543
transform 1 0 1708 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8007
timestamp 1682952543
transform 1 0 1716 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8008
timestamp 1682952543
transform 1 0 1724 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8040
timestamp 1682952543
transform 1 0 1756 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7978
timestamp 1682952543
transform 1 0 1796 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7979
timestamp 1682952543
transform 1 0 1828 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8005
timestamp 1682952543
transform 1 0 1812 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8006
timestamp 1682952543
transform 1 0 1844 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8007
timestamp 1682952543
transform 1 0 1860 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8079
timestamp 1682952543
transform 1 0 1772 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8080
timestamp 1682952543
transform 1 0 1788 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8081
timestamp 1682952543
transform 1 0 1812 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7890
timestamp 1682952543
transform 1 0 1764 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8135
timestamp 1682952543
transform 1 0 1740 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8025
timestamp 1682952543
transform 1 0 1884 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_8119
timestamp 1682952543
transform 1 0 1788 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7891
timestamp 1682952543
transform 1 0 1820 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7892
timestamp 1682952543
transform 1 0 1868 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8120
timestamp 1682952543
transform 1 0 1876 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8009
timestamp 1682952543
transform 1 0 1756 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8010
timestamp 1682952543
transform 1 0 1772 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8011
timestamp 1682952543
transform 1 0 1788 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8191
timestamp 1682952543
transform 1 0 1756 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8076
timestamp 1682952543
transform 1 0 1876 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_8192
timestamp 1682952543
transform 1 0 1876 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8082
timestamp 1682952543
transform 1 0 1900 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8136
timestamp 1682952543
transform 1 0 1892 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8026
timestamp 1682952543
transform 1 0 1924 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_7893
timestamp 1682952543
transform 1 0 1908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8077
timestamp 1682952543
transform 1 0 1892 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_8169
timestamp 1682952543
transform 1 0 1900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8121
timestamp 1682952543
transform 1 0 1916 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7894
timestamp 1682952543
transform 1 0 1940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8012
timestamp 1682952543
transform 1 0 1916 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8013
timestamp 1682952543
transform 1 0 1924 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8014
timestamp 1682952543
transform 1 0 1932 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8008
timestamp 1682952543
transform 1 0 1948 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7980
timestamp 1682952543
transform 1 0 1988 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8041
timestamp 1682952543
transform 1 0 1980 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8042
timestamp 1682952543
transform 1 0 2076 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7828
timestamp 1682952543
transform 1 0 1948 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_8083
timestamp 1682952543
transform 1 0 1956 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8084
timestamp 1682952543
transform 1 0 1972 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8085
timestamp 1682952543
transform 1 0 2060 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7895
timestamp 1682952543
transform 1 0 1964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7896
timestamp 1682952543
transform 1 0 2036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8015
timestamp 1682952543
transform 1 0 1972 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8016
timestamp 1682952543
transform 1 0 1988 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8137
timestamp 1682952543
transform 1 0 2028 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8170
timestamp 1682952543
transform 1 0 2012 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8193
timestamp 1682952543
transform 1 0 1988 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7981
timestamp 1682952543
transform 1 0 2100 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7982
timestamp 1682952543
transform 1 0 2116 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7983
timestamp 1682952543
transform 1 0 2140 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8009
timestamp 1682952543
transform 1 0 2092 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8086
timestamp 1682952543
transform 1 0 2084 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7829
timestamp 1682952543
transform 1 0 2092 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7897
timestamp 1682952543
transform 1 0 2084 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8043
timestamp 1682952543
transform 1 0 2124 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8087
timestamp 1682952543
transform 1 0 2132 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7898
timestamp 1682952543
transform 1 0 2108 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7899
timestamp 1682952543
transform 1 0 2124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7900
timestamp 1682952543
transform 1 0 2148 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8138
timestamp 1682952543
transform 1 0 2084 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8017
timestamp 1682952543
transform 1 0 2092 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8139
timestamp 1682952543
transform 1 0 2100 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7984
timestamp 1682952543
transform 1 0 2172 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_7901
timestamp 1682952543
transform 1 0 2164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8018
timestamp 1682952543
transform 1 0 2116 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8019
timestamp 1682952543
transform 1 0 2124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8020
timestamp 1682952543
transform 1 0 2140 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8021
timestamp 1682952543
transform 1 0 2156 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8171
timestamp 1682952543
transform 1 0 2116 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8172
timestamp 1682952543
transform 1 0 2148 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8194
timestamp 1682952543
transform 1 0 2116 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8195
timestamp 1682952543
transform 1 0 2148 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8196
timestamp 1682952543
transform 1 0 2172 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8022
timestamp 1682952543
transform 1 0 2188 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7985
timestamp 1682952543
transform 1 0 2228 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7986
timestamp 1682952543
transform 1 0 2284 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7987
timestamp 1682952543
transform 1 0 2316 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8010
timestamp 1682952543
transform 1 0 2244 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8011
timestamp 1682952543
transform 1 0 2276 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8088
timestamp 1682952543
transform 1 0 2228 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7902
timestamp 1682952543
transform 1 0 2228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8023
timestamp 1682952543
transform 1 0 2204 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8044
timestamp 1682952543
transform 1 0 2316 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8045
timestamp 1682952543
transform 1 0 2332 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8089
timestamp 1682952543
transform 1 0 2308 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8012
timestamp 1682952543
transform 1 0 2364 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8090
timestamp 1682952543
transform 1 0 2340 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7903
timestamp 1682952543
transform 1 0 2300 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7904
timestamp 1682952543
transform 1 0 2316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7905
timestamp 1682952543
transform 1 0 2332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7830
timestamp 1682952543
transform 1 0 2372 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7906
timestamp 1682952543
transform 1 0 2356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7907
timestamp 1682952543
transform 1 0 2372 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8024
timestamp 1682952543
transform 1 0 2308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8025
timestamp 1682952543
transform 1 0 2324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8026
timestamp 1682952543
transform 1 0 2340 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8027
timestamp 1682952543
transform 1 0 2348 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8173
timestamp 1682952543
transform 1 0 2284 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8174
timestamp 1682952543
transform 1 0 2324 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8091
timestamp 1682952543
transform 1 0 2396 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8028
timestamp 1682952543
transform 1 0 2372 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8140
timestamp 1682952543
transform 1 0 2380 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8029
timestamp 1682952543
transform 1 0 2388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8030
timestamp 1682952543
transform 1 0 2396 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8046
timestamp 1682952543
transform 1 0 2412 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8092
timestamp 1682952543
transform 1 0 2428 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8013
timestamp 1682952543
transform 1 0 2452 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_7908
timestamp 1682952543
transform 1 0 2404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7909
timestamp 1682952543
transform 1 0 2412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7910
timestamp 1682952543
transform 1 0 2428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7911
timestamp 1682952543
transform 1 0 2444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8031
timestamp 1682952543
transform 1 0 2412 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8197
timestamp 1682952543
transform 1 0 2412 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8078
timestamp 1682952543
transform 1 0 2468 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_8014
timestamp 1682952543
transform 1 0 2500 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8047
timestamp 1682952543
transform 1 0 2556 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8048
timestamp 1682952543
transform 1 0 2604 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7912
timestamp 1682952543
transform 1 0 2516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7913
timestamp 1682952543
transform 1 0 2564 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7914
timestamp 1682952543
transform 1 0 2572 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7915
timestamp 1682952543
transform 1 0 2588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7916
timestamp 1682952543
transform 1 0 2604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7917
timestamp 1682952543
transform 1 0 2628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8032
timestamp 1682952543
transform 1 0 2484 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8141
timestamp 1682952543
transform 1 0 2508 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8033
timestamp 1682952543
transform 1 0 2572 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8198
timestamp 1682952543
transform 1 0 2524 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8034
timestamp 1682952543
transform 1 0 2604 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8035
timestamp 1682952543
transform 1 0 2620 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8036
timestamp 1682952543
transform 1 0 2636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8037
timestamp 1682952543
transform 1 0 2644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8199
timestamp 1682952543
transform 1 0 2604 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_7918
timestamp 1682952543
transform 1 0 2660 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8142
timestamp 1682952543
transform 1 0 2668 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_7831
timestamp 1682952543
transform 1 0 2692 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7919
timestamp 1682952543
transform 1 0 2692 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8200
timestamp 1682952543
transform 1 0 2684 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8015
timestamp 1682952543
transform 1 0 2724 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8027
timestamp 1682952543
transform 1 0 2708 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_7821
timestamp 1682952543
transform 1 0 2708 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_8093
timestamp 1682952543
transform 1 0 2716 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7822
timestamp 1682952543
transform 1 0 2740 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_7832
timestamp 1682952543
transform 1 0 2724 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7833
timestamp 1682952543
transform 1 0 2732 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7920
timestamp 1682952543
transform 1 0 2716 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8122
timestamp 1682952543
transform 1 0 2740 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_8143
timestamp 1682952543
transform 1 0 2732 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8038
timestamp 1682952543
transform 1 0 2748 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8201
timestamp 1682952543
transform 1 0 2708 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8016
timestamp 1682952543
transform 1 0 2764 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_7834
timestamp 1682952543
transform 1 0 2764 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_8144
timestamp 1682952543
transform 1 0 2764 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8028
timestamp 1682952543
transform 1 0 2828 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_7921
timestamp 1682952543
transform 1 0 2804 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7922
timestamp 1682952543
transform 1 0 2860 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8039
timestamp 1682952543
transform 1 0 2780 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8145
timestamp 1682952543
transform 1 0 2804 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8029
timestamp 1682952543
transform 1 0 2884 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_8094
timestamp 1682952543
transform 1 0 2892 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7923
timestamp 1682952543
transform 1 0 2892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8040
timestamp 1682952543
transform 1 0 2876 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8041
timestamp 1682952543
transform 1 0 2884 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8202
timestamp 1682952543
transform 1 0 2884 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_7924
timestamp 1682952543
transform 1 0 2916 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7988
timestamp 1682952543
transform 1 0 2924 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8146
timestamp 1682952543
transform 1 0 2916 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_7925
timestamp 1682952543
transform 1 0 2948 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7926
timestamp 1682952543
transform 1 0 2964 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7989
timestamp 1682952543
transform 1 0 2988 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8030
timestamp 1682952543
transform 1 0 2988 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_8123
timestamp 1682952543
transform 1 0 2980 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8042
timestamp 1682952543
transform 1 0 2932 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8043
timestamp 1682952543
transform 1 0 2940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8044
timestamp 1682952543
transform 1 0 2956 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8147
timestamp 1682952543
transform 1 0 2972 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8017
timestamp 1682952543
transform 1 0 3012 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8049
timestamp 1682952543
transform 1 0 2996 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8095
timestamp 1682952543
transform 1 0 3004 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7927
timestamp 1682952543
transform 1 0 2996 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7928
timestamp 1682952543
transform 1 0 3004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7929
timestamp 1682952543
transform 1 0 3020 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8045
timestamp 1682952543
transform 1 0 2988 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8046
timestamp 1682952543
transform 1 0 2996 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8047
timestamp 1682952543
transform 1 0 3012 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8148
timestamp 1682952543
transform 1 0 3020 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_7930
timestamp 1682952543
transform 1 0 3036 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8048
timestamp 1682952543
transform 1 0 3028 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8018
timestamp 1682952543
transform 1 0 3044 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8019
timestamp 1682952543
transform 1 0 3156 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8031
timestamp 1682952543
transform 1 0 3164 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7990
timestamp 1682952543
transform 1 0 3220 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8050
timestamp 1682952543
transform 1 0 3204 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8051
timestamp 1682952543
transform 1 0 3236 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8096
timestamp 1682952543
transform 1 0 3156 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8097
timestamp 1682952543
transform 1 0 3180 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_8098
timestamp 1682952543
transform 1 0 3196 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7931
timestamp 1682952543
transform 1 0 3092 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7932
timestamp 1682952543
transform 1 0 3156 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7933
timestamp 1682952543
transform 1 0 3180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7934
timestamp 1682952543
transform 1 0 3196 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8149
timestamp 1682952543
transform 1 0 3092 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8150
timestamp 1682952543
transform 1 0 3108 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8049
timestamp 1682952543
transform 1 0 3140 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8050
timestamp 1682952543
transform 1 0 3156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8051
timestamp 1682952543
transform 1 0 3172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8052
timestamp 1682952543
transform 1 0 3188 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8099
timestamp 1682952543
transform 1 0 3228 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7991
timestamp 1682952543
transform 1 0 3332 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8020
timestamp 1682952543
transform 1 0 3276 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8032
timestamp 1682952543
transform 1 0 3332 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_8052
timestamp 1682952543
transform 1 0 3268 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8053
timestamp 1682952543
transform 1 0 3292 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8100
timestamp 1682952543
transform 1 0 3284 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7935
timestamp 1682952543
transform 1 0 3204 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7936
timestamp 1682952543
transform 1 0 3220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7937
timestamp 1682952543
transform 1 0 3236 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8124
timestamp 1682952543
transform 1 0 3244 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7992
timestamp 1682952543
transform 1 0 3404 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8054
timestamp 1682952543
transform 1 0 3380 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7938
timestamp 1682952543
transform 1 0 3252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7939
timestamp 1682952543
transform 1 0 3284 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7940
timestamp 1682952543
transform 1 0 3348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7941
timestamp 1682952543
transform 1 0 3380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8053
timestamp 1682952543
transform 1 0 3204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8054
timestamp 1682952543
transform 1 0 3212 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8055
timestamp 1682952543
transform 1 0 3228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8056
timestamp 1682952543
transform 1 0 3244 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8057
timestamp 1682952543
transform 1 0 3332 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8175
timestamp 1682952543
transform 1 0 3236 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8203
timestamp 1682952543
transform 1 0 3196 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8204
timestamp 1682952543
transform 1 0 3212 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8058
timestamp 1682952543
transform 1 0 3428 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8176
timestamp 1682952543
transform 1 0 3428 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8205
timestamp 1682952543
transform 1 0 3332 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8206
timestamp 1682952543
transform 1 0 3348 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8125
timestamp 1682952543
transform 1 0 3452 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7942
timestamp 1682952543
transform 1 0 3476 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7943
timestamp 1682952543
transform 1 0 3532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7944
timestamp 1682952543
transform 1 0 3596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8059
timestamp 1682952543
transform 1 0 3452 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8177
timestamp 1682952543
transform 1 0 3500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8178
timestamp 1682952543
transform 1 0 3524 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8207
timestamp 1682952543
transform 1 0 3484 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8060
timestamp 1682952543
transform 1 0 3548 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8179
timestamp 1682952543
transform 1 0 3596 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_7945
timestamp 1682952543
transform 1 0 3652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7946
timestamp 1682952543
transform 1 0 3676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7947
timestamp 1682952543
transform 1 0 3692 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8061
timestamp 1682952543
transform 1 0 3668 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8062
timestamp 1682952543
transform 1 0 3684 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8063
timestamp 1682952543
transform 1 0 3700 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8180
timestamp 1682952543
transform 1 0 3684 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8208
timestamp 1682952543
transform 1 0 3684 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8209
timestamp 1682952543
transform 1 0 3708 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8055
timestamp 1682952543
transform 1 0 3732 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8151
timestamp 1682952543
transform 1 0 3740 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7993
timestamp 1682952543
transform 1 0 3764 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_7823
timestamp 1682952543
transform 1 0 3764 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_8056
timestamp 1682952543
transform 1 0 3780 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_7835
timestamp 1682952543
transform 1 0 3756 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_8101
timestamp 1682952543
transform 1 0 3772 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7836
timestamp 1682952543
transform 1 0 3780 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_7948
timestamp 1682952543
transform 1 0 3772 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8057
timestamp 1682952543
transform 1 0 3804 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7994
timestamp 1682952543
transform 1 0 3836 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_8033
timestamp 1682952543
transform 1 0 3844 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_8102
timestamp 1682952543
transform 1 0 3828 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7949
timestamp 1682952543
transform 1 0 3812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7950
timestamp 1682952543
transform 1 0 3828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7951
timestamp 1682952543
transform 1 0 3844 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7952
timestamp 1682952543
transform 1 0 3852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8064
timestamp 1682952543
transform 1 0 3820 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8152
timestamp 1682952543
transform 1 0 3852 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8065
timestamp 1682952543
transform 1 0 3860 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8181
timestamp 1682952543
transform 1 0 3860 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8034
timestamp 1682952543
transform 1 0 3884 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_8058
timestamp 1682952543
transform 1 0 3916 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_8126
timestamp 1682952543
transform 1 0 3892 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_7953
timestamp 1682952543
transform 1 0 3916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7954
timestamp 1682952543
transform 1 0 3972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7955
timestamp 1682952543
transform 1 0 3980 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8066
timestamp 1682952543
transform 1 0 3876 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8067
timestamp 1682952543
transform 1 0 3892 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8153
timestamp 1682952543
transform 1 0 3916 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8154
timestamp 1682952543
transform 1 0 3964 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_8103
timestamp 1682952543
transform 1 0 4020 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7956
timestamp 1682952543
transform 1 0 4004 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7957
timestamp 1682952543
transform 1 0 4020 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_8021
timestamp 1682952543
transform 1 0 4044 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_8104
timestamp 1682952543
transform 1 0 4068 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_7958
timestamp 1682952543
transform 1 0 4068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7959
timestamp 1682952543
transform 1 0 4124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_7960
timestamp 1682952543
transform 1 0 4132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8068
timestamp 1682952543
transform 1 0 3988 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8069
timestamp 1682952543
transform 1 0 3996 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8070
timestamp 1682952543
transform 1 0 4012 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8071
timestamp 1682952543
transform 1 0 4028 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8072
timestamp 1682952543
transform 1 0 4044 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8210
timestamp 1682952543
transform 1 0 3884 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8182
timestamp 1682952543
transform 1 0 4020 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8211
timestamp 1682952543
transform 1 0 3996 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8073
timestamp 1682952543
transform 1 0 4148 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_8183
timestamp 1682952543
transform 1 0 4132 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_8212
timestamp 1682952543
transform 1 0 4044 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_8213
timestamp 1682952543
transform 1 0 4068 0 1 785
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_66
timestamp 1682952543
transform 1 0 48 0 1 770
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_491
timestamp 1682952543
transform 1 0 72 0 1 770
box -8 -3 104 105
use AOI22X1  AOI22X1_325
timestamp 1682952543
transform 1 0 168 0 1 770
box -8 -3 46 105
use FILL  FILL_3556
timestamp 1682952543
transform 1 0 208 0 1 770
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1682952543
transform 1 0 216 0 1 770
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1682952543
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1682952543
transform 1 0 232 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8214
timestamp 1682952543
transform 1 0 260 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_8215
timestamp 1682952543
transform 1 0 276 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_326
timestamp 1682952543
transform 1 0 240 0 1 770
box -8 -3 46 105
use FILL  FILL_3560
timestamp 1682952543
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1682952543
transform 1 0 288 0 1 770
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1682952543
transform 1 0 296 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8216
timestamp 1682952543
transform 1 0 324 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_352
timestamp 1682952543
transform 1 0 304 0 1 770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_494
timestamp 1682952543
transform 1 0 344 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_495
timestamp 1682952543
transform 1 0 440 0 1 770
box -8 -3 104 105
use INVX2  INVX2_566
timestamp 1682952543
transform -1 0 552 0 1 770
box -9 -3 26 105
use FILL  FILL_3564
timestamp 1682952543
transform 1 0 552 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_327
timestamp 1682952543
transform -1 0 600 0 1 770
box -8 -3 46 105
use FILL  FILL_3565
timestamp 1682952543
transform 1 0 600 0 1 770
box -8 -3 16 105
use FILL  FILL_3566
timestamp 1682952543
transform 1 0 608 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_496
timestamp 1682952543
transform 1 0 616 0 1 770
box -8 -3 104 105
use FILL  FILL_3567
timestamp 1682952543
transform 1 0 712 0 1 770
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1682952543
transform 1 0 720 0 1 770
box -8 -3 16 105
use INVX2  INVX2_567
timestamp 1682952543
transform -1 0 744 0 1 770
box -9 -3 26 105
use FILL  FILL_3569
timestamp 1682952543
transform 1 0 744 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_328
timestamp 1682952543
transform 1 0 752 0 1 770
box -8 -3 46 105
use FILL  FILL_3570
timestamp 1682952543
transform 1 0 792 0 1 770
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1682952543
transform 1 0 800 0 1 770
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1682952543
transform 1 0 808 0 1 770
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1682952543
transform 1 0 816 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_135
timestamp 1682952543
transform 1 0 824 0 1 770
box -8 -3 34 105
use M3_M2  M3_M2_8217
timestamp 1682952543
transform 1 0 868 0 1 775
box -3 -3 3 3
use FILL  FILL_3574
timestamp 1682952543
transform 1 0 856 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_95
timestamp 1682952543
transform 1 0 864 0 1 770
box -8 -3 32 105
use FILL  FILL_3575
timestamp 1682952543
transform 1 0 888 0 1 770
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1682952543
transform 1 0 896 0 1 770
box -8 -3 16 105
use FILL  FILL_3577
timestamp 1682952543
transform 1 0 904 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_96
timestamp 1682952543
transform 1 0 912 0 1 770
box -8 -3 32 105
use FILL  FILL_3578
timestamp 1682952543
transform 1 0 936 0 1 770
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1682952543
transform 1 0 944 0 1 770
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1682952543
transform 1 0 952 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_138
timestamp 1682952543
transform 1 0 960 0 1 770
box -8 -3 34 105
use FILL  FILL_3594
timestamp 1682952543
transform 1 0 992 0 1 770
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1682952543
transform 1 0 1000 0 1 770
box -8 -3 16 105
use FILL  FILL_3596
timestamp 1682952543
transform 1 0 1008 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_139
timestamp 1682952543
transform -1 0 1048 0 1 770
box -8 -3 34 105
use FILL  FILL_3597
timestamp 1682952543
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1682952543
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_3599
timestamp 1682952543
transform 1 0 1064 0 1 770
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1682952543
transform 1 0 1072 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8218
timestamp 1682952543
transform 1 0 1100 0 1 775
box -3 -3 3 3
use INVX2  INVX2_570
timestamp 1682952543
transform -1 0 1096 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_8219
timestamp 1682952543
transform 1 0 1124 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_8220
timestamp 1682952543
transform 1 0 1140 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_8221
timestamp 1682952543
transform 1 0 1188 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_499
timestamp 1682952543
transform -1 0 1192 0 1 770
box -8 -3 104 105
use OAI22X1  OAI22X1_355
timestamp 1682952543
transform -1 0 1232 0 1 770
box -8 -3 46 105
use FILL  FILL_3601
timestamp 1682952543
transform 1 0 1232 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_356
timestamp 1682952543
transform -1 0 1280 0 1 770
box -8 -3 46 105
use FILL  FILL_3602
timestamp 1682952543
transform 1 0 1280 0 1 770
box -8 -3 16 105
use INVX2  INVX2_571
timestamp 1682952543
transform -1 0 1304 0 1 770
box -9 -3 26 105
use FILL  FILL_3603
timestamp 1682952543
transform 1 0 1304 0 1 770
box -8 -3 16 105
use FILL  FILL_3604
timestamp 1682952543
transform 1 0 1312 0 1 770
box -8 -3 16 105
use INVX2  INVX2_572
timestamp 1682952543
transform -1 0 1336 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_8222
timestamp 1682952543
transform 1 0 1348 0 1 775
box -3 -3 3 3
use FILL  FILL_3605
timestamp 1682952543
transform 1 0 1336 0 1 770
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1682952543
transform 1 0 1344 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_357
timestamp 1682952543
transform -1 0 1392 0 1 770
box -8 -3 46 105
use FILL  FILL_3607
timestamp 1682952543
transform 1 0 1392 0 1 770
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1682952543
transform 1 0 1400 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8223
timestamp 1682952543
transform 1 0 1452 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_500
timestamp 1682952543
transform 1 0 1408 0 1 770
box -8 -3 104 105
use INVX2  INVX2_573
timestamp 1682952543
transform -1 0 1520 0 1 770
box -9 -3 26 105
use FILL  FILL_3609
timestamp 1682952543
transform 1 0 1520 0 1 770
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1682952543
transform 1 0 1528 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8224
timestamp 1682952543
transform 1 0 1548 0 1 775
box -3 -3 3 3
use FILL  FILL_3611
timestamp 1682952543
transform 1 0 1536 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_334
timestamp 1682952543
transform -1 0 1584 0 1 770
box -8 -3 46 105
use FILL  FILL_3612
timestamp 1682952543
transform 1 0 1584 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8225
timestamp 1682952543
transform 1 0 1652 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_501
timestamp 1682952543
transform 1 0 1592 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_8226
timestamp 1682952543
transform 1 0 1700 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_335
timestamp 1682952543
transform 1 0 1688 0 1 770
box -8 -3 46 105
use FILL  FILL_3613
timestamp 1682952543
transform 1 0 1728 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_358
timestamp 1682952543
transform 1 0 1736 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_8227
timestamp 1682952543
transform 1 0 1828 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_8228
timestamp 1682952543
transform 1 0 1876 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_502
timestamp 1682952543
transform 1 0 1776 0 1 770
box -8 -3 104 105
use NOR2X1  NOR2X1_97
timestamp 1682952543
transform 1 0 1872 0 1 770
box -8 -3 32 105
use FILL  FILL_3614
timestamp 1682952543
transform 1 0 1896 0 1 770
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1682952543
transform 1 0 1904 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_98
timestamp 1682952543
transform 1 0 1912 0 1 770
box -8 -3 32 105
use FILL  FILL_3616
timestamp 1682952543
transform 1 0 1936 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8229
timestamp 1682952543
transform 1 0 1964 0 1 775
box -3 -3 3 3
use OAI21X1  OAI21X1_140
timestamp 1682952543
transform -1 0 1976 0 1 770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_503
timestamp 1682952543
transform 1 0 1976 0 1 770
box -8 -3 104 105
use INVX2  INVX2_574
timestamp 1682952543
transform 1 0 2072 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_8230
timestamp 1682952543
transform 1 0 2108 0 1 775
box -3 -3 3 3
use OAI21X1  OAI21X1_141
timestamp 1682952543
transform -1 0 2120 0 1 770
box -8 -3 34 105
use OAI22X1  OAI22X1_359
timestamp 1682952543
transform 1 0 2120 0 1 770
box -8 -3 46 105
use FILL  FILL_3617
timestamp 1682952543
transform 1 0 2160 0 1 770
box -8 -3 16 105
use INVX2  INVX2_575
timestamp 1682952543
transform -1 0 2184 0 1 770
box -9 -3 26 105
use FILL  FILL_3618
timestamp 1682952543
transform 1 0 2184 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_504
timestamp 1682952543
transform 1 0 2192 0 1 770
box -8 -3 104 105
use INVX2  INVX2_576
timestamp 1682952543
transform 1 0 2288 0 1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_360
timestamp 1682952543
transform 1 0 2304 0 1 770
box -8 -3 46 105
use OAI21X1  OAI21X1_142
timestamp 1682952543
transform 1 0 2344 0 1 770
box -8 -3 34 105
use INVX2  INVX2_577
timestamp 1682952543
transform -1 0 2392 0 1 770
box -9 -3 26 105
use INVX2  INVX2_578
timestamp 1682952543
transform 1 0 2392 0 1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_336
timestamp 1682952543
transform 1 0 2408 0 1 770
box -8 -3 46 105
use FILL  FILL_3619
timestamp 1682952543
transform 1 0 2448 0 1 770
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1682952543
transform 1 0 2456 0 1 770
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1682952543
transform 1 0 2464 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8231
timestamp 1682952543
transform 1 0 2548 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_8232
timestamp 1682952543
transform 1 0 2564 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_505
timestamp 1682952543
transform 1 0 2472 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_8233
timestamp 1682952543
transform 1 0 2612 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_337
timestamp 1682952543
transform -1 0 2608 0 1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_338
timestamp 1682952543
transform 1 0 2608 0 1 770
box -8 -3 46 105
use FILL  FILL_3622
timestamp 1682952543
transform 1 0 2648 0 1 770
box -8 -3 16 105
use INVX2  INVX2_579
timestamp 1682952543
transform 1 0 2656 0 1 770
box -9 -3 26 105
use FILL  FILL_3623
timestamp 1682952543
transform 1 0 2672 0 1 770
box -8 -3 16 105
use FILL  FILL_3624
timestamp 1682952543
transform 1 0 2680 0 1 770
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1682952543
transform 1 0 2688 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_66
timestamp 1682952543
transform -1 0 2728 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_67
timestamp 1682952543
transform -1 0 2760 0 1 770
box -8 -3 40 105
use FILL  FILL_3626
timestamp 1682952543
transform 1 0 2760 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8234
timestamp 1682952543
transform 1 0 2788 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_8235
timestamp 1682952543
transform 1 0 2812 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_506
timestamp 1682952543
transform 1 0 2768 0 1 770
box -8 -3 104 105
use FILL  FILL_3627
timestamp 1682952543
transform 1 0 2864 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8236
timestamp 1682952543
transform 1 0 2892 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_339
timestamp 1682952543
transform 1 0 2872 0 1 770
box -8 -3 46 105
use FILL  FILL_3628
timestamp 1682952543
transform 1 0 2912 0 1 770
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1682952543
transform 1 0 2920 0 1 770
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1682952543
transform 1 0 2928 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8237
timestamp 1682952543
transform 1 0 2956 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_361
timestamp 1682952543
transform -1 0 2976 0 1 770
box -8 -3 46 105
use FILL  FILL_3631
timestamp 1682952543
transform 1 0 2976 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8238
timestamp 1682952543
transform 1 0 2996 0 1 775
box -3 -3 3 3
use FILL  FILL_3632
timestamp 1682952543
transform 1 0 2984 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_362
timestamp 1682952543
transform 1 0 2992 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_8239
timestamp 1682952543
transform 1 0 3044 0 1 775
box -3 -3 3 3
use FILL  FILL_3633
timestamp 1682952543
transform 1 0 3032 0 1 770
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1682952543
transform 1 0 3040 0 1 770
box -8 -3 16 105
use FILL  FILL_3635
timestamp 1682952543
transform 1 0 3048 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8240
timestamp 1682952543
transform 1 0 3140 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_507
timestamp 1682952543
transform -1 0 3152 0 1 770
box -8 -3 104 105
use OAI22X1  OAI22X1_363
timestamp 1682952543
transform 1 0 3152 0 1 770
box -8 -3 46 105
use INVX2  INVX2_580
timestamp 1682952543
transform -1 0 3208 0 1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_364
timestamp 1682952543
transform 1 0 3208 0 1 770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_508
timestamp 1682952543
transform -1 0 3344 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_509
timestamp 1682952543
transform -1 0 3440 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_8241
timestamp 1682952543
transform 1 0 3452 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_510
timestamp 1682952543
transform 1 0 3440 0 1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_511
timestamp 1682952543
transform 1 0 3536 0 1 770
box -8 -3 104 105
use FILL  FILL_3682
timestamp 1682952543
transform 1 0 3632 0 1 770
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1682952543
transform 1 0 3640 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8242
timestamp 1682952543
transform 1 0 3668 0 1 775
box -3 -3 3 3
use FILL  FILL_3684
timestamp 1682952543
transform 1 0 3648 0 1 770
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1682952543
transform 1 0 3656 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8243
timestamp 1682952543
transform 1 0 3700 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_372
timestamp 1682952543
transform -1 0 3704 0 1 770
box -8 -3 46 105
use FILL  FILL_3687
timestamp 1682952543
transform 1 0 3704 0 1 770
box -8 -3 16 105
use FILL  FILL_3690
timestamp 1682952543
transform 1 0 3712 0 1 770
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1682952543
transform 1 0 3720 0 1 770
box -8 -3 16 105
use FILL  FILL_3692
timestamp 1682952543
transform 1 0 3728 0 1 770
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1682952543
transform 1 0 3736 0 1 770
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1682952543
transform 1 0 3744 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_69
timestamp 1682952543
transform -1 0 3784 0 1 770
box -8 -3 40 105
use FILL  FILL_3695
timestamp 1682952543
transform 1 0 3784 0 1 770
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1682952543
transform 1 0 3792 0 1 770
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1682952543
transform 1 0 3800 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8244
timestamp 1682952543
transform 1 0 3820 0 1 775
box -3 -3 3 3
use AOI22X1  AOI22X1_346
timestamp 1682952543
transform 1 0 3808 0 1 770
box -8 -3 46 105
use FILL  FILL_3698
timestamp 1682952543
transform 1 0 3848 0 1 770
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1682952543
transform 1 0 3856 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_8245
timestamp 1682952543
transform 1 0 3900 0 1 775
box -3 -3 3 3
use INVX2  INVX2_594
timestamp 1682952543
transform -1 0 3880 0 1 770
box -9 -3 26 105
use M3_M2  M3_M2_8246
timestamp 1682952543
transform 1 0 3980 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_526
timestamp 1682952543
transform 1 0 3880 0 1 770
box -8 -3 104 105
use INVX2  INVX2_595
timestamp 1682952543
transform -1 0 3992 0 1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_374
timestamp 1682952543
transform 1 0 3992 0 1 770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_527
timestamp 1682952543
transform 1 0 4032 0 1 770
box -8 -3 104 105
use INVX2  INVX2_596
timestamp 1682952543
transform -1 0 4144 0 1 770
box -9 -3 26 105
use FILL  FILL_3700
timestamp 1682952543
transform 1 0 4144 0 1 770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_67
timestamp 1682952543
transform 1 0 4177 0 1 770
box -10 -3 10 3
use M2_M1  M2_M1_8082
timestamp 1682952543
transform 1 0 84 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8348
timestamp 1682952543
transform 1 0 148 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8302
timestamp 1682952543
transform 1 0 180 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8303
timestamp 1682952543
transform 1 0 212 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8304
timestamp 1682952543
transform 1 0 244 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8083
timestamp 1682952543
transform 1 0 180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8084
timestamp 1682952543
transform 1 0 268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8192
timestamp 1682952543
transform 1 0 124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8193
timestamp 1682952543
transform 1 0 164 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8383
timestamp 1682952543
transform 1 0 180 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8384
timestamp 1682952543
transform 1 0 204 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8349
timestamp 1682952543
transform 1 0 276 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8194
timestamp 1682952543
transform 1 0 228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8195
timestamp 1682952543
transform 1 0 260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8196
timestamp 1682952543
transform 1 0 268 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8422
timestamp 1682952543
transform 1 0 228 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8423
timestamp 1682952543
transform 1 0 268 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8247
timestamp 1682952543
transform 1 0 300 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8248
timestamp 1682952543
transform 1 0 356 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8305
timestamp 1682952543
transform 1 0 300 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8085
timestamp 1682952543
transform 1 0 300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8197
timestamp 1682952543
transform 1 0 348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8198
timestamp 1682952543
transform 1 0 380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8199
timestamp 1682952543
transform 1 0 388 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8200
timestamp 1682952543
transform 1 0 396 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8424
timestamp 1682952543
transform 1 0 348 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8425
timestamp 1682952543
transform 1 0 388 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8434
timestamp 1682952543
transform 1 0 380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8485
timestamp 1682952543
transform 1 0 396 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8086
timestamp 1682952543
transform 1 0 412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8087
timestamp 1682952543
transform 1 0 420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8088
timestamp 1682952543
transform 1 0 436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8201
timestamp 1682952543
transform 1 0 428 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8435
timestamp 1682952543
transform 1 0 420 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8466
timestamp 1682952543
transform 1 0 436 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8350
timestamp 1682952543
transform 1 0 460 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8306
timestamp 1682952543
transform 1 0 500 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8089
timestamp 1682952543
transform 1 0 476 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8351
timestamp 1682952543
transform 1 0 484 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8249
timestamp 1682952543
transform 1 0 580 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8270
timestamp 1682952543
transform 1 0 572 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8307
timestamp 1682952543
transform 1 0 556 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8090
timestamp 1682952543
transform 1 0 492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8091
timestamp 1682952543
transform 1 0 500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8092
timestamp 1682952543
transform 1 0 508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8093
timestamp 1682952543
transform 1 0 524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8094
timestamp 1682952543
transform 1 0 540 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8095
timestamp 1682952543
transform 1 0 548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8202
timestamp 1682952543
transform 1 0 468 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8385
timestamp 1682952543
transform 1 0 476 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8203
timestamp 1682952543
transform 1 0 484 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8386
timestamp 1682952543
transform 1 0 492 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8204
timestamp 1682952543
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8205
timestamp 1682952543
transform 1 0 532 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8387
timestamp 1682952543
transform 1 0 540 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8426
timestamp 1682952543
transform 1 0 516 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8436
timestamp 1682952543
transform 1 0 508 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8308
timestamp 1682952543
transform 1 0 596 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8309
timestamp 1682952543
transform 1 0 620 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8096
timestamp 1682952543
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8097
timestamp 1682952543
transform 1 0 596 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8098
timestamp 1682952543
transform 1 0 604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8206
timestamp 1682952543
transform 1 0 564 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8388
timestamp 1682952543
transform 1 0 572 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8352
timestamp 1682952543
transform 1 0 612 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8099
timestamp 1682952543
transform 1 0 620 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8207
timestamp 1682952543
transform 1 0 580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8208
timestamp 1682952543
transform 1 0 588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8209
timestamp 1682952543
transform 1 0 612 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8427
timestamp 1682952543
transform 1 0 580 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8437
timestamp 1682952543
transform 1 0 564 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8467
timestamp 1682952543
transform 1 0 564 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8468
timestamp 1682952543
transform 1 0 604 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8210
timestamp 1682952543
transform 1 0 636 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8486
timestamp 1682952543
transform 1 0 636 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8100
timestamp 1682952543
transform 1 0 660 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8353
timestamp 1682952543
transform 1 0 708 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8354
timestamp 1682952543
transform 1 0 748 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8211
timestamp 1682952543
transform 1 0 708 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8389
timestamp 1682952543
transform 1 0 732 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8212
timestamp 1682952543
transform 1 0 740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8213
timestamp 1682952543
transform 1 0 748 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8469
timestamp 1682952543
transform 1 0 676 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8470
timestamp 1682952543
transform 1 0 700 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8487
timestamp 1682952543
transform 1 0 732 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8355
timestamp 1682952543
transform 1 0 772 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8214
timestamp 1682952543
transform 1 0 772 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8101
timestamp 1682952543
transform 1 0 788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8102
timestamp 1682952543
transform 1 0 796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8103
timestamp 1682952543
transform 1 0 812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8104
timestamp 1682952543
transform 1 0 820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8105
timestamp 1682952543
transform 1 0 828 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8390
timestamp 1682952543
transform 1 0 796 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8215
timestamp 1682952543
transform 1 0 804 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8391
timestamp 1682952543
transform 1 0 828 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8438
timestamp 1682952543
transform 1 0 820 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8471
timestamp 1682952543
transform 1 0 812 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8271
timestamp 1682952543
transform 1 0 852 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8310
timestamp 1682952543
transform 1 0 852 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8216
timestamp 1682952543
transform 1 0 844 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8272
timestamp 1682952543
transform 1 0 868 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8311
timestamp 1682952543
transform 1 0 884 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8106
timestamp 1682952543
transform 1 0 876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8107
timestamp 1682952543
transform 1 0 884 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8356
timestamp 1682952543
transform 1 0 908 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8108
timestamp 1682952543
transform 1 0 916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8217
timestamp 1682952543
transform 1 0 876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8218
timestamp 1682952543
transform 1 0 892 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8219
timestamp 1682952543
transform 1 0 908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8308
timestamp 1682952543
transform 1 0 868 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8439
timestamp 1682952543
transform 1 0 900 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8472
timestamp 1682952543
transform 1 0 884 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8357
timestamp 1682952543
transform 1 0 932 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8109
timestamp 1682952543
transform 1 0 948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8220
timestamp 1682952543
transform 1 0 932 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8473
timestamp 1682952543
transform 1 0 940 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8110
timestamp 1682952543
transform 1 0 956 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8358
timestamp 1682952543
transform 1 0 972 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8309
timestamp 1682952543
transform 1 0 972 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8273
timestamp 1682952543
transform 1 0 1012 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8312
timestamp 1682952543
transform 1 0 996 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8274
timestamp 1682952543
transform 1 0 1036 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8313
timestamp 1682952543
transform 1 0 1028 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8111
timestamp 1682952543
transform 1 0 1012 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8359
timestamp 1682952543
transform 1 0 1020 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8112
timestamp 1682952543
transform 1 0 1036 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8392
timestamp 1682952543
transform 1 0 980 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8221
timestamp 1682952543
transform 1 0 996 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8393
timestamp 1682952543
transform 1 0 1004 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8222
timestamp 1682952543
transform 1 0 1012 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8223
timestamp 1682952543
transform 1 0 1028 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8224
timestamp 1682952543
transform 1 0 1036 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8310
timestamp 1682952543
transform 1 0 980 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8440
timestamp 1682952543
transform 1 0 972 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8474
timestamp 1682952543
transform 1 0 972 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8311
timestamp 1682952543
transform 1 0 1012 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8475
timestamp 1682952543
transform 1 0 996 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8394
timestamp 1682952543
transform 1 0 1044 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8312
timestamp 1682952543
transform 1 0 1044 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8441
timestamp 1682952543
transform 1 0 1036 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8314
timestamp 1682952543
transform 1 0 1076 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8113
timestamp 1682952543
transform 1 0 1076 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8225
timestamp 1682952543
transform 1 0 1068 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8476
timestamp 1682952543
transform 1 0 1060 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8360
timestamp 1682952543
transform 1 0 1084 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8114
timestamp 1682952543
transform 1 0 1092 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8226
timestamp 1682952543
transform 1 0 1084 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8315
timestamp 1682952543
transform 1 0 1132 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8080
timestamp 1682952543
transform 1 0 1180 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_8115
timestamp 1682952543
transform 1 0 1124 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8116
timestamp 1682952543
transform 1 0 1140 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8361
timestamp 1682952543
transform 1 0 1148 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8117
timestamp 1682952543
transform 1 0 1156 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8362
timestamp 1682952543
transform 1 0 1180 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8316
timestamp 1682952543
transform 1 0 1204 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8118
timestamp 1682952543
transform 1 0 1188 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8119
timestamp 1682952543
transform 1 0 1204 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8227
timestamp 1682952543
transform 1 0 1132 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8395
timestamp 1682952543
transform 1 0 1140 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8228
timestamp 1682952543
transform 1 0 1148 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8363
timestamp 1682952543
transform 1 0 1212 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8229
timestamp 1682952543
transform 1 0 1180 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8396
timestamp 1682952543
transform 1 0 1188 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8230
timestamp 1682952543
transform 1 0 1196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8231
timestamp 1682952543
transform 1 0 1212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8120
timestamp 1682952543
transform 1 0 1228 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8317
timestamp 1682952543
transform 1 0 1244 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8121
timestamp 1682952543
transform 1 0 1244 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8275
timestamp 1682952543
transform 1 0 1348 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8318
timestamp 1682952543
transform 1 0 1412 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8122
timestamp 1682952543
transform 1 0 1412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8232
timestamp 1682952543
transform 1 0 1268 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8233
timestamp 1682952543
transform 1 0 1324 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8234
timestamp 1682952543
transform 1 0 1332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8235
timestamp 1682952543
transform 1 0 1372 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8319
timestamp 1682952543
transform 1 0 1460 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8320
timestamp 1682952543
transform 1 0 1516 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8123
timestamp 1682952543
transform 1 0 1436 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8364
timestamp 1682952543
transform 1 0 1484 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8236
timestamp 1682952543
transform 1 0 1484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8237
timestamp 1682952543
transform 1 0 1516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8238
timestamp 1682952543
transform 1 0 1524 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8442
timestamp 1682952543
transform 1 0 1484 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8488
timestamp 1682952543
transform 1 0 1508 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8443
timestamp 1682952543
transform 1 0 1524 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8489
timestamp 1682952543
transform 1 0 1524 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8397
timestamp 1682952543
transform 1 0 1540 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8321
timestamp 1682952543
transform 1 0 1580 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8124
timestamp 1682952543
transform 1 0 1556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8125
timestamp 1682952543
transform 1 0 1564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8126
timestamp 1682952543
transform 1 0 1580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8127
timestamp 1682952543
transform 1 0 1588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8239
timestamp 1682952543
transform 1 0 1548 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8398
timestamp 1682952543
transform 1 0 1556 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8240
timestamp 1682952543
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8399
timestamp 1682952543
transform 1 0 1580 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8241
timestamp 1682952543
transform 1 0 1588 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8444
timestamp 1682952543
transform 1 0 1564 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8400
timestamp 1682952543
transform 1 0 1596 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8128
timestamp 1682952543
transform 1 0 1612 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8445
timestamp 1682952543
transform 1 0 1612 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8446
timestamp 1682952543
transform 1 0 1628 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8276
timestamp 1682952543
transform 1 0 1652 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8129
timestamp 1682952543
transform 1 0 1644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8130
timestamp 1682952543
transform 1 0 1652 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8131
timestamp 1682952543
transform 1 0 1668 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8132
timestamp 1682952543
transform 1 0 1676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8242
timestamp 1682952543
transform 1 0 1636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8243
timestamp 1682952543
transform 1 0 1644 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8244
timestamp 1682952543
transform 1 0 1660 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8401
timestamp 1682952543
transform 1 0 1668 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8245
timestamp 1682952543
transform 1 0 1676 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8447
timestamp 1682952543
transform 1 0 1668 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8490
timestamp 1682952543
transform 1 0 1644 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8477
timestamp 1682952543
transform 1 0 1676 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8277
timestamp 1682952543
transform 1 0 1692 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8322
timestamp 1682952543
transform 1 0 1724 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8133
timestamp 1682952543
transform 1 0 1796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8246
timestamp 1682952543
transform 1 0 1708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8247
timestamp 1682952543
transform 1 0 1716 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8448
timestamp 1682952543
transform 1 0 1708 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8402
timestamp 1682952543
transform 1 0 1724 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8248
timestamp 1682952543
transform 1 0 1748 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8449
timestamp 1682952543
transform 1 0 1748 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8478
timestamp 1682952543
transform 1 0 1732 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8134
timestamp 1682952543
transform 1 0 1828 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8135
timestamp 1682952543
transform 1 0 1836 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8249
timestamp 1682952543
transform 1 0 1820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8250
timestamp 1682952543
transform 1 0 1828 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8403
timestamp 1682952543
transform 1 0 1836 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8323
timestamp 1682952543
transform 1 0 1868 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8324
timestamp 1682952543
transform 1 0 1892 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8136
timestamp 1682952543
transform 1 0 1868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8137
timestamp 1682952543
transform 1 0 1876 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8138
timestamp 1682952543
transform 1 0 1892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8251
timestamp 1682952543
transform 1 0 1844 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8252
timestamp 1682952543
transform 1 0 1860 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8491
timestamp 1682952543
transform 1 0 1828 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8404
timestamp 1682952543
transform 1 0 1876 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8139
timestamp 1682952543
transform 1 0 1916 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8253
timestamp 1682952543
transform 1 0 1900 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8479
timestamp 1682952543
transform 1 0 1884 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8325
timestamp 1682952543
transform 1 0 1964 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8254
timestamp 1682952543
transform 1 0 1956 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8313
timestamp 1682952543
transform 1 0 1940 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8492
timestamp 1682952543
transform 1 0 1948 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8140
timestamp 1682952543
transform 1 0 1988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8141
timestamp 1682952543
transform 1 0 1996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8142
timestamp 1682952543
transform 1 0 2012 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8405
timestamp 1682952543
transform 1 0 1988 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8314
timestamp 1682952543
transform 1 0 1988 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8255
timestamp 1682952543
transform 1 0 2004 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8256
timestamp 1682952543
transform 1 0 2020 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8406
timestamp 1682952543
transform 1 0 2028 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8257
timestamp 1682952543
transform 1 0 2036 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8450
timestamp 1682952543
transform 1 0 2004 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8493
timestamp 1682952543
transform 1 0 2028 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8278
timestamp 1682952543
transform 1 0 2044 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8143
timestamp 1682952543
transform 1 0 2044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8315
timestamp 1682952543
transform 1 0 2060 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8279
timestamp 1682952543
transform 1 0 2068 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8144
timestamp 1682952543
transform 1 0 2084 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8451
timestamp 1682952543
transform 1 0 2076 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8280
timestamp 1682952543
transform 1 0 2156 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8145
timestamp 1682952543
transform 1 0 2116 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8258
timestamp 1682952543
transform 1 0 2140 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8259
timestamp 1682952543
transform 1 0 2196 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8407
timestamp 1682952543
transform 1 0 2204 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8281
timestamp 1682952543
transform 1 0 2292 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8365
timestamp 1682952543
transform 1 0 2268 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8146
timestamp 1682952543
transform 1 0 2292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8260
timestamp 1682952543
transform 1 0 2212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8261
timestamp 1682952543
transform 1 0 2268 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8480
timestamp 1682952543
transform 1 0 2196 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8408
timestamp 1682952543
transform 1 0 2292 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8452
timestamp 1682952543
transform 1 0 2212 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8453
timestamp 1682952543
transform 1 0 2252 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8481
timestamp 1682952543
transform 1 0 2260 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8147
timestamp 1682952543
transform 1 0 2316 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8262
timestamp 1682952543
transform 1 0 2308 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8366
timestamp 1682952543
transform 1 0 2324 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8148
timestamp 1682952543
transform 1 0 2332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8149
timestamp 1682952543
transform 1 0 2348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8263
timestamp 1682952543
transform 1 0 2340 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8282
timestamp 1682952543
transform 1 0 2380 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8150
timestamp 1682952543
transform 1 0 2380 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8151
timestamp 1682952543
transform 1 0 2468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8264
timestamp 1682952543
transform 1 0 2404 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8482
timestamp 1682952543
transform 1 0 2396 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8494
timestamp 1682952543
transform 1 0 2380 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8495
timestamp 1682952543
transform 1 0 2436 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8265
timestamp 1682952543
transform 1 0 2476 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8316
timestamp 1682952543
transform 1 0 2492 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8283
timestamp 1682952543
transform 1 0 2516 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8081
timestamp 1682952543
transform 1 0 2516 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_8250
timestamp 1682952543
transform 1 0 2540 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8152
timestamp 1682952543
transform 1 0 2516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8153
timestamp 1682952543
transform 1 0 2532 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8266
timestamp 1682952543
transform 1 0 2524 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8428
timestamp 1682952543
transform 1 0 2524 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8483
timestamp 1682952543
transform 1 0 2516 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8367
timestamp 1682952543
transform 1 0 2548 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8284
timestamp 1682952543
transform 1 0 2572 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8154
timestamp 1682952543
transform 1 0 2556 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8155
timestamp 1682952543
transform 1 0 2572 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8368
timestamp 1682952543
transform 1 0 2580 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8285
timestamp 1682952543
transform 1 0 2628 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8286
timestamp 1682952543
transform 1 0 2660 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8287
timestamp 1682952543
transform 1 0 2676 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8288
timestamp 1682952543
transform 1 0 2740 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8289
timestamp 1682952543
transform 1 0 2780 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8326
timestamp 1682952543
transform 1 0 2700 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8327
timestamp 1682952543
transform 1 0 2756 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8328
timestamp 1682952543
transform 1 0 2772 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8156
timestamp 1682952543
transform 1 0 2588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8157
timestamp 1682952543
transform 1 0 2676 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8369
timestamp 1682952543
transform 1 0 2692 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8370
timestamp 1682952543
transform 1 0 2724 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8371
timestamp 1682952543
transform 1 0 2748 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8158
timestamp 1682952543
transform 1 0 2772 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8159
timestamp 1682952543
transform 1 0 2788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8160
timestamp 1682952543
transform 1 0 2796 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8161
timestamp 1682952543
transform 1 0 2812 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8162
timestamp 1682952543
transform 1 0 2820 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8267
timestamp 1682952543
transform 1 0 2564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8268
timestamp 1682952543
transform 1 0 2580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8269
timestamp 1682952543
transform 1 0 2588 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8270
timestamp 1682952543
transform 1 0 2636 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8409
timestamp 1682952543
transform 1 0 2644 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8271
timestamp 1682952543
transform 1 0 2692 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8410
timestamp 1682952543
transform 1 0 2708 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8272
timestamp 1682952543
transform 1 0 2724 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8411
timestamp 1682952543
transform 1 0 2788 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8273
timestamp 1682952543
transform 1 0 2804 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8454
timestamp 1682952543
transform 1 0 2564 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8455
timestamp 1682952543
transform 1 0 2596 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8456
timestamp 1682952543
transform 1 0 2652 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8457
timestamp 1682952543
transform 1 0 2692 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8496
timestamp 1682952543
transform 1 0 2724 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8412
timestamp 1682952543
transform 1 0 2820 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8458
timestamp 1682952543
transform 1 0 2804 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8251
timestamp 1682952543
transform 1 0 2844 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8252
timestamp 1682952543
transform 1 0 2884 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8329
timestamp 1682952543
transform 1 0 2844 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8163
timestamp 1682952543
transform 1 0 2844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8274
timestamp 1682952543
transform 1 0 2892 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8413
timestamp 1682952543
transform 1 0 2908 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8459
timestamp 1682952543
transform 1 0 2828 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8460
timestamp 1682952543
transform 1 0 2876 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8497
timestamp 1682952543
transform 1 0 2924 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8253
timestamp 1682952543
transform 1 0 2940 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8254
timestamp 1682952543
transform 1 0 2980 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8290
timestamp 1682952543
transform 1 0 2948 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8291
timestamp 1682952543
transform 1 0 2964 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8330
timestamp 1682952543
transform 1 0 2972 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8164
timestamp 1682952543
transform 1 0 2972 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8372
timestamp 1682952543
transform 1 0 2980 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8292
timestamp 1682952543
transform 1 0 3020 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8331
timestamp 1682952543
transform 1 0 3028 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8165
timestamp 1682952543
transform 1 0 2988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8166
timestamp 1682952543
transform 1 0 2996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8167
timestamp 1682952543
transform 1 0 3004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8168
timestamp 1682952543
transform 1 0 3020 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8169
timestamp 1682952543
transform 1 0 3036 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8275
timestamp 1682952543
transform 1 0 2956 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8276
timestamp 1682952543
transform 1 0 2964 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8414
timestamp 1682952543
transform 1 0 2972 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8277
timestamp 1682952543
transform 1 0 2980 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8461
timestamp 1682952543
transform 1 0 2964 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8373
timestamp 1682952543
transform 1 0 3044 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8278
timestamp 1682952543
transform 1 0 3012 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8415
timestamp 1682952543
transform 1 0 3020 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8279
timestamp 1682952543
transform 1 0 3028 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8280
timestamp 1682952543
transform 1 0 3044 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8462
timestamp 1682952543
transform 1 0 3028 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8498
timestamp 1682952543
transform 1 0 3004 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8499
timestamp 1682952543
transform 1 0 3036 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_8332
timestamp 1682952543
transform 1 0 3092 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8333
timestamp 1682952543
transform 1 0 3140 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8170
timestamp 1682952543
transform 1 0 3140 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8416
timestamp 1682952543
transform 1 0 3068 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8281
timestamp 1682952543
transform 1 0 3092 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8463
timestamp 1682952543
transform 1 0 3076 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8255
timestamp 1682952543
transform 1 0 3172 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8256
timestamp 1682952543
transform 1 0 3196 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8257
timestamp 1682952543
transform 1 0 3220 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8293
timestamp 1682952543
transform 1 0 3244 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8334
timestamp 1682952543
transform 1 0 3164 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8335
timestamp 1682952543
transform 1 0 3188 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8171
timestamp 1682952543
transform 1 0 3164 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8374
timestamp 1682952543
transform 1 0 3188 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8375
timestamp 1682952543
transform 1 0 3204 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8376
timestamp 1682952543
transform 1 0 3244 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8282
timestamp 1682952543
transform 1 0 3196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8283
timestamp 1682952543
transform 1 0 3244 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8284
timestamp 1682952543
transform 1 0 3252 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8258
timestamp 1682952543
transform 1 0 3276 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8294
timestamp 1682952543
transform 1 0 3316 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8172
timestamp 1682952543
transform 1 0 3300 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8377
timestamp 1682952543
transform 1 0 3308 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8336
timestamp 1682952543
transform 1 0 3340 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8173
timestamp 1682952543
transform 1 0 3332 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8285
timestamp 1682952543
transform 1 0 3308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8286
timestamp 1682952543
transform 1 0 3324 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8417
timestamp 1682952543
transform 1 0 3332 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8378
timestamp 1682952543
transform 1 0 3364 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8287
timestamp 1682952543
transform 1 0 3364 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8317
timestamp 1682952543
transform 1 0 3348 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8319
timestamp 1682952543
transform 1 0 3356 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_8484
timestamp 1682952543
transform 1 0 3356 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_8259
timestamp 1682952543
transform 1 0 3396 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8295
timestamp 1682952543
transform 1 0 3388 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8337
timestamp 1682952543
transform 1 0 3380 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8174
timestamp 1682952543
transform 1 0 3380 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8338
timestamp 1682952543
transform 1 0 3412 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8260
timestamp 1682952543
transform 1 0 3436 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8175
timestamp 1682952543
transform 1 0 3412 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8176
timestamp 1682952543
transform 1 0 3428 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8418
timestamp 1682952543
transform 1 0 3396 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8288
timestamp 1682952543
transform 1 0 3404 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8289
timestamp 1682952543
transform 1 0 3420 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8290
timestamp 1682952543
transform 1 0 3428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8318
timestamp 1682952543
transform 1 0 3388 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_8464
timestamp 1682952543
transform 1 0 3388 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8261
timestamp 1682952543
transform 1 0 3452 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8262
timestamp 1682952543
transform 1 0 3516 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8339
timestamp 1682952543
transform 1 0 3476 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8177
timestamp 1682952543
transform 1 0 3524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8291
timestamp 1682952543
transform 1 0 3476 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8465
timestamp 1682952543
transform 1 0 3452 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_8263
timestamp 1682952543
transform 1 0 3628 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8340
timestamp 1682952543
transform 1 0 3596 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8178
timestamp 1682952543
transform 1 0 3548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8292
timestamp 1682952543
transform 1 0 3596 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8429
timestamp 1682952543
transform 1 0 3628 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8264
timestamp 1682952543
transform 1 0 3660 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8296
timestamp 1682952543
transform 1 0 3668 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8297
timestamp 1682952543
transform 1 0 3692 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8341
timestamp 1682952543
transform 1 0 3676 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8179
timestamp 1682952543
transform 1 0 3660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8180
timestamp 1682952543
transform 1 0 3676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8181
timestamp 1682952543
transform 1 0 3692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8182
timestamp 1682952543
transform 1 0 3700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8293
timestamp 1682952543
transform 1 0 3660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8294
timestamp 1682952543
transform 1 0 3668 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8295
timestamp 1682952543
transform 1 0 3684 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8430
timestamp 1682952543
transform 1 0 3660 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8431
timestamp 1682952543
transform 1 0 3684 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8296
timestamp 1682952543
transform 1 0 3700 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8265
timestamp 1682952543
transform 1 0 3716 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8342
timestamp 1682952543
transform 1 0 3732 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8183
timestamp 1682952543
transform 1 0 3716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8184
timestamp 1682952543
transform 1 0 3732 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8185
timestamp 1682952543
transform 1 0 3748 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8419
timestamp 1682952543
transform 1 0 3716 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8297
timestamp 1682952543
transform 1 0 3724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8298
timestamp 1682952543
transform 1 0 3740 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8298
timestamp 1682952543
transform 1 0 3772 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8299
timestamp 1682952543
transform 1 0 3788 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8343
timestamp 1682952543
transform 1 0 3796 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8186
timestamp 1682952543
transform 1 0 3772 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8379
timestamp 1682952543
transform 1 0 3836 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8420
timestamp 1682952543
transform 1 0 3772 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8299
timestamp 1682952543
transform 1 0 3796 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8421
timestamp 1682952543
transform 1 0 3804 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_8432
timestamp 1682952543
transform 1 0 3804 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_8266
timestamp 1682952543
transform 1 0 3868 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8079
timestamp 1682952543
transform 1 0 3868 0 1 755
box -2 -2 2 2
use M3_M2  M3_M2_8267
timestamp 1682952543
transform 1 0 3884 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8300
timestamp 1682952543
transform 1 0 3892 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8344
timestamp 1682952543
transform 1 0 3892 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8380
timestamp 1682952543
transform 1 0 3876 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8187
timestamp 1682952543
transform 1 0 3892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8300
timestamp 1682952543
transform 1 0 3868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8301
timestamp 1682952543
transform 1 0 3876 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8302
timestamp 1682952543
transform 1 0 3884 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8303
timestamp 1682952543
transform 1 0 3900 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8433
timestamp 1682952543
transform 1 0 3860 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8188
timestamp 1682952543
transform 1 0 3916 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8268
timestamp 1682952543
transform 1 0 3940 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_8269
timestamp 1682952543
transform 1 0 3980 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8189
timestamp 1682952543
transform 1 0 3932 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8301
timestamp 1682952543
transform 1 0 3948 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_8345
timestamp 1682952543
transform 1 0 3972 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_8346
timestamp 1682952543
transform 1 0 4012 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8190
timestamp 1682952543
transform 1 0 3948 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_8381
timestamp 1682952543
transform 1 0 3988 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_8382
timestamp 1682952543
transform 1 0 4028 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8304
timestamp 1682952543
transform 1 0 3972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8305
timestamp 1682952543
transform 1 0 4028 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_8347
timestamp 1682952543
transform 1 0 4092 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8191
timestamp 1682952543
transform 1 0 4068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8306
timestamp 1682952543
transform 1 0 4092 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8307
timestamp 1682952543
transform 1 0 4148 0 1 725
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_68
timestamp 1682952543
transform 1 0 24 0 1 670
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_492
timestamp 1682952543
transform 1 0 72 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_493
timestamp 1682952543
transform 1 0 168 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_565
timestamp 1682952543
transform 1 0 264 0 -1 770
box -9 -3 26 105
use FILL  FILL_3561
timestamp 1682952543
transform 1 0 280 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_497
timestamp 1682952543
transform 1 0 288 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_568
timestamp 1682952543
transform -1 0 400 0 -1 770
box -9 -3 26 105
use FILL  FILL_3581
timestamp 1682952543
transform 1 0 400 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_329
timestamp 1682952543
transform -1 0 448 0 -1 770
box -8 -3 46 105
use FILL  FILL_3582
timestamp 1682952543
transform 1 0 448 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_8500
timestamp 1682952543
transform 1 0 468 0 1 675
box -3 -3 3 3
use FILL  FILL_3583
timestamp 1682952543
transform 1 0 456 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_330
timestamp 1682952543
transform 1 0 464 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_353
timestamp 1682952543
transform 1 0 504 0 -1 770
box -8 -3 46 105
use FILL  FILL_3584
timestamp 1682952543
transform 1 0 544 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_354
timestamp 1682952543
transform -1 0 592 0 -1 770
box -8 -3 46 105
use AOI22X1  AOI22X1_331
timestamp 1682952543
transform 1 0 592 0 -1 770
box -8 -3 46 105
use FILL  FILL_3585
timestamp 1682952543
transform 1 0 632 0 -1 770
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1682952543
transform 1 0 640 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_498
timestamp 1682952543
transform 1 0 648 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_569
timestamp 1682952543
transform -1 0 760 0 -1 770
box -9 -3 26 105
use FILL  FILL_3587
timestamp 1682952543
transform 1 0 760 0 -1 770
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1682952543
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1682952543
transform 1 0 776 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_332
timestamp 1682952543
transform -1 0 824 0 -1 770
box -8 -3 46 105
use FILL  FILL_3590
timestamp 1682952543
transform 1 0 824 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_136
timestamp 1682952543
transform 1 0 832 0 -1 770
box -8 -3 34 105
use M3_M2  M3_M2_8501
timestamp 1682952543
transform 1 0 876 0 1 675
box -3 -3 3 3
use FILL  FILL_3591
timestamp 1682952543
transform 1 0 864 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_333
timestamp 1682952543
transform 1 0 872 0 -1 770
box -8 -3 46 105
use FILL  FILL_3592
timestamp 1682952543
transform 1 0 912 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_137
timestamp 1682952543
transform 1 0 920 0 -1 770
box -8 -3 34 105
use FILL  FILL_3593
timestamp 1682952543
transform 1 0 952 0 -1 770
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1682952543
transform 1 0 960 0 -1 770
box -8 -3 16 105
use FILL  FILL_3637
timestamp 1682952543
transform 1 0 968 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_143
timestamp 1682952543
transform -1 0 1008 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_144
timestamp 1682952543
transform -1 0 1040 0 -1 770
box -8 -3 34 105
use FILL  FILL_3638
timestamp 1682952543
transform 1 0 1040 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_145
timestamp 1682952543
transform -1 0 1080 0 -1 770
box -8 -3 34 105
use FILL  FILL_3639
timestamp 1682952543
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1682952543
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1682952543
transform 1 0 1096 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_8502
timestamp 1682952543
transform 1 0 1116 0 1 675
box -3 -3 3 3
use INVX2  INVX2_581
timestamp 1682952543
transform 1 0 1104 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_582
timestamp 1682952543
transform 1 0 1120 0 -1 770
box -9 -3 26 105
use OAI22X1  OAI22X1_365
timestamp 1682952543
transform -1 0 1176 0 -1 770
box -8 -3 46 105
use FILL  FILL_3642
timestamp 1682952543
transform 1 0 1176 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_366
timestamp 1682952543
transform -1 0 1224 0 -1 770
box -8 -3 46 105
use FILL  FILL_3643
timestamp 1682952543
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_512
timestamp 1682952543
transform 1 0 1232 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_513
timestamp 1682952543
transform -1 0 1424 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_514
timestamp 1682952543
transform 1 0 1424 0 -1 770
box -8 -3 104 105
use FILL  FILL_3644
timestamp 1682952543
transform 1 0 1520 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_583
timestamp 1682952543
transform -1 0 1544 0 -1 770
box -9 -3 26 105
use FILL  FILL_3645
timestamp 1682952543
transform 1 0 1544 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_340
timestamp 1682952543
transform 1 0 1552 0 -1 770
box -8 -3 46 105
use FILL  FILL_3646
timestamp 1682952543
transform 1 0 1592 0 -1 770
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1682952543
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_584
timestamp 1682952543
transform 1 0 1608 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_585
timestamp 1682952543
transform -1 0 1640 0 -1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_341
timestamp 1682952543
transform 1 0 1640 0 -1 770
box -8 -3 46 105
use FILL  FILL_3648
timestamp 1682952543
transform 1 0 1680 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_586
timestamp 1682952543
transform 1 0 1688 0 -1 770
box -9 -3 26 105
use FILL  FILL_3649
timestamp 1682952543
transform 1 0 1704 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_8503
timestamp 1682952543
transform 1 0 1796 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_515
timestamp 1682952543
transform -1 0 1808 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_587
timestamp 1682952543
transform -1 0 1824 0 -1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_342
timestamp 1682952543
transform 1 0 1824 0 -1 770
box -8 -3 46 105
use FILL  FILL_3650
timestamp 1682952543
transform 1 0 1864 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_588
timestamp 1682952543
transform 1 0 1872 0 -1 770
box -9 -3 26 105
use OAI21X1  OAI21X1_146
timestamp 1682952543
transform 1 0 1888 0 -1 770
box -8 -3 34 105
use FILL  FILL_3651
timestamp 1682952543
transform 1 0 1920 0 -1 770
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1682952543
transform 1 0 1928 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_147
timestamp 1682952543
transform -1 0 1968 0 -1 770
box -8 -3 34 105
use FILL  FILL_3653
timestamp 1682952543
transform 1 0 1968 0 -1 770
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1682952543
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1682952543
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_367
timestamp 1682952543
transform 1 0 1992 0 -1 770
box -8 -3 46 105
use FILL  FILL_3656
timestamp 1682952543
transform 1 0 2032 0 -1 770
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1682952543
transform 1 0 2040 0 -1 770
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1682952543
transform 1 0 2048 0 -1 770
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1682952543
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1682952543
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_589
timestamp 1682952543
transform -1 0 2088 0 -1 770
box -9 -3 26 105
use FILL  FILL_3661
timestamp 1682952543
transform 1 0 2088 0 -1 770
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1682952543
transform 1 0 2096 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_516
timestamp 1682952543
transform 1 0 2104 0 -1 770
box -8 -3 104 105
use FILL  FILL_3663
timestamp 1682952543
transform 1 0 2200 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_517
timestamp 1682952543
transform -1 0 2304 0 -1 770
box -8 -3 104 105
use FILL  FILL_3664
timestamp 1682952543
transform 1 0 2304 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_368
timestamp 1682952543
transform 1 0 2312 0 -1 770
box -8 -3 46 105
use FILL  FILL_3665
timestamp 1682952543
transform 1 0 2352 0 -1 770
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1682952543
transform 1 0 2360 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_518
timestamp 1682952543
transform 1 0 2368 0 -1 770
box -8 -3 104 105
use OAI21X1  OAI21X1_148
timestamp 1682952543
transform 1 0 2464 0 -1 770
box -8 -3 34 105
use NOR2X1  NOR2X1_99
timestamp 1682952543
transform -1 0 2520 0 -1 770
box -8 -3 32 105
use INVX2  INVX2_590
timestamp 1682952543
transform -1 0 2536 0 -1 770
box -9 -3 26 105
use FILL  FILL_3667
timestamp 1682952543
transform 1 0 2536 0 -1 770
box -8 -3 16 105
use FILL  FILL_3668
timestamp 1682952543
transform 1 0 2544 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_369
timestamp 1682952543
transform -1 0 2592 0 -1 770
box -8 -3 46 105
use M3_M2  M3_M2_8504
timestamp 1682952543
transform 1 0 2684 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_519
timestamp 1682952543
transform -1 0 2688 0 -1 770
box -8 -3 104 105
use M3_M2  M3_M2_8505
timestamp 1682952543
transform 1 0 2700 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_520
timestamp 1682952543
transform -1 0 2784 0 -1 770
box -8 -3 104 105
use AOI22X1  AOI22X1_343
timestamp 1682952543
transform 1 0 2784 0 -1 770
box -8 -3 46 105
use FILL  FILL_3669
timestamp 1682952543
transform 1 0 2824 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_521
timestamp 1682952543
transform 1 0 2832 0 -1 770
box -8 -3 104 105
use FILL  FILL_3670
timestamp 1682952543
transform 1 0 2928 0 -1 770
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1682952543
transform 1 0 2936 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_591
timestamp 1682952543
transform 1 0 2944 0 -1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_344
timestamp 1682952543
transform 1 0 2960 0 -1 770
box -8 -3 46 105
use OAI22X1  OAI22X1_370
timestamp 1682952543
transform 1 0 3000 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_592
timestamp 1682952543
transform -1 0 3056 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_522
timestamp 1682952543
transform -1 0 3152 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_523
timestamp 1682952543
transform 1 0 3152 0 -1 770
box -8 -3 104 105
use FILL  FILL_3672
timestamp 1682952543
transform 1 0 3248 0 -1 770
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1682952543
transform 1 0 3256 0 -1 770
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1682952543
transform 1 0 3264 0 -1 770
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1682952543
transform 1 0 3272 0 -1 770
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1682952543
transform 1 0 3280 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_345
timestamp 1682952543
transform -1 0 3328 0 -1 770
box -8 -3 46 105
use FILL  FILL_3677
timestamp 1682952543
transform 1 0 3328 0 -1 770
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1682952543
transform 1 0 3336 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_68
timestamp 1682952543
transform -1 0 3376 0 -1 770
box -8 -3 40 105
use FILL  FILL_3679
timestamp 1682952543
transform 1 0 3376 0 -1 770
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1682952543
transform 1 0 3384 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_371
timestamp 1682952543
transform -1 0 3432 0 -1 770
box -8 -3 46 105
use FILL  FILL_3681
timestamp 1682952543
transform 1 0 3432 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_524
timestamp 1682952543
transform -1 0 3536 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_525
timestamp 1682952543
transform 1 0 3536 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_593
timestamp 1682952543
transform 1 0 3632 0 -1 770
box -9 -3 26 105
use FILL  FILL_3685
timestamp 1682952543
transform 1 0 3648 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_373
timestamp 1682952543
transform 1 0 3656 0 -1 770
box -8 -3 46 105
use FILL  FILL_3688
timestamp 1682952543
transform 1 0 3696 0 -1 770
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1682952543
transform 1 0 3704 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_8506
timestamp 1682952543
transform 1 0 3756 0 1 675
box -3 -3 3 3
use OAI22X1  OAI22X1_375
timestamp 1682952543
transform 1 0 3712 0 -1 770
box -8 -3 46 105
use FILL  FILL_3701
timestamp 1682952543
transform 1 0 3752 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_528
timestamp 1682952543
transform 1 0 3760 0 -1 770
box -8 -3 104 105
use FILL  FILL_3702
timestamp 1682952543
transform 1 0 3856 0 -1 770
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1682952543
transform 1 0 3864 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_376
timestamp 1682952543
transform 1 0 3872 0 -1 770
box -8 -3 46 105
use FILL  FILL_3704
timestamp 1682952543
transform 1 0 3912 0 -1 770
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1682952543
transform 1 0 3920 0 -1 770
box -8 -3 16 105
use FILL  FILL_3706
timestamp 1682952543
transform 1 0 3928 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_529
timestamp 1682952543
transform 1 0 3936 0 -1 770
box -8 -3 104 105
use FILL  FILL_3707
timestamp 1682952543
transform 1 0 4032 0 -1 770
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1682952543
transform 1 0 4040 0 -1 770
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1682952543
transform 1 0 4048 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_530
timestamp 1682952543
transform 1 0 4056 0 -1 770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_69
timestamp 1682952543
transform 1 0 4201 0 1 670
box -10 -3 10 3
use M2_M1  M2_M1_8331
timestamp 1682952543
transform 1 0 124 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8688
timestamp 1682952543
transform 1 0 116 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8581
timestamp 1682952543
transform 1 0 148 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8332
timestamp 1682952543
transform 1 0 140 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8667
timestamp 1682952543
transform 1 0 140 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8460
timestamp 1682952543
transform 1 0 148 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8532
timestamp 1682952543
transform 1 0 188 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8582
timestamp 1682952543
transform 1 0 172 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8639
timestamp 1682952543
transform 1 0 164 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8533
timestamp 1682952543
transform 1 0 284 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8534
timestamp 1682952543
transform 1 0 300 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8551
timestamp 1682952543
transform 1 0 252 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8583
timestamp 1682952543
transform 1 0 252 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8584
timestamp 1682952543
transform 1 0 292 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8333
timestamp 1682952543
transform 1 0 172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8334
timestamp 1682952543
transform 1 0 188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8335
timestamp 1682952543
transform 1 0 252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8336
timestamp 1682952543
transform 1 0 284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8337
timestamp 1682952543
transform 1 0 292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8338
timestamp 1682952543
transform 1 0 300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8461
timestamp 1682952543
transform 1 0 164 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8668
timestamp 1682952543
transform 1 0 172 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8462
timestamp 1682952543
transform 1 0 188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8463
timestamp 1682952543
transform 1 0 204 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8689
timestamp 1682952543
transform 1 0 252 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8690
timestamp 1682952543
transform 1 0 284 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8552
timestamp 1682952543
transform 1 0 324 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8553
timestamp 1682952543
transform 1 0 356 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8585
timestamp 1682952543
transform 1 0 348 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8339
timestamp 1682952543
transform 1 0 332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8340
timestamp 1682952543
transform 1 0 348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8464
timestamp 1682952543
transform 1 0 316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8465
timestamp 1682952543
transform 1 0 324 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8466
timestamp 1682952543
transform 1 0 340 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8691
timestamp 1682952543
transform 1 0 340 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8467
timestamp 1682952543
transform 1 0 356 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8554
timestamp 1682952543
transform 1 0 436 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8586
timestamp 1682952543
transform 1 0 396 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8587
timestamp 1682952543
transform 1 0 444 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8588
timestamp 1682952543
transform 1 0 484 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8341
timestamp 1682952543
transform 1 0 444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8342
timestamp 1682952543
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8343
timestamp 1682952543
transform 1 0 484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8468
timestamp 1682952543
transform 1 0 396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8469
timestamp 1682952543
transform 1 0 484 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8470
timestamp 1682952543
transform 1 0 500 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8692
timestamp 1682952543
transform 1 0 500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8589
timestamp 1682952543
transform 1 0 532 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8344
timestamp 1682952543
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8345
timestamp 1682952543
transform 1 0 532 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8640
timestamp 1682952543
transform 1 0 540 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8669
timestamp 1682952543
transform 1 0 516 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8471
timestamp 1682952543
transform 1 0 524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8472
timestamp 1682952543
transform 1 0 540 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8473
timestamp 1682952543
transform 1 0 548 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8670
timestamp 1682952543
transform 1 0 556 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8507
timestamp 1682952543
transform 1 0 572 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8516
timestamp 1682952543
transform 1 0 588 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8590
timestamp 1682952543
transform 1 0 572 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8346
timestamp 1682952543
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8347
timestamp 1682952543
transform 1 0 588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8474
timestamp 1682952543
transform 1 0 580 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8671
timestamp 1682952543
transform 1 0 588 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8475
timestamp 1682952543
transform 1 0 596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8476
timestamp 1682952543
transform 1 0 604 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8693
timestamp 1682952543
transform 1 0 580 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8591
timestamp 1682952543
transform 1 0 620 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8517
timestamp 1682952543
transform 1 0 692 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8592
timestamp 1682952543
transform 1 0 660 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8348
timestamp 1682952543
transform 1 0 620 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8349
timestamp 1682952543
transform 1 0 628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8350
timestamp 1682952543
transform 1 0 660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8477
timestamp 1682952543
transform 1 0 708 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8730
timestamp 1682952543
transform 1 0 668 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8535
timestamp 1682952543
transform 1 0 732 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8351
timestamp 1682952543
transform 1 0 732 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8555
timestamp 1682952543
transform 1 0 764 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8641
timestamp 1682952543
transform 1 0 748 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8352
timestamp 1682952543
transform 1 0 756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8353
timestamp 1682952543
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8478
timestamp 1682952543
transform 1 0 748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8479
timestamp 1682952543
transform 1 0 764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8480
timestamp 1682952543
transform 1 0 772 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8731
timestamp 1682952543
transform 1 0 764 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8354
timestamp 1682952543
transform 1 0 788 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8585
timestamp 1682952543
transform 1 0 796 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_8642
timestamp 1682952543
transform 1 0 812 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8556
timestamp 1682952543
transform 1 0 828 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8557
timestamp 1682952543
transform 1 0 844 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8593
timestamp 1682952543
transform 1 0 836 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8536
timestamp 1682952543
transform 1 0 884 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8320
timestamp 1682952543
transform 1 0 868 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_8594
timestamp 1682952543
transform 1 0 868 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8355
timestamp 1682952543
transform 1 0 836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8356
timestamp 1682952543
transform 1 0 844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8357
timestamp 1682952543
transform 1 0 860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8481
timestamp 1682952543
transform 1 0 820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8482
timestamp 1682952543
transform 1 0 828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8483
timestamp 1682952543
transform 1 0 836 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8643
timestamp 1682952543
transform 1 0 876 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8484
timestamp 1682952543
transform 1 0 868 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8672
timestamp 1682952543
transform 1 0 876 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8586
timestamp 1682952543
transform 1 0 876 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_8537
timestamp 1682952543
transform 1 0 908 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8558
timestamp 1682952543
transform 1 0 932 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8595
timestamp 1682952543
transform 1 0 908 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8596
timestamp 1682952543
transform 1 0 948 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8358
timestamp 1682952543
transform 1 0 892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8359
timestamp 1682952543
transform 1 0 908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8360
timestamp 1682952543
transform 1 0 916 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8361
timestamp 1682952543
transform 1 0 948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8485
timestamp 1682952543
transform 1 0 900 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8486
timestamp 1682952543
transform 1 0 996 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8694
timestamp 1682952543
transform 1 0 980 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8644
timestamp 1682952543
transform 1 0 1012 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8487
timestamp 1682952543
transform 1 0 1012 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8597
timestamp 1682952543
transform 1 0 1028 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8322
timestamp 1682952543
transform 1 0 1044 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_8559
timestamp 1682952543
transform 1 0 1068 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8598
timestamp 1682952543
transform 1 0 1068 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8362
timestamp 1682952543
transform 1 0 1068 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8695
timestamp 1682952543
transform 1 0 1052 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8560
timestamp 1682952543
transform 1 0 1124 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8363
timestamp 1682952543
transform 1 0 1092 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8364
timestamp 1682952543
transform 1 0 1148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8488
timestamp 1682952543
transform 1 0 1084 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8673
timestamp 1682952543
transform 1 0 1092 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8489
timestamp 1682952543
transform 1 0 1172 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8696
timestamp 1682952543
transform 1 0 1140 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8365
timestamp 1682952543
transform 1 0 1196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8490
timestamp 1682952543
transform 1 0 1188 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8697
timestamp 1682952543
transform 1 0 1188 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8366
timestamp 1682952543
transform 1 0 1212 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8674
timestamp 1682952543
transform 1 0 1212 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8367
timestamp 1682952543
transform 1 0 1300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8491
timestamp 1682952543
transform 1 0 1252 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8675
timestamp 1682952543
transform 1 0 1300 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8599
timestamp 1682952543
transform 1 0 1396 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8368
timestamp 1682952543
transform 1 0 1348 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8369
timestamp 1682952543
transform 1 0 1364 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8370
timestamp 1682952543
transform 1 0 1380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8371
timestamp 1682952543
transform 1 0 1396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8492
timestamp 1682952543
transform 1 0 1356 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8676
timestamp 1682952543
transform 1 0 1364 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8493
timestamp 1682952543
transform 1 0 1372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8494
timestamp 1682952543
transform 1 0 1388 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8677
timestamp 1682952543
transform 1 0 1396 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8561
timestamp 1682952543
transform 1 0 1484 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8600
timestamp 1682952543
transform 1 0 1468 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8601
timestamp 1682952543
transform 1 0 1508 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8562
timestamp 1682952543
transform 1 0 1532 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8508
timestamp 1682952543
transform 1 0 1588 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8518
timestamp 1682952543
transform 1 0 1572 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8602
timestamp 1682952543
transform 1 0 1532 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8603
timestamp 1682952543
transform 1 0 1564 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8604
timestamp 1682952543
transform 1 0 1588 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8372
timestamp 1682952543
transform 1 0 1468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8373
timestamp 1682952543
transform 1 0 1500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8374
timestamp 1682952543
transform 1 0 1508 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8495
timestamp 1682952543
transform 1 0 1404 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8496
timestamp 1682952543
transform 1 0 1420 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8645
timestamp 1682952543
transform 1 0 1516 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8375
timestamp 1682952543
transform 1 0 1524 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8646
timestamp 1682952543
transform 1 0 1532 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8519
timestamp 1682952543
transform 1 0 1612 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8605
timestamp 1682952543
transform 1 0 1628 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8376
timestamp 1682952543
transform 1 0 1540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8377
timestamp 1682952543
transform 1 0 1556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8378
timestamp 1682952543
transform 1 0 1564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8379
timestamp 1682952543
transform 1 0 1572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8380
timestamp 1682952543
transform 1 0 1588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8497
timestamp 1682952543
transform 1 0 1524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8498
timestamp 1682952543
transform 1 0 1532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8499
timestamp 1682952543
transform 1 0 1548 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8698
timestamp 1682952543
transform 1 0 1500 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8699
timestamp 1682952543
transform 1 0 1548 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8647
timestamp 1682952543
transform 1 0 1604 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8381
timestamp 1682952543
transform 1 0 1612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8382
timestamp 1682952543
transform 1 0 1628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8500
timestamp 1682952543
transform 1 0 1580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8501
timestamp 1682952543
transform 1 0 1596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8502
timestamp 1682952543
transform 1 0 1604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8503
timestamp 1682952543
transform 1 0 1620 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8504
timestamp 1682952543
transform 1 0 1636 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8505
timestamp 1682952543
transform 1 0 1644 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8732
timestamp 1682952543
transform 1 0 1580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8700
timestamp 1682952543
transform 1 0 1636 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8606
timestamp 1682952543
transform 1 0 1652 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8607
timestamp 1682952543
transform 1 0 1676 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8383
timestamp 1682952543
transform 1 0 1652 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8384
timestamp 1682952543
transform 1 0 1660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8385
timestamp 1682952543
transform 1 0 1700 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8648
timestamp 1682952543
transform 1 0 1716 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8506
timestamp 1682952543
transform 1 0 1740 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8701
timestamp 1682952543
transform 1 0 1660 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8520
timestamp 1682952543
transform 1 0 1804 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8521
timestamp 1682952543
transform 1 0 1820 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8386
timestamp 1682952543
transform 1 0 1804 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8507
timestamp 1682952543
transform 1 0 1764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8387
timestamp 1682952543
transform 1 0 1868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8388
timestamp 1682952543
transform 1 0 1876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8323
timestamp 1682952543
transform 1 0 1908 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_8649
timestamp 1682952543
transform 1 0 1908 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8587
timestamp 1682952543
transform 1 0 1900 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_8733
timestamp 1682952543
transform 1 0 1900 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8508
timestamp 1682952543
transform 1 0 1916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8324
timestamp 1682952543
transform 1 0 1940 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8389
timestamp 1682952543
transform 1 0 1932 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8650
timestamp 1682952543
transform 1 0 1940 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8509
timestamp 1682952543
transform 1 0 1940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8588
timestamp 1682952543
transform 1 0 1964 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_8734
timestamp 1682952543
transform 1 0 1956 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8325
timestamp 1682952543
transform 1 0 1972 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8390
timestamp 1682952543
transform 1 0 1988 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8702
timestamp 1682952543
transform 1 0 1972 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8735
timestamp 1682952543
transform 1 0 1988 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8510
timestamp 1682952543
transform 1 0 2004 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8703
timestamp 1682952543
transform 1 0 2004 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8391
timestamp 1682952543
transform 1 0 2020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8511
timestamp 1682952543
transform 1 0 2044 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8736
timestamp 1682952543
transform 1 0 2044 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8608
timestamp 1682952543
transform 1 0 2076 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8609
timestamp 1682952543
transform 1 0 2140 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8610
timestamp 1682952543
transform 1 0 2188 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8392
timestamp 1682952543
transform 1 0 2060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8393
timestamp 1682952543
transform 1 0 2076 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8394
timestamp 1682952543
transform 1 0 2084 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8395
timestamp 1682952543
transform 1 0 2124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8396
timestamp 1682952543
transform 1 0 2188 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8512
timestamp 1682952543
transform 1 0 2068 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8678
timestamp 1682952543
transform 1 0 2076 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8513
timestamp 1682952543
transform 1 0 2084 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8514
timestamp 1682952543
transform 1 0 2172 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8515
timestamp 1682952543
transform 1 0 2188 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8704
timestamp 1682952543
transform 1 0 2068 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8705
timestamp 1682952543
transform 1 0 2124 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8737
timestamp 1682952543
transform 1 0 2100 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8738
timestamp 1682952543
transform 1 0 2188 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8679
timestamp 1682952543
transform 1 0 2204 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8563
timestamp 1682952543
transform 1 0 2244 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8397
timestamp 1682952543
transform 1 0 2236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8516
timestamp 1682952543
transform 1 0 2212 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8517
timestamp 1682952543
transform 1 0 2228 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8518
timestamp 1682952543
transform 1 0 2244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8519
timestamp 1682952543
transform 1 0 2252 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8706
timestamp 1682952543
transform 1 0 2236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8739
timestamp 1682952543
transform 1 0 2244 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8520
timestamp 1682952543
transform 1 0 2268 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8707
timestamp 1682952543
transform 1 0 2268 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8611
timestamp 1682952543
transform 1 0 2292 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8564
timestamp 1682952543
transform 1 0 2316 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8538
timestamp 1682952543
transform 1 0 2332 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8565
timestamp 1682952543
transform 1 0 2356 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8326
timestamp 1682952543
transform 1 0 2316 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_8612
timestamp 1682952543
transform 1 0 2324 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8613
timestamp 1682952543
transform 1 0 2340 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8327
timestamp 1682952543
transform 1 0 2356 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8398
timestamp 1682952543
transform 1 0 2292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8399
timestamp 1682952543
transform 1 0 2300 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8400
timestamp 1682952543
transform 1 0 2316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8521
timestamp 1682952543
transform 1 0 2316 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8708
timestamp 1682952543
transform 1 0 2308 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8401
timestamp 1682952543
transform 1 0 2340 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8522
timestamp 1682952543
transform 1 0 2324 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8740
timestamp 1682952543
transform 1 0 2348 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8651
timestamp 1682952543
transform 1 0 2372 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8539
timestamp 1682952543
transform 1 0 2420 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8402
timestamp 1682952543
transform 1 0 2388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8403
timestamp 1682952543
transform 1 0 2412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8404
timestamp 1682952543
transform 1 0 2428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8523
timestamp 1682952543
transform 1 0 2372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8524
timestamp 1682952543
transform 1 0 2380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8525
timestamp 1682952543
transform 1 0 2396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8526
timestamp 1682952543
transform 1 0 2404 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8709
timestamp 1682952543
transform 1 0 2380 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8710
timestamp 1682952543
transform 1 0 2412 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8741
timestamp 1682952543
transform 1 0 2396 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8405
timestamp 1682952543
transform 1 0 2444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8527
timestamp 1682952543
transform 1 0 2444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8328
timestamp 1682952543
transform 1 0 2476 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8406
timestamp 1682952543
transform 1 0 2460 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8652
timestamp 1682952543
transform 1 0 2492 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8509
timestamp 1682952543
transform 1 0 2516 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8510
timestamp 1682952543
transform 1 0 2540 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8540
timestamp 1682952543
transform 1 0 2524 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8566
timestamp 1682952543
transform 1 0 2532 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8653
timestamp 1682952543
transform 1 0 2508 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8511
timestamp 1682952543
transform 1 0 2580 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8541
timestamp 1682952543
transform 1 0 2572 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8567
timestamp 1682952543
transform 1 0 2564 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8542
timestamp 1682952543
transform 1 0 2604 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8614
timestamp 1682952543
transform 1 0 2556 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8615
timestamp 1682952543
transform 1 0 2588 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8407
timestamp 1682952543
transform 1 0 2516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8408
timestamp 1682952543
transform 1 0 2532 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8409
timestamp 1682952543
transform 1 0 2548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8410
timestamp 1682952543
transform 1 0 2564 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8528
timestamp 1682952543
transform 1 0 2500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8529
timestamp 1682952543
transform 1 0 2508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8530
timestamp 1682952543
transform 1 0 2524 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8711
timestamp 1682952543
transform 1 0 2500 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8411
timestamp 1682952543
transform 1 0 2604 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8654
timestamp 1682952543
transform 1 0 2612 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8568
timestamp 1682952543
transform 1 0 2684 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8616
timestamp 1682952543
transform 1 0 2660 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8412
timestamp 1682952543
transform 1 0 2628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8413
timestamp 1682952543
transform 1 0 2636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8414
timestamp 1682952543
transform 1 0 2660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8531
timestamp 1682952543
transform 1 0 2556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8532
timestamp 1682952543
transform 1 0 2572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8533
timestamp 1682952543
transform 1 0 2580 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8534
timestamp 1682952543
transform 1 0 2596 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8535
timestamp 1682952543
transform 1 0 2612 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8536
timestamp 1682952543
transform 1 0 2620 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8712
timestamp 1682952543
transform 1 0 2540 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8713
timestamp 1682952543
transform 1 0 2564 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8742
timestamp 1682952543
transform 1 0 2580 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8714
timestamp 1682952543
transform 1 0 2620 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8537
timestamp 1682952543
transform 1 0 2644 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8743
timestamp 1682952543
transform 1 0 2628 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8512
timestamp 1682952543
transform 1 0 2732 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8513
timestamp 1682952543
transform 1 0 2764 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8514
timestamp 1682952543
transform 1 0 2796 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8522
timestamp 1682952543
transform 1 0 2740 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8523
timestamp 1682952543
transform 1 0 2796 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8543
timestamp 1682952543
transform 1 0 2708 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8544
timestamp 1682952543
transform 1 0 2772 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8617
timestamp 1682952543
transform 1 0 2692 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8415
timestamp 1682952543
transform 1 0 2692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8538
timestamp 1682952543
transform 1 0 2684 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8618
timestamp 1682952543
transform 1 0 2772 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8416
timestamp 1682952543
transform 1 0 2772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8539
timestamp 1682952543
transform 1 0 2708 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8540
timestamp 1682952543
transform 1 0 2724 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8715
timestamp 1682952543
transform 1 0 2708 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8744
timestamp 1682952543
transform 1 0 2756 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8524
timestamp 1682952543
transform 1 0 2828 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8545
timestamp 1682952543
transform 1 0 2820 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8546
timestamp 1682952543
transform 1 0 2836 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8619
timestamp 1682952543
transform 1 0 2844 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8417
timestamp 1682952543
transform 1 0 2820 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8418
timestamp 1682952543
transform 1 0 2836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8541
timestamp 1682952543
transform 1 0 2828 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8542
timestamp 1682952543
transform 1 0 2844 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8680
timestamp 1682952543
transform 1 0 2852 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8419
timestamp 1682952543
transform 1 0 2868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8543
timestamp 1682952543
transform 1 0 2860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8544
timestamp 1682952543
transform 1 0 2868 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8525
timestamp 1682952543
transform 1 0 2884 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8655
timestamp 1682952543
transform 1 0 2908 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8420
timestamp 1682952543
transform 1 0 2916 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8545
timestamp 1682952543
transform 1 0 2908 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8620
timestamp 1682952543
transform 1 0 2932 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8421
timestamp 1682952543
transform 1 0 2932 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8656
timestamp 1682952543
transform 1 0 2940 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8422
timestamp 1682952543
transform 1 0 2948 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8546
timestamp 1682952543
transform 1 0 2940 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8681
timestamp 1682952543
transform 1 0 2948 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8547
timestamp 1682952543
transform 1 0 2956 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8716
timestamp 1682952543
transform 1 0 2948 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8515
timestamp 1682952543
transform 1 0 2996 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_8526
timestamp 1682952543
transform 1 0 3004 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8547
timestamp 1682952543
transform 1 0 2996 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8621
timestamp 1682952543
transform 1 0 2988 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8622
timestamp 1682952543
transform 1 0 3004 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8423
timestamp 1682952543
transform 1 0 2996 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8424
timestamp 1682952543
transform 1 0 3020 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8548
timestamp 1682952543
transform 1 0 2988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8549
timestamp 1682952543
transform 1 0 3004 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8745
timestamp 1682952543
transform 1 0 2988 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8548
timestamp 1682952543
transform 1 0 3044 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8657
timestamp 1682952543
transform 1 0 3036 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8425
timestamp 1682952543
transform 1 0 3044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8550
timestamp 1682952543
transform 1 0 3036 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8527
timestamp 1682952543
transform 1 0 3060 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8746
timestamp 1682952543
transform 1 0 3052 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8623
timestamp 1682952543
transform 1 0 3100 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8426
timestamp 1682952543
transform 1 0 3100 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8551
timestamp 1682952543
transform 1 0 3148 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8528
timestamp 1682952543
transform 1 0 3260 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8549
timestamp 1682952543
transform 1 0 3252 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8569
timestamp 1682952543
transform 1 0 3172 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8570
timestamp 1682952543
transform 1 0 3212 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8571
timestamp 1682952543
transform 1 0 3244 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8624
timestamp 1682952543
transform 1 0 3212 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8427
timestamp 1682952543
transform 1 0 3212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8552
timestamp 1682952543
transform 1 0 3172 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8717
timestamp 1682952543
transform 1 0 3220 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8718
timestamp 1682952543
transform 1 0 3236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8625
timestamp 1682952543
transform 1 0 3292 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8428
timestamp 1682952543
transform 1 0 3268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8429
timestamp 1682952543
transform 1 0 3276 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8658
timestamp 1682952543
transform 1 0 3284 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8430
timestamp 1682952543
transform 1 0 3300 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8682
timestamp 1682952543
transform 1 0 3268 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8553
timestamp 1682952543
transform 1 0 3276 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8554
timestamp 1682952543
transform 1 0 3292 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8683
timestamp 1682952543
transform 1 0 3300 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8719
timestamp 1682952543
transform 1 0 3276 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8555
timestamp 1682952543
transform 1 0 3316 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8572
timestamp 1682952543
transform 1 0 3324 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8659
timestamp 1682952543
transform 1 0 3324 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8431
timestamp 1682952543
transform 1 0 3332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8556
timestamp 1682952543
transform 1 0 3332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8626
timestamp 1682952543
transform 1 0 3364 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8660
timestamp 1682952543
transform 1 0 3372 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8573
timestamp 1682952543
transform 1 0 3388 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8432
timestamp 1682952543
transform 1 0 3380 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8433
timestamp 1682952543
transform 1 0 3404 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8627
timestamp 1682952543
transform 1 0 3420 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8557
timestamp 1682952543
transform 1 0 3372 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8558
timestamp 1682952543
transform 1 0 3380 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8559
timestamp 1682952543
transform 1 0 3396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8560
timestamp 1682952543
transform 1 0 3412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8561
timestamp 1682952543
transform 1 0 3420 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8720
timestamp 1682952543
transform 1 0 3380 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8721
timestamp 1682952543
transform 1 0 3412 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8661
timestamp 1682952543
transform 1 0 3428 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8529
timestamp 1682952543
transform 1 0 3468 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8574
timestamp 1682952543
transform 1 0 3444 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8575
timestamp 1682952543
transform 1 0 3476 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8628
timestamp 1682952543
transform 1 0 3460 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8629
timestamp 1682952543
transform 1 0 3500 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8630
timestamp 1682952543
transform 1 0 3516 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8434
timestamp 1682952543
transform 1 0 3436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8435
timestamp 1682952543
transform 1 0 3452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8436
timestamp 1682952543
transform 1 0 3468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8437
timestamp 1682952543
transform 1 0 3484 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8662
timestamp 1682952543
transform 1 0 3492 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8438
timestamp 1682952543
transform 1 0 3500 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8439
timestamp 1682952543
transform 1 0 3516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8562
timestamp 1682952543
transform 1 0 3444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8563
timestamp 1682952543
transform 1 0 3460 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8684
timestamp 1682952543
transform 1 0 3468 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8564
timestamp 1682952543
transform 1 0 3476 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8685
timestamp 1682952543
transform 1 0 3484 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8565
timestamp 1682952543
transform 1 0 3492 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8566
timestamp 1682952543
transform 1 0 3508 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8747
timestamp 1682952543
transform 1 0 3444 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8748
timestamp 1682952543
transform 1 0 3476 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8440
timestamp 1682952543
transform 1 0 3588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8567
timestamp 1682952543
transform 1 0 3524 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8568
timestamp 1682952543
transform 1 0 3540 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8722
timestamp 1682952543
transform 1 0 3588 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8530
timestamp 1682952543
transform 1 0 3652 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_8631
timestamp 1682952543
transform 1 0 3660 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8632
timestamp 1682952543
transform 1 0 3684 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8441
timestamp 1682952543
transform 1 0 3660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8442
timestamp 1682952543
transform 1 0 3668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8443
timestamp 1682952543
transform 1 0 3684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8569
timestamp 1682952543
transform 1 0 3660 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8570
timestamp 1682952543
transform 1 0 3676 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8686
timestamp 1682952543
transform 1 0 3684 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8633
timestamp 1682952543
transform 1 0 3716 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8444
timestamp 1682952543
transform 1 0 3708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8571
timestamp 1682952543
transform 1 0 3692 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8723
timestamp 1682952543
transform 1 0 3676 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8687
timestamp 1682952543
transform 1 0 3700 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_8749
timestamp 1682952543
transform 1 0 3692 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8572
timestamp 1682952543
transform 1 0 3716 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8724
timestamp 1682952543
transform 1 0 3708 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8531
timestamp 1682952543
transform 1 0 3756 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8445
timestamp 1682952543
transform 1 0 3740 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8663
timestamp 1682952543
transform 1 0 3748 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8576
timestamp 1682952543
transform 1 0 3764 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8321
timestamp 1682952543
transform 1 0 3780 0 1 635
box -2 -2 2 2
use M2_M1  M2_M1_8446
timestamp 1682952543
transform 1 0 3756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8573
timestamp 1682952543
transform 1 0 3748 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8725
timestamp 1682952543
transform 1 0 3732 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8329
timestamp 1682952543
transform 1 0 3772 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_8634
timestamp 1682952543
transform 1 0 3788 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8330
timestamp 1682952543
transform 1 0 3796 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8447
timestamp 1682952543
transform 1 0 3788 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8664
timestamp 1682952543
transform 1 0 3796 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_8550
timestamp 1682952543
transform 1 0 3844 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_8635
timestamp 1682952543
transform 1 0 3828 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8448
timestamp 1682952543
transform 1 0 3812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8449
timestamp 1682952543
transform 1 0 3828 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8665
timestamp 1682952543
transform 1 0 3836 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8450
timestamp 1682952543
transform 1 0 3844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8451
timestamp 1682952543
transform 1 0 3852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8574
timestamp 1682952543
transform 1 0 3820 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8575
timestamp 1682952543
transform 1 0 3836 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8577
timestamp 1682952543
transform 1 0 3900 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8578
timestamp 1682952543
transform 1 0 3948 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8579
timestamp 1682952543
transform 1 0 3964 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8580
timestamp 1682952543
transform 1 0 3988 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_8636
timestamp 1682952543
transform 1 0 3884 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_8637
timestamp 1682952543
transform 1 0 3940 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8452
timestamp 1682952543
transform 1 0 3876 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8453
timestamp 1682952543
transform 1 0 3892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8454
timestamp 1682952543
transform 1 0 3908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8455
timestamp 1682952543
transform 1 0 3940 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8456
timestamp 1682952543
transform 1 0 4012 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_8666
timestamp 1682952543
transform 1 0 4020 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8457
timestamp 1682952543
transform 1 0 4028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8458
timestamp 1682952543
transform 1 0 4076 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8576
timestamp 1682952543
transform 1 0 3860 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8577
timestamp 1682952543
transform 1 0 3868 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8578
timestamp 1682952543
transform 1 0 3884 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8579
timestamp 1682952543
transform 1 0 3900 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8580
timestamp 1682952543
transform 1 0 3988 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8581
timestamp 1682952543
transform 1 0 4004 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8582
timestamp 1682952543
transform 1 0 4020 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8583
timestamp 1682952543
transform 1 0 4036 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8584
timestamp 1682952543
transform 1 0 4052 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_8726
timestamp 1682952543
transform 1 0 3860 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8750
timestamp 1682952543
transform 1 0 3820 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8751
timestamp 1682952543
transform 1 0 3852 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8727
timestamp 1682952543
transform 1 0 3908 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8752
timestamp 1682952543
transform 1 0 3876 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8753
timestamp 1682952543
transform 1 0 3900 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8728
timestamp 1682952543
transform 1 0 4020 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8754
timestamp 1682952543
transform 1 0 4004 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_8729
timestamp 1682952543
transform 1 0 4076 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_8638
timestamp 1682952543
transform 1 0 4148 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8459
timestamp 1682952543
transform 1 0 4148 0 1 615
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_70
timestamp 1682952543
transform 1 0 48 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_8755
timestamp 1682952543
transform 1 0 84 0 1 575
box -3 -3 3 3
use FILL  FILL_3710
timestamp 1682952543
transform 1 0 72 0 1 570
box -8 -3 16 105
use FILL  FILL_3711
timestamp 1682952543
transform 1 0 80 0 1 570
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1682952543
transform 1 0 88 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8756
timestamp 1682952543
transform 1 0 108 0 1 575
box -3 -3 3 3
use FILL  FILL_3713
timestamp 1682952543
transform 1 0 96 0 1 570
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1682952543
transform 1 0 104 0 1 570
box -8 -3 16 105
use FILL  FILL_3715
timestamp 1682952543
transform 1 0 112 0 1 570
box -8 -3 16 105
use INVX2  INVX2_597
timestamp 1682952543
transform -1 0 136 0 1 570
box -9 -3 26 105
use FILL  FILL_3716
timestamp 1682952543
transform 1 0 136 0 1 570
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1682952543
transform 1 0 144 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_347
timestamp 1682952543
transform -1 0 192 0 1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_531
timestamp 1682952543
transform 1 0 192 0 1 570
box -8 -3 104 105
use INVX2  INVX2_598
timestamp 1682952543
transform -1 0 304 0 1 570
box -9 -3 26 105
use FILL  FILL_3718
timestamp 1682952543
transform 1 0 304 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_348
timestamp 1682952543
transform 1 0 312 0 1 570
box -8 -3 46 105
use FILL  FILL_3719
timestamp 1682952543
transform 1 0 352 0 1 570
box -8 -3 16 105
use INVX2  INVX2_599
timestamp 1682952543
transform 1 0 360 0 1 570
box -9 -3 26 105
use FILL  FILL_3720
timestamp 1682952543
transform 1 0 376 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8757
timestamp 1682952543
transform 1 0 396 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_532
timestamp 1682952543
transform 1 0 384 0 1 570
box -8 -3 104 105
use INVX2  INVX2_600
timestamp 1682952543
transform 1 0 480 0 1 570
box -9 -3 26 105
use FILL  FILL_3721
timestamp 1682952543
transform 1 0 496 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8758
timestamp 1682952543
transform 1 0 524 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_377
timestamp 1682952543
transform 1 0 504 0 1 570
box -8 -3 46 105
use FILL  FILL_3722
timestamp 1682952543
transform 1 0 544 0 1 570
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1682952543
transform 1 0 552 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_378
timestamp 1682952543
transform -1 0 600 0 1 570
box -8 -3 46 105
use INVX2  INVX2_601
timestamp 1682952543
transform 1 0 600 0 1 570
box -9 -3 26 105
use FILL  FILL_3724
timestamp 1682952543
transform 1 0 616 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_533
timestamp 1682952543
transform -1 0 720 0 1 570
box -8 -3 104 105
use FILL  FILL_3725
timestamp 1682952543
transform 1 0 720 0 1 570
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1682952543
transform 1 0 728 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_349
timestamp 1682952543
transform 1 0 736 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_8759
timestamp 1682952543
transform 1 0 796 0 1 575
box -3 -3 3 3
use INVX2  INVX2_602
timestamp 1682952543
transform 1 0 776 0 1 570
box -9 -3 26 105
use FILL  FILL_3727
timestamp 1682952543
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_3728
timestamp 1682952543
transform 1 0 800 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_100
timestamp 1682952543
transform 1 0 808 0 1 570
box -8 -3 32 105
use M3_M2  M3_M2_8760
timestamp 1682952543
transform 1 0 860 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_149
timestamp 1682952543
transform 1 0 832 0 1 570
box -8 -3 34 105
use FILL  FILL_3729
timestamp 1682952543
transform 1 0 864 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_101
timestamp 1682952543
transform 1 0 872 0 1 570
box -8 -3 32 105
use INVX2  INVX2_603
timestamp 1682952543
transform 1 0 896 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_534
timestamp 1682952543
transform -1 0 1008 0 1 570
box -8 -3 104 105
use FILL  FILL_3730
timestamp 1682952543
transform 1 0 1008 0 1 570
box -8 -3 16 105
use FILL  FILL_3731
timestamp 1682952543
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1682952543
transform 1 0 1024 0 1 570
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1682952543
transform 1 0 1032 0 1 570
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1682952543
transform 1 0 1040 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_150
timestamp 1682952543
transform -1 0 1080 0 1 570
box -8 -3 34 105
use FILL  FILL_3735
timestamp 1682952543
transform 1 0 1080 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_535
timestamp 1682952543
transform -1 0 1184 0 1 570
box -8 -3 104 105
use FILL  FILL_3736
timestamp 1682952543
transform 1 0 1184 0 1 570
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1682952543
transform 1 0 1192 0 1 570
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1682952543
transform 1 0 1200 0 1 570
box -8 -3 16 105
use INVX2  INVX2_604
timestamp 1682952543
transform 1 0 1208 0 1 570
box -9 -3 26 105
use FILL  FILL_3739
timestamp 1682952543
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1682952543
transform 1 0 1232 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_536
timestamp 1682952543
transform 1 0 1240 0 1 570
box -8 -3 104 105
use INVX2  INVX2_605
timestamp 1682952543
transform 1 0 1336 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_8761
timestamp 1682952543
transform 1 0 1380 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_379
timestamp 1682952543
transform -1 0 1392 0 1 570
box -8 -3 46 105
use INVX2  INVX2_606
timestamp 1682952543
transform -1 0 1408 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_537
timestamp 1682952543
transform 1 0 1408 0 1 570
box -8 -3 104 105
use INVX2  INVX2_607
timestamp 1682952543
transform -1 0 1520 0 1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_350
timestamp 1682952543
transform 1 0 1520 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_380
timestamp 1682952543
transform 1 0 1560 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_8762
timestamp 1682952543
transform 1 0 1628 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_381
timestamp 1682952543
transform 1 0 1600 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_8763
timestamp 1682952543
transform 1 0 1668 0 1 575
box -3 -3 3 3
use INVX2  INVX2_608
timestamp 1682952543
transform 1 0 1640 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_8764
timestamp 1682952543
transform 1 0 1740 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_538
timestamp 1682952543
transform -1 0 1752 0 1 570
box -8 -3 104 105
use M3_M2  M3_M2_8765
timestamp 1682952543
transform 1 0 1780 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_8766
timestamp 1682952543
transform 1 0 1796 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_539
timestamp 1682952543
transform 1 0 1752 0 1 570
box -8 -3 104 105
use FILL  FILL_3741
timestamp 1682952543
transform 1 0 1848 0 1 570
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1682952543
transform 1 0 1856 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_151
timestamp 1682952543
transform 1 0 1864 0 1 570
box -8 -3 34 105
use FILL  FILL_3743
timestamp 1682952543
transform 1 0 1896 0 1 570
box -8 -3 16 105
use FILL  FILL_3744
timestamp 1682952543
transform 1 0 1904 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_103
timestamp 1682952543
transform 1 0 1912 0 1 570
box -8 -3 32 105
use FILL  FILL_3776
timestamp 1682952543
transform 1 0 1936 0 1 570
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1682952543
transform 1 0 1944 0 1 570
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1682952543
transform 1 0 1952 0 1 570
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1682952543
transform 1 0 1960 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_158
timestamp 1682952543
transform -1 0 2000 0 1 570
box -8 -3 34 105
use FILL  FILL_3780
timestamp 1682952543
transform 1 0 2000 0 1 570
box -8 -3 16 105
use INVX2  INVX2_617
timestamp 1682952543
transform 1 0 2008 0 1 570
box -9 -3 26 105
use FILL  FILL_3781
timestamp 1682952543
transform 1 0 2024 0 1 570
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1682952543
transform 1 0 2032 0 1 570
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1682952543
transform 1 0 2040 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_386
timestamp 1682952543
transform -1 0 2088 0 1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_548
timestamp 1682952543
transform -1 0 2184 0 1 570
box -8 -3 104 105
use INVX2  INVX2_618
timestamp 1682952543
transform 1 0 2184 0 1 570
box -9 -3 26 105
use FILL  FILL_3784
timestamp 1682952543
transform 1 0 2200 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_387
timestamp 1682952543
transform 1 0 2208 0 1 570
box -8 -3 46 105
use INVX2  INVX2_619
timestamp 1682952543
transform 1 0 2248 0 1 570
box -9 -3 26 105
use FILL  FILL_3785
timestamp 1682952543
transform 1 0 2264 0 1 570
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1682952543
transform 1 0 2272 0 1 570
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1682952543
transform 1 0 2280 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8767
timestamp 1682952543
transform 1 0 2316 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_159
timestamp 1682952543
transform 1 0 2288 0 1 570
box -8 -3 34 105
use FILL  FILL_3788
timestamp 1682952543
transform 1 0 2320 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_160
timestamp 1682952543
transform 1 0 2328 0 1 570
box -8 -3 34 105
use FILL  FILL_3789
timestamp 1682952543
transform 1 0 2360 0 1 570
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1682952543
transform 1 0 2368 0 1 570
box -8 -3 16 105
use INVX2  INVX2_620
timestamp 1682952543
transform 1 0 2376 0 1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_359
timestamp 1682952543
transform 1 0 2392 0 1 570
box -8 -3 46 105
use FILL  FILL_3791
timestamp 1682952543
transform 1 0 2432 0 1 570
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1682952543
transform 1 0 2440 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8768
timestamp 1682952543
transform 1 0 2476 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_161
timestamp 1682952543
transform 1 0 2448 0 1 570
box -8 -3 34 105
use FILL  FILL_3793
timestamp 1682952543
transform 1 0 2480 0 1 570
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1682952543
transform 1 0 2488 0 1 570
box -8 -3 16 105
use FILL  FILL_3796
timestamp 1682952543
transform 1 0 2496 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_389
timestamp 1682952543
transform 1 0 2504 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_360
timestamp 1682952543
transform -1 0 2584 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_361
timestamp 1682952543
transform 1 0 2584 0 1 570
box -8 -3 46 105
use INVX2  INVX2_623
timestamp 1682952543
transform 1 0 2624 0 1 570
box -9 -3 26 105
use BUFX2  BUFX2_102
timestamp 1682952543
transform -1 0 2664 0 1 570
box -5 -3 28 105
use BUFX2  BUFX2_103
timestamp 1682952543
transform 1 0 2664 0 1 570
box -5 -3 28 105
use BUFX2  BUFX2_104
timestamp 1682952543
transform 1 0 2688 0 1 570
box -5 -3 28 105
use M3_M2  M3_M2_8769
timestamp 1682952543
transform 1 0 2748 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_553
timestamp 1682952543
transform 1 0 2712 0 1 570
box -8 -3 104 105
use INVX2  INVX2_625
timestamp 1682952543
transform 1 0 2808 0 1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_391
timestamp 1682952543
transform -1 0 2864 0 1 570
box -8 -3 46 105
use FILL  FILL_3806
timestamp 1682952543
transform 1 0 2864 0 1 570
box -8 -3 16 105
use FILL  FILL_3807
timestamp 1682952543
transform 1 0 2872 0 1 570
box -8 -3 16 105
use FILL  FILL_3808
timestamp 1682952543
transform 1 0 2880 0 1 570
box -8 -3 16 105
use INVX2  INVX2_626
timestamp 1682952543
transform 1 0 2888 0 1 570
box -9 -3 26 105
use FILL  FILL_3809
timestamp 1682952543
transform 1 0 2904 0 1 570
box -8 -3 16 105
use FILL  FILL_3810
timestamp 1682952543
transform 1 0 2912 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_392
timestamp 1682952543
transform -1 0 2960 0 1 570
box -8 -3 46 105
use FILL  FILL_3811
timestamp 1682952543
transform 1 0 2960 0 1 570
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1682952543
transform 1 0 2968 0 1 570
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1682952543
transform 1 0 2976 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_393
timestamp 1682952543
transform -1 0 3024 0 1 570
box -8 -3 46 105
use FILL  FILL_3814
timestamp 1682952543
transform 1 0 3024 0 1 570
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1682952543
transform 1 0 3032 0 1 570
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1682952543
transform 1 0 3040 0 1 570
box -8 -3 16 105
use INVX2  INVX2_627
timestamp 1682952543
transform -1 0 3064 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_554
timestamp 1682952543
transform -1 0 3160 0 1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_555
timestamp 1682952543
transform 1 0 3160 0 1 570
box -8 -3 104 105
use INVX2  INVX2_628
timestamp 1682952543
transform 1 0 3256 0 1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_394
timestamp 1682952543
transform 1 0 3272 0 1 570
box -8 -3 46 105
use FILL  FILL_3817
timestamp 1682952543
transform 1 0 3312 0 1 570
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1682952543
transform 1 0 3320 0 1 570
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1682952543
transform 1 0 3328 0 1 570
box -8 -3 16 105
use INVX2  INVX2_629
timestamp 1682952543
transform -1 0 3352 0 1 570
box -9 -3 26 105
use FILL  FILL_3820
timestamp 1682952543
transform 1 0 3352 0 1 570
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1682952543
transform 1 0 3360 0 1 570
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1682952543
transform 1 0 3368 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_396
timestamp 1682952543
transform 1 0 3376 0 1 570
box -8 -3 46 105
use FILL  FILL_3841
timestamp 1682952543
transform 1 0 3416 0 1 570
box -8 -3 16 105
use FILL  FILL_3842
timestamp 1682952543
transform 1 0 3424 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_363
timestamp 1682952543
transform 1 0 3432 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_397
timestamp 1682952543
transform 1 0 3472 0 1 570
box -8 -3 46 105
use INVX2  INVX2_634
timestamp 1682952543
transform -1 0 3528 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_558
timestamp 1682952543
transform 1 0 3528 0 1 570
box -8 -3 104 105
use INVX2  INVX2_635
timestamp 1682952543
transform 1 0 3624 0 1 570
box -9 -3 26 105
use FILL  FILL_3843
timestamp 1682952543
transform 1 0 3640 0 1 570
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1682952543
transform 1 0 3648 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_398
timestamp 1682952543
transform 1 0 3656 0 1 570
box -8 -3 46 105
use FILL  FILL_3845
timestamp 1682952543
transform 1 0 3696 0 1 570
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1682952543
transform 1 0 3704 0 1 570
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1682952543
transform 1 0 3712 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_8770
timestamp 1682952543
transform 1 0 3780 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_364
timestamp 1682952543
transform 1 0 3720 0 1 570
box -8 -3 46 105
use FILL  FILL_3848
timestamp 1682952543
transform 1 0 3760 0 1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_71
timestamp 1682952543
transform -1 0 3800 0 1 570
box -8 -3 40 105
use FILL  FILL_3849
timestamp 1682952543
transform 1 0 3800 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_365
timestamp 1682952543
transform 1 0 3808 0 1 570
box -8 -3 46 105
use INVX2  INVX2_636
timestamp 1682952543
transform -1 0 3864 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_8771
timestamp 1682952543
transform 1 0 3884 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_399
timestamp 1682952543
transform -1 0 3904 0 1 570
box -8 -3 46 105
use M3_M2  M3_M2_8772
timestamp 1682952543
transform 1 0 3924 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_559
timestamp 1682952543
transform -1 0 4000 0 1 570
box -8 -3 104 105
use OAI22X1  OAI22X1_400
timestamp 1682952543
transform 1 0 4000 0 1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_560
timestamp 1682952543
transform 1 0 4040 0 1 570
box -8 -3 104 105
use INVX2  INVX2_637
timestamp 1682952543
transform 1 0 4136 0 1 570
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_71
timestamp 1682952543
transform 1 0 4177 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_8773
timestamp 1682952543
transform 1 0 172 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8825
timestamp 1682952543
transform 1 0 164 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8826
timestamp 1682952543
transform 1 0 180 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8774
timestamp 1682952543
transform 1 0 220 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8593
timestamp 1682952543
transform 1 0 84 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8594
timestamp 1682952543
transform 1 0 172 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8595
timestamp 1682952543
transform 1 0 180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8596
timestamp 1682952543
transform 1 0 196 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8858
timestamp 1682952543
transform 1 0 204 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8597
timestamp 1682952543
transform 1 0 212 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8827
timestamp 1682952543
transform 1 0 228 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8598
timestamp 1682952543
transform 1 0 228 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8859
timestamp 1682952543
transform 1 0 236 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8701
timestamp 1682952543
transform 1 0 132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8702
timestamp 1682952543
transform 1 0 164 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8703
timestamp 1682952543
transform 1 0 188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8704
timestamp 1682952543
transform 1 0 204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8705
timestamp 1682952543
transform 1 0 220 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8918
timestamp 1682952543
transform 1 0 132 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8919
timestamp 1682952543
transform 1 0 172 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8920
timestamp 1682952543
transform 1 0 204 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8775
timestamp 1682952543
transform 1 0 268 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8599
timestamp 1682952543
transform 1 0 260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8706
timestamp 1682952543
transform 1 0 252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8707
timestamp 1682952543
transform 1 0 276 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8860
timestamp 1682952543
transform 1 0 308 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8796
timestamp 1682952543
transform 1 0 340 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8797
timestamp 1682952543
transform 1 0 356 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8600
timestamp 1682952543
transform 1 0 316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8601
timestamp 1682952543
transform 1 0 340 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8861
timestamp 1682952543
transform 1 0 348 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8708
timestamp 1682952543
transform 1 0 308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8709
timestamp 1682952543
transform 1 0 324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8710
timestamp 1682952543
transform 1 0 340 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8921
timestamp 1682952543
transform 1 0 340 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8798
timestamp 1682952543
transform 1 0 444 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8602
timestamp 1682952543
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8711
timestamp 1682952543
transform 1 0 412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8712
timestamp 1682952543
transform 1 0 444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8713
timestamp 1682952543
transform 1 0 452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8714
timestamp 1682952543
transform 1 0 460 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8922
timestamp 1682952543
transform 1 0 412 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8923
timestamp 1682952543
transform 1 0 452 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8799
timestamp 1682952543
transform 1 0 500 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8603
timestamp 1682952543
transform 1 0 476 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8604
timestamp 1682952543
transform 1 0 484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8605
timestamp 1682952543
transform 1 0 500 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8606
timestamp 1682952543
transform 1 0 516 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8715
timestamp 1682952543
transform 1 0 476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8716
timestamp 1682952543
transform 1 0 492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8717
timestamp 1682952543
transform 1 0 508 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8924
timestamp 1682952543
transform 1 0 476 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8800
timestamp 1682952543
transform 1 0 548 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8607
timestamp 1682952543
transform 1 0 548 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8718
timestamp 1682952543
transform 1 0 540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8719
timestamp 1682952543
transform 1 0 556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8720
timestamp 1682952543
transform 1 0 564 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8980
timestamp 1682952543
transform 1 0 548 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_8608
timestamp 1682952543
transform 1 0 580 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8828
timestamp 1682952543
transform 1 0 604 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8862
timestamp 1682952543
transform 1 0 596 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8609
timestamp 1682952543
transform 1 0 620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8610
timestamp 1682952543
transform 1 0 628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8721
timestamp 1682952543
transform 1 0 596 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8722
timestamp 1682952543
transform 1 0 612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8889
timestamp 1682952543
transform 1 0 620 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8723
timestamp 1682952543
transform 1 0 628 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8925
timestamp 1682952543
transform 1 0 596 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8801
timestamp 1682952543
transform 1 0 708 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8802
timestamp 1682952543
transform 1 0 740 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8611
timestamp 1682952543
transform 1 0 740 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8724
timestamp 1682952543
transform 1 0 652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8725
timestamp 1682952543
transform 1 0 660 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8890
timestamp 1682952543
transform 1 0 668 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8726
timestamp 1682952543
transform 1 0 692 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8926
timestamp 1682952543
transform 1 0 652 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8927
timestamp 1682952543
transform 1 0 692 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8981
timestamp 1682952543
transform 1 0 708 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8982
timestamp 1682952543
transform 1 0 732 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8829
timestamp 1682952543
transform 1 0 812 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8612
timestamp 1682952543
transform 1 0 764 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8727
timestamp 1682952543
transform 1 0 788 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8728
timestamp 1682952543
transform 1 0 844 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8957
timestamp 1682952543
transform 1 0 836 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8971
timestamp 1682952543
transform 1 0 836 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8803
timestamp 1682952543
transform 1 0 860 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8804
timestamp 1682952543
transform 1 0 892 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8830
timestamp 1682952543
transform 1 0 868 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8613
timestamp 1682952543
transform 1 0 860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8614
timestamp 1682952543
transform 1 0 868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8615
timestamp 1682952543
transform 1 0 892 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8616
timestamp 1682952543
transform 1 0 900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8729
timestamp 1682952543
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8730
timestamp 1682952543
transform 1 0 892 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8928
timestamp 1682952543
transform 1 0 876 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8617
timestamp 1682952543
transform 1 0 924 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8776
timestamp 1682952543
transform 1 0 956 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8805
timestamp 1682952543
transform 1 0 948 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8618
timestamp 1682952543
transform 1 0 948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8731
timestamp 1682952543
transform 1 0 924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8732
timestamp 1682952543
transform 1 0 932 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8929
timestamp 1682952543
transform 1 0 900 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8930
timestamp 1682952543
transform 1 0 932 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8589
timestamp 1682952543
transform 1 0 956 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_8891
timestamp 1682952543
transform 1 0 956 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8619
timestamp 1682952543
transform 1 0 972 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8931
timestamp 1682952543
transform 1 0 964 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8824
timestamp 1682952543
transform 1 0 972 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8958
timestamp 1682952543
transform 1 0 972 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8777
timestamp 1682952543
transform 1 0 988 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8863
timestamp 1682952543
transform 1 0 1004 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8778
timestamp 1682952543
transform 1 0 1044 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8620
timestamp 1682952543
transform 1 0 1012 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8892
timestamp 1682952543
transform 1 0 996 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8733
timestamp 1682952543
transform 1 0 1004 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8959
timestamp 1682952543
transform 1 0 988 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8864
timestamp 1682952543
transform 1 0 1028 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8621
timestamp 1682952543
transform 1 0 1036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8622
timestamp 1682952543
transform 1 0 1044 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8865
timestamp 1682952543
transform 1 0 1060 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8623
timestamp 1682952543
transform 1 0 1068 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8624
timestamp 1682952543
transform 1 0 1076 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8734
timestamp 1682952543
transform 1 0 1020 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8893
timestamp 1682952543
transform 1 0 1036 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8735
timestamp 1682952543
transform 1 0 1060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8825
timestamp 1682952543
transform 1 0 1036 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8866
timestamp 1682952543
transform 1 0 1092 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8625
timestamp 1682952543
transform 1 0 1100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8626
timestamp 1682952543
transform 1 0 1108 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8736
timestamp 1682952543
transform 1 0 1092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8826
timestamp 1682952543
transform 1 0 1044 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8932
timestamp 1682952543
transform 1 0 1068 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8827
timestamp 1682952543
transform 1 0 1076 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8960
timestamp 1682952543
transform 1 0 1044 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8961
timestamp 1682952543
transform 1 0 1076 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8894
timestamp 1682952543
transform 1 0 1108 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8831
timestamp 1682952543
transform 1 0 1220 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8627
timestamp 1682952543
transform 1 0 1132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8628
timestamp 1682952543
transform 1 0 1220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8737
timestamp 1682952543
transform 1 0 1124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8738
timestamp 1682952543
transform 1 0 1140 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8739
timestamp 1682952543
transform 1 0 1196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8828
timestamp 1682952543
transform 1 0 1108 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8962
timestamp 1682952543
transform 1 0 1108 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8983
timestamp 1682952543
transform 1 0 1084 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8963
timestamp 1682952543
transform 1 0 1132 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8832
timestamp 1682952543
transform 1 0 1244 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8629
timestamp 1682952543
transform 1 0 1244 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8867
timestamp 1682952543
transform 1 0 1292 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8740
timestamp 1682952543
transform 1 0 1292 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8964
timestamp 1682952543
transform 1 0 1228 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8630
timestamp 1682952543
transform 1 0 1348 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8868
timestamp 1682952543
transform 1 0 1356 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8631
timestamp 1682952543
transform 1 0 1364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8632
timestamp 1682952543
transform 1 0 1380 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8741
timestamp 1682952543
transform 1 0 1340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8742
timestamp 1682952543
transform 1 0 1356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8743
timestamp 1682952543
transform 1 0 1372 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8933
timestamp 1682952543
transform 1 0 1340 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8779
timestamp 1682952543
transform 1 0 1404 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8780
timestamp 1682952543
transform 1 0 1508 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8633
timestamp 1682952543
transform 1 0 1412 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8869
timestamp 1682952543
transform 1 0 1492 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8895
timestamp 1682952543
transform 1 0 1412 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8896
timestamp 1682952543
transform 1 0 1452 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8744
timestamp 1682952543
transform 1 0 1460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8745
timestamp 1682952543
transform 1 0 1492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8746
timestamp 1682952543
transform 1 0 1500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8747
timestamp 1682952543
transform 1 0 1508 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8934
timestamp 1682952543
transform 1 0 1460 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8935
timestamp 1682952543
transform 1 0 1500 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8984
timestamp 1682952543
transform 1 0 1436 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8897
timestamp 1682952543
transform 1 0 1516 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8833
timestamp 1682952543
transform 1 0 1556 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8834
timestamp 1682952543
transform 1 0 1604 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8634
timestamp 1682952543
transform 1 0 1532 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8635
timestamp 1682952543
transform 1 0 1540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8636
timestamp 1682952543
transform 1 0 1556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8637
timestamp 1682952543
transform 1 0 1572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8638
timestamp 1682952543
transform 1 0 1588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8748
timestamp 1682952543
transform 1 0 1548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8749
timestamp 1682952543
transform 1 0 1564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8750
timestamp 1682952543
transform 1 0 1580 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8751
timestamp 1682952543
transform 1 0 1596 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8898
timestamp 1682952543
transform 1 0 1604 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8752
timestamp 1682952543
transform 1 0 1612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8936
timestamp 1682952543
transform 1 0 1596 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8781
timestamp 1682952543
transform 1 0 1620 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8639
timestamp 1682952543
transform 1 0 1620 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8640
timestamp 1682952543
transform 1 0 1644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8641
timestamp 1682952543
transform 1 0 1660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8642
timestamp 1682952543
transform 1 0 1668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8753
timestamp 1682952543
transform 1 0 1636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8754
timestamp 1682952543
transform 1 0 1652 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8937
timestamp 1682952543
transform 1 0 1644 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8965
timestamp 1682952543
transform 1 0 1636 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8755
timestamp 1682952543
transform 1 0 1676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8756
timestamp 1682952543
transform 1 0 1700 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8806
timestamp 1682952543
transform 1 0 1724 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8643
timestamp 1682952543
transform 1 0 1724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8757
timestamp 1682952543
transform 1 0 1724 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8938
timestamp 1682952543
transform 1 0 1724 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8807
timestamp 1682952543
transform 1 0 1844 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8835
timestamp 1682952543
transform 1 0 1740 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8836
timestamp 1682952543
transform 1 0 1764 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8837
timestamp 1682952543
transform 1 0 1820 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8644
timestamp 1682952543
transform 1 0 1740 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8870
timestamp 1682952543
transform 1 0 1772 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8899
timestamp 1682952543
transform 1 0 1740 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8758
timestamp 1682952543
transform 1 0 1764 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8900
timestamp 1682952543
transform 1 0 1780 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8838
timestamp 1682952543
transform 1 0 1860 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8645
timestamp 1682952543
transform 1 0 1836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8646
timestamp 1682952543
transform 1 0 1860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8759
timestamp 1682952543
transform 1 0 1820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8760
timestamp 1682952543
transform 1 0 1828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8761
timestamp 1682952543
transform 1 0 1844 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8939
timestamp 1682952543
transform 1 0 1764 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8966
timestamp 1682952543
transform 1 0 1828 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8762
timestamp 1682952543
transform 1 0 1868 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8763
timestamp 1682952543
transform 1 0 1876 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8782
timestamp 1682952543
transform 1 0 1908 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8590
timestamp 1682952543
transform 1 0 1908 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8647
timestamp 1682952543
transform 1 0 1916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8648
timestamp 1682952543
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8649
timestamp 1682952543
transform 1 0 1940 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8901
timestamp 1682952543
transform 1 0 1908 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8764
timestamp 1682952543
transform 1 0 1932 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8829
timestamp 1682952543
transform 1 0 1908 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8902
timestamp 1682952543
transform 1 0 1940 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8839
timestamp 1682952543
transform 1 0 2052 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8650
timestamp 1682952543
transform 1 0 1964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8651
timestamp 1682952543
transform 1 0 2052 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8765
timestamp 1682952543
transform 1 0 1956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8766
timestamp 1682952543
transform 1 0 1972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8767
timestamp 1682952543
transform 1 0 2012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8830
timestamp 1682952543
transform 1 0 1940 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8940
timestamp 1682952543
transform 1 0 1964 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8967
timestamp 1682952543
transform 1 0 1948 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8972
timestamp 1682952543
transform 1 0 1924 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8973
timestamp 1682952543
transform 1 0 1940 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8840
timestamp 1682952543
transform 1 0 2076 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8841
timestamp 1682952543
transform 1 0 2108 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8652
timestamp 1682952543
transform 1 0 2076 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8768
timestamp 1682952543
transform 1 0 2124 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8941
timestamp 1682952543
transform 1 0 2116 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8974
timestamp 1682952543
transform 1 0 1980 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8975
timestamp 1682952543
transform 1 0 2028 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8976
timestamp 1682952543
transform 1 0 2068 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8842
timestamp 1682952543
transform 1 0 2172 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8653
timestamp 1682952543
transform 1 0 2180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8769
timestamp 1682952543
transform 1 0 2172 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8942
timestamp 1682952543
transform 1 0 2172 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8808
timestamp 1682952543
transform 1 0 2212 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8809
timestamp 1682952543
transform 1 0 2300 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8843
timestamp 1682952543
transform 1 0 2212 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8654
timestamp 1682952543
transform 1 0 2212 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8770
timestamp 1682952543
transform 1 0 2196 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8771
timestamp 1682952543
transform 1 0 2236 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8943
timestamp 1682952543
transform 1 0 2196 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8783
timestamp 1682952543
transform 1 0 2364 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8810
timestamp 1682952543
transform 1 0 2356 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8811
timestamp 1682952543
transform 1 0 2396 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8655
timestamp 1682952543
transform 1 0 2316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8656
timestamp 1682952543
transform 1 0 2332 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8871
timestamp 1682952543
transform 1 0 2340 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8844
timestamp 1682952543
transform 1 0 2364 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8657
timestamp 1682952543
transform 1 0 2348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8658
timestamp 1682952543
transform 1 0 2364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8772
timestamp 1682952543
transform 1 0 2308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8773
timestamp 1682952543
transform 1 0 2316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8774
timestamp 1682952543
transform 1 0 2340 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8977
timestamp 1682952543
transform 1 0 2324 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8985
timestamp 1682952543
transform 1 0 2300 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8872
timestamp 1682952543
transform 1 0 2436 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8659
timestamp 1682952543
transform 1 0 2452 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8903
timestamp 1682952543
transform 1 0 2364 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8812
timestamp 1682952543
transform 1 0 2492 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8845
timestamp 1682952543
transform 1 0 2484 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8775
timestamp 1682952543
transform 1 0 2388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8776
timestamp 1682952543
transform 1 0 2444 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8777
timestamp 1682952543
transform 1 0 2460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8660
timestamp 1682952543
transform 1 0 2484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8778
timestamp 1682952543
transform 1 0 2484 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8831
timestamp 1682952543
transform 1 0 2476 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8944
timestamp 1682952543
transform 1 0 2484 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8591
timestamp 1682952543
transform 1 0 2524 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_8873
timestamp 1682952543
transform 1 0 2516 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8661
timestamp 1682952543
transform 1 0 2524 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8904
timestamp 1682952543
transform 1 0 2524 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8779
timestamp 1682952543
transform 1 0 2540 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8784
timestamp 1682952543
transform 1 0 2596 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8662
timestamp 1682952543
transform 1 0 2580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8663
timestamp 1682952543
transform 1 0 2588 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8978
timestamp 1682952543
transform 1 0 2580 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_8780
timestamp 1682952543
transform 1 0 2604 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8785
timestamp 1682952543
transform 1 0 2620 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8874
timestamp 1682952543
transform 1 0 2620 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8781
timestamp 1682952543
transform 1 0 2620 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8945
timestamp 1682952543
transform 1 0 2620 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8592
timestamp 1682952543
transform 1 0 2692 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8664
timestamp 1682952543
transform 1 0 2644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8665
timestamp 1682952543
transform 1 0 2652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8666
timestamp 1682952543
transform 1 0 2668 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8875
timestamp 1682952543
transform 1 0 2684 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8846
timestamp 1682952543
transform 1 0 2708 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8667
timestamp 1682952543
transform 1 0 2692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8668
timestamp 1682952543
transform 1 0 2700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8782
timestamp 1682952543
transform 1 0 2660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8783
timestamp 1682952543
transform 1 0 2676 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8784
timestamp 1682952543
transform 1 0 2708 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8785
timestamp 1682952543
transform 1 0 2716 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8946
timestamp 1682952543
transform 1 0 2716 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8786
timestamp 1682952543
transform 1 0 2780 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8786
timestamp 1682952543
transform 1 0 2812 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8669
timestamp 1682952543
transform 1 0 2812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8670
timestamp 1682952543
transform 1 0 2836 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8905
timestamp 1682952543
transform 1 0 2812 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8787
timestamp 1682952543
transform 1 0 2820 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8906
timestamp 1682952543
transform 1 0 2828 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8813
timestamp 1682952543
transform 1 0 2860 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8671
timestamp 1682952543
transform 1 0 2860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8788
timestamp 1682952543
transform 1 0 2844 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8947
timestamp 1682952543
transform 1 0 2820 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8907
timestamp 1682952543
transform 1 0 2852 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8876
timestamp 1682952543
transform 1 0 2916 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8847
timestamp 1682952543
transform 1 0 2988 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8672
timestamp 1682952543
transform 1 0 2948 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8673
timestamp 1682952543
transform 1 0 2964 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8789
timestamp 1682952543
transform 1 0 2868 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8790
timestamp 1682952543
transform 1 0 2924 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8986
timestamp 1682952543
transform 1 0 2940 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8877
timestamp 1682952543
transform 1 0 2972 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8674
timestamp 1682952543
transform 1 0 2980 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8675
timestamp 1682952543
transform 1 0 2996 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8676
timestamp 1682952543
transform 1 0 3012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8791
timestamp 1682952543
transform 1 0 2972 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8792
timestamp 1682952543
transform 1 0 2988 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8793
timestamp 1682952543
transform 1 0 3004 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8794
timestamp 1682952543
transform 1 0 3044 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8832
timestamp 1682952543
transform 1 0 3028 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8948
timestamp 1682952543
transform 1 0 3044 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8836
timestamp 1682952543
transform 1 0 3036 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_8979
timestamp 1682952543
transform 1 0 3036 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8908
timestamp 1682952543
transform 1 0 3076 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8814
timestamp 1682952543
transform 1 0 3100 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8677
timestamp 1682952543
transform 1 0 3100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8795
timestamp 1682952543
transform 1 0 3084 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8833
timestamp 1682952543
transform 1 0 3076 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8878
timestamp 1682952543
transform 1 0 3116 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8848
timestamp 1682952543
transform 1 0 3132 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8678
timestamp 1682952543
transform 1 0 3124 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8679
timestamp 1682952543
transform 1 0 3132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8796
timestamp 1682952543
transform 1 0 3108 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8909
timestamp 1682952543
transform 1 0 3124 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8797
timestamp 1682952543
transform 1 0 3132 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8815
timestamp 1682952543
transform 1 0 3148 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8798
timestamp 1682952543
transform 1 0 3164 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8910
timestamp 1682952543
transform 1 0 3172 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8949
timestamp 1682952543
transform 1 0 3164 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8849
timestamp 1682952543
transform 1 0 3196 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8879
timestamp 1682952543
transform 1 0 3188 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8680
timestamp 1682952543
transform 1 0 3196 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8880
timestamp 1682952543
transform 1 0 3204 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8799
timestamp 1682952543
transform 1 0 3204 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8968
timestamp 1682952543
transform 1 0 3196 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8681
timestamp 1682952543
transform 1 0 3220 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8881
timestamp 1682952543
transform 1 0 3252 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8800
timestamp 1682952543
transform 1 0 3268 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8950
timestamp 1682952543
transform 1 0 3268 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8850
timestamp 1682952543
transform 1 0 3316 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8851
timestamp 1682952543
transform 1 0 3340 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8682
timestamp 1682952543
transform 1 0 3332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8801
timestamp 1682952543
transform 1 0 3316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8802
timestamp 1682952543
transform 1 0 3324 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8911
timestamp 1682952543
transform 1 0 3332 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8951
timestamp 1682952543
transform 1 0 3332 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8683
timestamp 1682952543
transform 1 0 3348 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8912
timestamp 1682952543
transform 1 0 3356 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8803
timestamp 1682952543
transform 1 0 3364 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8969
timestamp 1682952543
transform 1 0 3348 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8787
timestamp 1682952543
transform 1 0 3380 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8684
timestamp 1682952543
transform 1 0 3380 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8913
timestamp 1682952543
transform 1 0 3380 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8804
timestamp 1682952543
transform 1 0 3404 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8970
timestamp 1682952543
transform 1 0 3404 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8788
timestamp 1682952543
transform 1 0 3540 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8816
timestamp 1682952543
transform 1 0 3508 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8817
timestamp 1682952543
transform 1 0 3540 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8852
timestamp 1682952543
transform 1 0 3492 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8853
timestamp 1682952543
transform 1 0 3516 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8685
timestamp 1682952543
transform 1 0 3492 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8882
timestamp 1682952543
transform 1 0 3524 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8883
timestamp 1682952543
transform 1 0 3572 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8805
timestamp 1682952543
transform 1 0 3476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8806
timestamp 1682952543
transform 1 0 3516 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8807
timestamp 1682952543
transform 1 0 3572 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8952
timestamp 1682952543
transform 1 0 3516 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8953
timestamp 1682952543
transform 1 0 3564 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8834
timestamp 1682952543
transform 1 0 3580 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8789
timestamp 1682952543
transform 1 0 3596 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8808
timestamp 1682952543
transform 1 0 3612 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8954
timestamp 1682952543
transform 1 0 3612 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8837
timestamp 1682952543
transform 1 0 3604 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_8884
timestamp 1682952543
transform 1 0 3628 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8790
timestamp 1682952543
transform 1 0 3644 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8791
timestamp 1682952543
transform 1 0 3676 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8686
timestamp 1682952543
transform 1 0 3644 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8885
timestamp 1682952543
transform 1 0 3652 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8818
timestamp 1682952543
transform 1 0 3700 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8854
timestamp 1682952543
transform 1 0 3692 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_8792
timestamp 1682952543
transform 1 0 3764 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8819
timestamp 1682952543
transform 1 0 3748 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8855
timestamp 1682952543
transform 1 0 3740 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8687
timestamp 1682952543
transform 1 0 3660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8688
timestamp 1682952543
transform 1 0 3668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8689
timestamp 1682952543
transform 1 0 3676 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8690
timestamp 1682952543
transform 1 0 3692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8691
timestamp 1682952543
transform 1 0 3708 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8692
timestamp 1682952543
transform 1 0 3724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8809
timestamp 1682952543
transform 1 0 3636 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8810
timestamp 1682952543
transform 1 0 3652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8835
timestamp 1682952543
transform 1 0 3628 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8914
timestamp 1682952543
transform 1 0 3676 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8811
timestamp 1682952543
transform 1 0 3684 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8812
timestamp 1682952543
transform 1 0 3700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8813
timestamp 1682952543
transform 1 0 3748 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8820
timestamp 1682952543
transform 1 0 3820 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8814
timestamp 1682952543
transform 1 0 3820 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8815
timestamp 1682952543
transform 1 0 3828 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8793
timestamp 1682952543
transform 1 0 3868 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8794
timestamp 1682952543
transform 1 0 3900 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8795
timestamp 1682952543
transform 1 0 3916 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8821
timestamp 1682952543
transform 1 0 3892 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8693
timestamp 1682952543
transform 1 0 3844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8694
timestamp 1682952543
transform 1 0 3852 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8695
timestamp 1682952543
transform 1 0 3860 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8886
timestamp 1682952543
transform 1 0 3868 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8915
timestamp 1682952543
transform 1 0 3860 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8822
timestamp 1682952543
transform 1 0 3916 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8823
timestamp 1682952543
transform 1 0 3932 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_8856
timestamp 1682952543
transform 1 0 3916 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8696
timestamp 1682952543
transform 1 0 3892 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8697
timestamp 1682952543
transform 1 0 3900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8698
timestamp 1682952543
transform 1 0 3916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8699
timestamp 1682952543
transform 1 0 3932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8816
timestamp 1682952543
transform 1 0 3868 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8817
timestamp 1682952543
transform 1 0 3884 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8955
timestamp 1682952543
transform 1 0 3860 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8916
timestamp 1682952543
transform 1 0 3900 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_8818
timestamp 1682952543
transform 1 0 3908 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8819
timestamp 1682952543
transform 1 0 3924 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8956
timestamp 1682952543
transform 1 0 3948 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8857
timestamp 1682952543
transform 1 0 3988 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8700
timestamp 1682952543
transform 1 0 3964 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8887
timestamp 1682952543
transform 1 0 4028 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8820
timestamp 1682952543
transform 1 0 3988 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8917
timestamp 1682952543
transform 1 0 4052 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8888
timestamp 1682952543
transform 1 0 4068 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8821
timestamp 1682952543
transform 1 0 4060 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8822
timestamp 1682952543
transform 1 0 4068 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8824
timestamp 1682952543
transform 1 0 4100 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8823
timestamp 1682952543
transform 1 0 4148 0 1 525
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_72
timestamp 1682952543
transform 1 0 24 0 1 470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_540
timestamp 1682952543
transform 1 0 72 0 -1 570
box -8 -3 104 105
use AOI22X1  AOI22X1_351
timestamp 1682952543
transform -1 0 208 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_609
timestamp 1682952543
transform 1 0 208 0 -1 570
box -9 -3 26 105
use FILL  FILL_3745
timestamp 1682952543
transform 1 0 224 0 -1 570
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1682952543
transform 1 0 232 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_382
timestamp 1682952543
transform -1 0 280 0 -1 570
box -8 -3 46 105
use FILL  FILL_3747
timestamp 1682952543
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1682952543
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1682952543
transform 1 0 296 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_352
timestamp 1682952543
transform -1 0 344 0 -1 570
box -8 -3 46 105
use FILL  FILL_3750
timestamp 1682952543
transform 1 0 344 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_541
timestamp 1682952543
transform 1 0 352 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_610
timestamp 1682952543
transform -1 0 464 0 -1 570
box -9 -3 26 105
use FILL  FILL_3751
timestamp 1682952543
transform 1 0 464 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_353
timestamp 1682952543
transform 1 0 472 0 -1 570
box -8 -3 46 105
use FILL  FILL_3752
timestamp 1682952543
transform 1 0 512 0 -1 570
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1682952543
transform 1 0 520 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_383
timestamp 1682952543
transform -1 0 568 0 -1 570
box -8 -3 46 105
use FILL  FILL_3754
timestamp 1682952543
transform 1 0 568 0 -1 570
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1682952543
transform 1 0 576 0 -1 570
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1682952543
transform 1 0 584 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_354
timestamp 1682952543
transform 1 0 592 0 -1 570
box -8 -3 46 105
use FILL  FILL_3757
timestamp 1682952543
transform 1 0 632 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_611
timestamp 1682952543
transform 1 0 640 0 -1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_542
timestamp 1682952543
transform -1 0 752 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_543
timestamp 1682952543
transform 1 0 752 0 -1 570
box -8 -3 104 105
use FILL  FILL_3758
timestamp 1682952543
transform 1 0 848 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_355
timestamp 1682952543
transform 1 0 856 0 -1 570
box -8 -3 46 105
use FILL  FILL_3759
timestamp 1682952543
transform 1 0 896 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_612
timestamp 1682952543
transform 1 0 904 0 -1 570
box -9 -3 26 105
use OAI21X1  OAI21X1_152
timestamp 1682952543
transform 1 0 920 0 -1 570
box -8 -3 34 105
use FILL  FILL_3760
timestamp 1682952543
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_3761
timestamp 1682952543
transform 1 0 960 0 -1 570
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1682952543
transform 1 0 968 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_102
timestamp 1682952543
transform 1 0 976 0 -1 570
box -8 -3 32 105
use FILL  FILL_3763
timestamp 1682952543
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_153
timestamp 1682952543
transform 1 0 1008 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_154
timestamp 1682952543
transform -1 0 1072 0 -1 570
box -8 -3 34 105
use M3_M2  M3_M2_8987
timestamp 1682952543
transform 1 0 1100 0 1 475
box -3 -3 3 3
use OAI21X1  OAI21X1_155
timestamp 1682952543
transform -1 0 1104 0 -1 570
box -8 -3 34 105
use OAI21X1  OAI21X1_156
timestamp 1682952543
transform -1 0 1136 0 -1 570
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_544
timestamp 1682952543
transform -1 0 1232 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_545
timestamp 1682952543
transform 1 0 1232 0 -1 570
box -8 -3 104 105
use M3_M2  M3_M2_8988
timestamp 1682952543
transform 1 0 1340 0 1 475
box -3 -3 3 3
use INVX2  INVX2_613
timestamp 1682952543
transform 1 0 1328 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_384
timestamp 1682952543
transform -1 0 1384 0 -1 570
box -8 -3 46 105
use FILL  FILL_3764
timestamp 1682952543
transform 1 0 1384 0 -1 570
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1682952543
transform 1 0 1392 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_546
timestamp 1682952543
transform 1 0 1400 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_614
timestamp 1682952543
transform -1 0 1512 0 -1 570
box -9 -3 26 105
use FILL  FILL_3766
timestamp 1682952543
transform 1 0 1512 0 -1 570
box -8 -3 16 105
use FILL  FILL_3767
timestamp 1682952543
transform 1 0 1520 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8989
timestamp 1682952543
transform 1 0 1540 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_356
timestamp 1682952543
transform 1 0 1528 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_8990
timestamp 1682952543
transform 1 0 1580 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_385
timestamp 1682952543
transform 1 0 1568 0 -1 570
box -8 -3 46 105
use M3_M2  M3_M2_8991
timestamp 1682952543
transform 1 0 1620 0 1 475
box -3 -3 3 3
use FILL  FILL_3768
timestamp 1682952543
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_3769
timestamp 1682952543
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1682952543
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8992
timestamp 1682952543
transform 1 0 1644 0 1 475
box -3 -3 3 3
use AOI22X1  AOI22X1_357
timestamp 1682952543
transform 1 0 1632 0 -1 570
box -8 -3 46 105
use FILL  FILL_3771
timestamp 1682952543
transform 1 0 1672 0 -1 570
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1682952543
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_615
timestamp 1682952543
transform 1 0 1688 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_616
timestamp 1682952543
transform -1 0 1720 0 -1 570
box -9 -3 26 105
use FILL  FILL_3773
timestamp 1682952543
transform 1 0 1720 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_547
timestamp 1682952543
transform 1 0 1728 0 -1 570
box -8 -3 104 105
use AOI22X1  AOI22X1_358
timestamp 1682952543
transform 1 0 1824 0 -1 570
box -8 -3 46 105
use FILL  FILL_3774
timestamp 1682952543
transform 1 0 1864 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_157
timestamp 1682952543
transform 1 0 1872 0 -1 570
box -8 -3 34 105
use FILL  FILL_3775
timestamp 1682952543
transform 1 0 1904 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_104
timestamp 1682952543
transform 1 0 1912 0 -1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_162
timestamp 1682952543
transform -1 0 1968 0 -1 570
box -8 -3 34 105
use M3_M2  M3_M2_8993
timestamp 1682952543
transform 1 0 1996 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_8994
timestamp 1682952543
transform 1 0 2052 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_8995
timestamp 1682952543
transform 1 0 2068 0 1 475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_549
timestamp 1682952543
transform -1 0 2064 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_550
timestamp 1682952543
transform 1 0 2064 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_621
timestamp 1682952543
transform 1 0 2160 0 -1 570
box -9 -3 26 105
use BUFX2  BUFX2_101
timestamp 1682952543
transform -1 0 2200 0 -1 570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_551
timestamp 1682952543
transform 1 0 2200 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_622
timestamp 1682952543
transform 1 0 2296 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_388
timestamp 1682952543
transform 1 0 2312 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_552
timestamp 1682952543
transform 1 0 2352 0 -1 570
box -8 -3 104 105
use OAI21X1  OAI21X1_163
timestamp 1682952543
transform 1 0 2448 0 -1 570
box -8 -3 34 105
use FILL  FILL_3794
timestamp 1682952543
transform 1 0 2480 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_105
timestamp 1682952543
transform 1 0 2488 0 -1 570
box -5 -3 28 105
use FILL  FILL_3797
timestamp 1682952543
transform 1 0 2512 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_105
timestamp 1682952543
transform 1 0 2520 0 -1 570
box -8 -3 32 105
use FILL  FILL_3798
timestamp 1682952543
transform 1 0 2544 0 -1 570
box -8 -3 16 105
use FILL  FILL_3799
timestamp 1682952543
transform 1 0 2552 0 -1 570
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1682952543
transform 1 0 2560 0 -1 570
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1682952543
transform 1 0 2568 0 -1 570
box -8 -3 16 105
use FILL  FILL_3802
timestamp 1682952543
transform 1 0 2576 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_624
timestamp 1682952543
transform 1 0 2584 0 -1 570
box -9 -3 26 105
use FILL  FILL_3803
timestamp 1682952543
transform 1 0 2600 0 -1 570
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1682952543
transform 1 0 2608 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_106
timestamp 1682952543
transform 1 0 2616 0 -1 570
box -5 -3 28 105
use FILL  FILL_3805
timestamp 1682952543
transform 1 0 2640 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_390
timestamp 1682952543
transform -1 0 2688 0 -1 570
box -8 -3 46 105
use NOR2X1  NOR2X1_106
timestamp 1682952543
transform 1 0 2688 0 -1 570
box -8 -3 32 105
use M3_M2  M3_M2_8996
timestamp 1682952543
transform 1 0 2724 0 1 475
box -3 -3 3 3
use FILL  FILL_3822
timestamp 1682952543
transform 1 0 2712 0 -1 570
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1682952543
transform 1 0 2720 0 -1 570
box -8 -3 16 105
use FILL  FILL_3824
timestamp 1682952543
transform 1 0 2728 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8997
timestamp 1682952543
transform 1 0 2756 0 1 475
box -3 -3 3 3
use BUFX2  BUFX2_107
timestamp 1682952543
transform 1 0 2736 0 -1 570
box -5 -3 28 105
use M3_M2  M3_M2_8998
timestamp 1682952543
transform 1 0 2772 0 1 475
box -3 -3 3 3
use FILL  FILL_3825
timestamp 1682952543
transform 1 0 2760 0 -1 570
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1682952543
transform 1 0 2768 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8999
timestamp 1682952543
transform 1 0 2788 0 1 475
box -3 -3 3 3
use FILL  FILL_3827
timestamp 1682952543
transform 1 0 2776 0 -1 570
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1682952543
transform 1 0 2784 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_108
timestamp 1682952543
transform 1 0 2792 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_109
timestamp 1682952543
transform 1 0 2816 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_110
timestamp 1682952543
transform 1 0 2840 0 -1 570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_556
timestamp 1682952543
transform -1 0 2960 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_630
timestamp 1682952543
transform 1 0 2960 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_395
timestamp 1682952543
transform -1 0 3016 0 -1 570
box -8 -3 46 105
use FILL  FILL_3829
timestamp 1682952543
transform 1 0 3016 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_70
timestamp 1682952543
transform -1 0 3056 0 -1 570
box -8 -3 40 105
use FILL  FILL_3830
timestamp 1682952543
transform 1 0 3056 0 -1 570
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1682952543
transform 1 0 3064 0 -1 570
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1682952543
transform 1 0 3072 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_111
timestamp 1682952543
transform 1 0 3080 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_112
timestamp 1682952543
transform 1 0 3104 0 -1 570
box -5 -3 28 105
use FILL  FILL_3833
timestamp 1682952543
transform 1 0 3128 0 -1 570
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1682952543
transform 1 0 3136 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_362
timestamp 1682952543
transform 1 0 3144 0 -1 570
box -8 -3 46 105
use FILL  FILL_3835
timestamp 1682952543
transform 1 0 3184 0 -1 570
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1682952543
transform 1 0 3192 0 -1 570
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1682952543
transform 1 0 3200 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_557
timestamp 1682952543
transform 1 0 3208 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_631
timestamp 1682952543
transform 1 0 3304 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_632
timestamp 1682952543
transform -1 0 3336 0 -1 570
box -9 -3 26 105
use FILL  FILL_3838
timestamp 1682952543
transform 1 0 3336 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_633
timestamp 1682952543
transform 1 0 3344 0 -1 570
box -9 -3 26 105
use FILL  FILL_3839
timestamp 1682952543
transform 1 0 3360 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_9000
timestamp 1682952543
transform 1 0 3380 0 1 475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_561
timestamp 1682952543
transform 1 0 3368 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_638
timestamp 1682952543
transform 1 0 3464 0 -1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_562
timestamp 1682952543
transform 1 0 3480 0 -1 570
box -8 -3 104 105
use FILL  FILL_3850
timestamp 1682952543
transform 1 0 3576 0 -1 570
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1682952543
transform 1 0 3584 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_72
timestamp 1682952543
transform -1 0 3624 0 -1 570
box -8 -3 40 105
use FILL  FILL_3852
timestamp 1682952543
transform 1 0 3624 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_366
timestamp 1682952543
transform 1 0 3632 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_401
timestamp 1682952543
transform 1 0 3672 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_563
timestamp 1682952543
transform 1 0 3712 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_639
timestamp 1682952543
transform 1 0 3808 0 -1 570
box -9 -3 26 105
use FILL  FILL_3853
timestamp 1682952543
transform 1 0 3824 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_640
timestamp 1682952543
transform -1 0 3848 0 -1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_367
timestamp 1682952543
transform -1 0 3888 0 -1 570
box -8 -3 46 105
use FILL  FILL_3854
timestamp 1682952543
transform 1 0 3888 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_402
timestamp 1682952543
transform -1 0 3936 0 -1 570
box -8 -3 46 105
use FILL  FILL_3855
timestamp 1682952543
transform 1 0 3936 0 -1 570
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1682952543
transform 1 0 3944 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_564
timestamp 1682952543
transform 1 0 3952 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_641
timestamp 1682952543
transform 1 0 4048 0 -1 570
box -9 -3 26 105
use FILL  FILL_3857
timestamp 1682952543
transform 1 0 4064 0 -1 570
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1682952543
transform 1 0 4072 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_642
timestamp 1682952543
transform -1 0 4096 0 -1 570
box -9 -3 26 105
use FILL  FILL_3859
timestamp 1682952543
transform 1 0 4096 0 -1 570
box -8 -3 16 105
use FILL  FILL_3860
timestamp 1682952543
transform 1 0 4104 0 -1 570
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1682952543
transform 1 0 4112 0 -1 570
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1682952543
transform 1 0 4120 0 -1 570
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1682952543
transform 1 0 4128 0 -1 570
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1682952543
transform 1 0 4136 0 -1 570
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1682952543
transform 1 0 4144 0 -1 570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_73
timestamp 1682952543
transform 1 0 4201 0 1 470
box -10 -3 10 3
use M2_M1  M2_M1_8849
timestamp 1682952543
transform 1 0 108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8850
timestamp 1682952543
transform 1 0 164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8851
timestamp 1682952543
transform 1 0 172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8972
timestamp 1682952543
transform 1 0 84 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9132
timestamp 1682952543
transform 1 0 132 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9154
timestamp 1682952543
transform 1 0 164 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9073
timestamp 1682952543
transform 1 0 196 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9074
timestamp 1682952543
transform 1 0 220 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9075
timestamp 1682952543
transform 1 0 284 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9076
timestamp 1682952543
transform 1 0 324 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8852
timestamp 1682952543
transform 1 0 188 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8853
timestamp 1682952543
transform 1 0 204 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9107
timestamp 1682952543
transform 1 0 212 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8854
timestamp 1682952543
transform 1 0 220 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8855
timestamp 1682952543
transform 1 0 284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8856
timestamp 1682952543
transform 1 0 316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8857
timestamp 1682952543
transform 1 0 324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8973
timestamp 1682952543
transform 1 0 180 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8974
timestamp 1682952543
transform 1 0 188 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9133
timestamp 1682952543
transform 1 0 204 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_8975
timestamp 1682952543
transform 1 0 212 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9155
timestamp 1682952543
transform 1 0 188 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_8976
timestamp 1682952543
transform 1 0 236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8977
timestamp 1682952543
transform 1 0 324 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9156
timestamp 1682952543
transform 1 0 300 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_8978
timestamp 1682952543
transform 1 0 340 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9157
timestamp 1682952543
transform 1 0 340 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9024
timestamp 1682952543
transform 1 0 468 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9044
timestamp 1682952543
transform 1 0 444 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9077
timestamp 1682952543
transform 1 0 412 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9078
timestamp 1682952543
transform 1 0 452 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9045
timestamp 1682952543
transform 1 0 492 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8858
timestamp 1682952543
transform 1 0 348 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8859
timestamp 1682952543
transform 1 0 412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8860
timestamp 1682952543
transform 1 0 444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8861
timestamp 1682952543
transform 1 0 452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8979
timestamp 1682952543
transform 1 0 364 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9108
timestamp 1682952543
transform 1 0 460 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8862
timestamp 1682952543
transform 1 0 468 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9109
timestamp 1682952543
transform 1 0 476 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8863
timestamp 1682952543
transform 1 0 484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8864
timestamp 1682952543
transform 1 0 508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8980
timestamp 1682952543
transform 1 0 468 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8981
timestamp 1682952543
transform 1 0 476 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8982
timestamp 1682952543
transform 1 0 492 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8983
timestamp 1682952543
transform 1 0 500 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9158
timestamp 1682952543
transform 1 0 436 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9046
timestamp 1682952543
transform 1 0 516 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9001
timestamp 1682952543
transform 1 0 556 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9025
timestamp 1682952543
transform 1 0 556 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9079
timestamp 1682952543
transform 1 0 540 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9026
timestamp 1682952543
transform 1 0 596 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9047
timestamp 1682952543
transform 1 0 580 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9080
timestamp 1682952543
transform 1 0 572 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8865
timestamp 1682952543
transform 1 0 548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8866
timestamp 1682952543
transform 1 0 556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8867
timestamp 1682952543
transform 1 0 572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8868
timestamp 1682952543
transform 1 0 596 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8984
timestamp 1682952543
transform 1 0 532 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8985
timestamp 1682952543
transform 1 0 540 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9159
timestamp 1682952543
transform 1 0 532 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9134
timestamp 1682952543
transform 1 0 548 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_8986
timestamp 1682952543
transform 1 0 564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8987
timestamp 1682952543
transform 1 0 580 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8988
timestamp 1682952543
transform 1 0 596 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9160
timestamp 1682952543
transform 1 0 572 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9027
timestamp 1682952543
transform 1 0 628 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9048
timestamp 1682952543
transform 1 0 612 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9081
timestamp 1682952543
transform 1 0 604 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9082
timestamp 1682952543
transform 1 0 668 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8869
timestamp 1682952543
transform 1 0 604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8870
timestamp 1682952543
transform 1 0 612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8871
timestamp 1682952543
transform 1 0 644 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9110
timestamp 1682952543
transform 1 0 692 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_9135
timestamp 1682952543
transform 1 0 644 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_8989
timestamp 1682952543
transform 1 0 692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8840
timestamp 1682952543
transform 1 0 732 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_8990
timestamp 1682952543
transform 1 0 716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9077
timestamp 1682952543
transform 1 0 708 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_9205
timestamp 1682952543
transform 1 0 660 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9206
timestamp 1682952543
transform 1 0 708 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9002
timestamp 1682952543
transform 1 0 780 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9009
timestamp 1682952543
transform 1 0 756 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9111
timestamp 1682952543
transform 1 0 740 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_9083
timestamp 1682952543
transform 1 0 780 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9003
timestamp 1682952543
transform 1 0 844 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9004
timestamp 1682952543
transform 1 0 868 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9028
timestamp 1682952543
transform 1 0 820 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_8872
timestamp 1682952543
transform 1 0 756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8873
timestamp 1682952543
transform 1 0 764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8874
timestamp 1682952543
transform 1 0 780 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9112
timestamp 1682952543
transform 1 0 788 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8875
timestamp 1682952543
transform 1 0 796 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8876
timestamp 1682952543
transform 1 0 820 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8991
timestamp 1682952543
transform 1 0 756 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8992
timestamp 1682952543
transform 1 0 780 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8993
timestamp 1682952543
transform 1 0 788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8994
timestamp 1682952543
transform 1 0 804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8995
timestamp 1682952543
transform 1 0 820 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9161
timestamp 1682952543
transform 1 0 756 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9207
timestamp 1682952543
transform 1 0 740 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9010
timestamp 1682952543
transform 1 0 940 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9029
timestamp 1682952543
transform 1 0 868 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9030
timestamp 1682952543
transform 1 0 892 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9031
timestamp 1682952543
transform 1 0 908 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9032
timestamp 1682952543
transform 1 0 972 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9049
timestamp 1682952543
transform 1 0 876 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9050
timestamp 1682952543
transform 1 0 916 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8877
timestamp 1682952543
transform 1 0 828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8878
timestamp 1682952543
transform 1 0 836 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9113
timestamp 1682952543
transform 1 0 844 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8879
timestamp 1682952543
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8880
timestamp 1682952543
transform 1 0 868 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8881
timestamp 1682952543
transform 1 0 876 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9162
timestamp 1682952543
transform 1 0 804 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9163
timestamp 1682952543
transform 1 0 820 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9114
timestamp 1682952543
transform 1 0 916 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8882
timestamp 1682952543
transform 1 0 924 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8883
timestamp 1682952543
transform 1 0 972 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8996
timestamp 1682952543
transform 1 0 844 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8997
timestamp 1682952543
transform 1 0 868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8998
timestamp 1682952543
transform 1 0 956 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_8999
timestamp 1682952543
transform 1 0 972 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9164
timestamp 1682952543
transform 1 0 852 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9165
timestamp 1682952543
transform 1 0 868 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9166
timestamp 1682952543
transform 1 0 916 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9167
timestamp 1682952543
transform 1 0 956 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9005
timestamp 1682952543
transform 1 0 1020 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9006
timestamp 1682952543
transform 1 0 1052 0 1 465
box -3 -3 3 3
use M2_M1  M2_M1_8884
timestamp 1682952543
transform 1 0 996 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9115
timestamp 1682952543
transform 1 0 1012 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8885
timestamp 1682952543
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8886
timestamp 1682952543
transform 1 0 1092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9000
timestamp 1682952543
transform 1 0 988 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9136
timestamp 1682952543
transform 1 0 996 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9001
timestamp 1682952543
transform 1 0 1012 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9137
timestamp 1682952543
transform 1 0 1036 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9168
timestamp 1682952543
transform 1 0 1012 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9033
timestamp 1682952543
transform 1 0 1124 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9034
timestamp 1682952543
transform 1 0 1172 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_8887
timestamp 1682952543
transform 1 0 1116 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8888
timestamp 1682952543
transform 1 0 1180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9002
timestamp 1682952543
transform 1 0 1108 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9078
timestamp 1682952543
transform 1 0 1100 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_9003
timestamp 1682952543
transform 1 0 1132 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9138
timestamp 1682952543
transform 1 0 1180 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9208
timestamp 1682952543
transform 1 0 1132 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9209
timestamp 1682952543
transform 1 0 1164 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9051
timestamp 1682952543
transform 1 0 1228 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8889
timestamp 1682952543
transform 1 0 1228 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8890
timestamp 1682952543
transform 1 0 1292 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9004
timestamp 1682952543
transform 1 0 1244 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9169
timestamp 1682952543
transform 1 0 1292 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9210
timestamp 1682952543
transform 1 0 1228 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_8891
timestamp 1682952543
transform 1 0 1340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8892
timestamp 1682952543
transform 1 0 1356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8893
timestamp 1682952543
transform 1 0 1372 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9116
timestamp 1682952543
transform 1 0 1380 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9005
timestamp 1682952543
transform 1 0 1348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9006
timestamp 1682952543
transform 1 0 1364 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9007
timestamp 1682952543
transform 1 0 1380 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9008
timestamp 1682952543
transform 1 0 1388 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9170
timestamp 1682952543
transform 1 0 1364 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9052
timestamp 1682952543
transform 1 0 1412 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8894
timestamp 1682952543
transform 1 0 1396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8895
timestamp 1682952543
transform 1 0 1412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8896
timestamp 1682952543
transform 1 0 1428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9009
timestamp 1682952543
transform 1 0 1404 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9139
timestamp 1682952543
transform 1 0 1412 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9053
timestamp 1682952543
transform 1 0 1532 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8897
timestamp 1682952543
transform 1 0 1500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8898
timestamp 1682952543
transform 1 0 1532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8899
timestamp 1682952543
transform 1 0 1540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9010
timestamp 1682952543
transform 1 0 1420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9011
timestamp 1682952543
transform 1 0 1436 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9012
timestamp 1682952543
transform 1 0 1452 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9171
timestamp 1682952543
transform 1 0 1396 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9172
timestamp 1682952543
transform 1 0 1428 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9211
timestamp 1682952543
transform 1 0 1380 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9140
timestamp 1682952543
transform 1 0 1500 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9141
timestamp 1682952543
transform 1 0 1540 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9212
timestamp 1682952543
transform 1 0 1484 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9011
timestamp 1682952543
transform 1 0 1588 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9054
timestamp 1682952543
transform 1 0 1564 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9084
timestamp 1682952543
transform 1 0 1588 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8900
timestamp 1682952543
transform 1 0 1556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8901
timestamp 1682952543
transform 1 0 1572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8902
timestamp 1682952543
transform 1 0 1588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9013
timestamp 1682952543
transform 1 0 1556 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9014
timestamp 1682952543
transform 1 0 1564 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9015
timestamp 1682952543
transform 1 0 1580 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9055
timestamp 1682952543
transform 1 0 1620 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9085
timestamp 1682952543
transform 1 0 1604 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9086
timestamp 1682952543
transform 1 0 1636 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9056
timestamp 1682952543
transform 1 0 1692 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8903
timestamp 1682952543
transform 1 0 1612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8904
timestamp 1682952543
transform 1 0 1620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8905
timestamp 1682952543
transform 1 0 1636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8906
timestamp 1682952543
transform 1 0 1660 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8907
timestamp 1682952543
transform 1 0 1692 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9016
timestamp 1682952543
transform 1 0 1604 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9142
timestamp 1682952543
transform 1 0 1612 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9017
timestamp 1682952543
transform 1 0 1620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9018
timestamp 1682952543
transform 1 0 1644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9019
timestamp 1682952543
transform 1 0 1652 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9143
timestamp 1682952543
transform 1 0 1692 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9020
timestamp 1682952543
transform 1 0 1740 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9057
timestamp 1682952543
transform 1 0 1796 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9087
timestamp 1682952543
transform 1 0 1804 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9035
timestamp 1682952543
transform 1 0 1876 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9058
timestamp 1682952543
transform 1 0 1868 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9088
timestamp 1682952543
transform 1 0 1860 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8908
timestamp 1682952543
transform 1 0 1804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8909
timestamp 1682952543
transform 1 0 1844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8910
timestamp 1682952543
transform 1 0 1860 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9021
timestamp 1682952543
transform 1 0 1764 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9012
timestamp 1682952543
transform 1 0 1900 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9059
timestamp 1682952543
transform 1 0 1884 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8911
timestamp 1682952543
transform 1 0 1876 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9022
timestamp 1682952543
transform 1 0 1868 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9023
timestamp 1682952543
transform 1 0 1876 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9173
timestamp 1682952543
transform 1 0 1844 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9174
timestamp 1682952543
transform 1 0 1860 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9175
timestamp 1682952543
transform 1 0 1876 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9013
timestamp 1682952543
transform 1 0 1924 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9060
timestamp 1682952543
transform 1 0 1908 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8841
timestamp 1682952543
transform 1 0 1908 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9024
timestamp 1682952543
transform 1 0 1916 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9079
timestamp 1682952543
transform 1 0 1908 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_9061
timestamp 1682952543
transform 1 0 1940 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8912
timestamp 1682952543
transform 1 0 1932 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9025
timestamp 1682952543
transform 1 0 1932 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9026
timestamp 1682952543
transform 1 0 1940 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9176
timestamp 1682952543
transform 1 0 1932 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9036
timestamp 1682952543
transform 1 0 1956 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_8842
timestamp 1682952543
transform 1 0 1948 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_8913
timestamp 1682952543
transform 1 0 1964 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9177
timestamp 1682952543
transform 1 0 1956 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9027
timestamp 1682952543
transform 1 0 1980 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9178
timestamp 1682952543
transform 1 0 1980 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_8914
timestamp 1682952543
transform 1 0 2036 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9028
timestamp 1682952543
transform 1 0 1996 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9144
timestamp 1682952543
transform 1 0 2020 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9179
timestamp 1682952543
transform 1 0 2044 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_8915
timestamp 1682952543
transform 1 0 2092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9029
timestamp 1682952543
transform 1 0 2100 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9180
timestamp 1682952543
transform 1 0 2092 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_8916
timestamp 1682952543
transform 1 0 2116 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8917
timestamp 1682952543
transform 1 0 2132 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9117
timestamp 1682952543
transform 1 0 2140 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9030
timestamp 1682952543
transform 1 0 2124 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9031
timestamp 1682952543
transform 1 0 2140 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9089
timestamp 1682952543
transform 1 0 2156 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8918
timestamp 1682952543
transform 1 0 2156 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9090
timestamp 1682952543
transform 1 0 2180 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8919
timestamp 1682952543
transform 1 0 2180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9032
timestamp 1682952543
transform 1 0 2172 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9091
timestamp 1682952543
transform 1 0 2260 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8920
timestamp 1682952543
transform 1 0 2260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9033
timestamp 1682952543
transform 1 0 2196 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9034
timestamp 1682952543
transform 1 0 2212 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9092
timestamp 1682952543
transform 1 0 2332 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8921
timestamp 1682952543
transform 1 0 2340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8843
timestamp 1682952543
transform 1 0 2380 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_8922
timestamp 1682952543
transform 1 0 2364 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9014
timestamp 1682952543
transform 1 0 2396 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9007
timestamp 1682952543
transform 1 0 2460 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_9015
timestamp 1682952543
transform 1 0 2460 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9016
timestamp 1682952543
transform 1 0 2492 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9017
timestamp 1682952543
transform 1 0 2516 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9062
timestamp 1682952543
transform 1 0 2420 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9063
timestamp 1682952543
transform 1 0 2436 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8844
timestamp 1682952543
transform 1 0 2388 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_9093
timestamp 1682952543
transform 1 0 2396 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9118
timestamp 1682952543
transform 1 0 2388 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_9094
timestamp 1682952543
transform 1 0 2532 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8923
timestamp 1682952543
transform 1 0 2396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8924
timestamp 1682952543
transform 1 0 2412 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8925
timestamp 1682952543
transform 1 0 2428 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8926
timestamp 1682952543
transform 1 0 2436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8927
timestamp 1682952543
transform 1 0 2468 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9119
timestamp 1682952543
transform 1 0 2476 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_9095
timestamp 1682952543
transform 1 0 2572 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9096
timestamp 1682952543
transform 1 0 2612 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8928
timestamp 1682952543
transform 1 0 2532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8929
timestamp 1682952543
transform 1 0 2548 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9035
timestamp 1682952543
transform 1 0 2388 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9036
timestamp 1682952543
transform 1 0 2404 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9037
timestamp 1682952543
transform 1 0 2420 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9145
timestamp 1682952543
transform 1 0 2436 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9146
timestamp 1682952543
transform 1 0 2468 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9038
timestamp 1682952543
transform 1 0 2516 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9181
timestamp 1682952543
transform 1 0 2452 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9182
timestamp 1682952543
transform 1 0 2492 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9213
timestamp 1682952543
transform 1 0 2444 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9214
timestamp 1682952543
transform 1 0 2468 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9120
timestamp 1682952543
transform 1 0 2556 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8930
timestamp 1682952543
transform 1 0 2564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8931
timestamp 1682952543
transform 1 0 2572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8932
timestamp 1682952543
transform 1 0 2604 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9121
timestamp 1682952543
transform 1 0 2652 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9039
timestamp 1682952543
transform 1 0 2540 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9147
timestamp 1682952543
transform 1 0 2548 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9040
timestamp 1682952543
transform 1 0 2564 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9148
timestamp 1682952543
transform 1 0 2572 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9041
timestamp 1682952543
transform 1 0 2652 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9183
timestamp 1682952543
transform 1 0 2628 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9184
timestamp 1682952543
transform 1 0 2652 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9064
timestamp 1682952543
transform 1 0 2684 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8933
timestamp 1682952543
transform 1 0 2684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8934
timestamp 1682952543
transform 1 0 2700 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9122
timestamp 1682952543
transform 1 0 2708 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_9018
timestamp 1682952543
transform 1 0 2740 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_8935
timestamp 1682952543
transform 1 0 2724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8936
timestamp 1682952543
transform 1 0 2732 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9149
timestamp 1682952543
transform 1 0 2684 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9042
timestamp 1682952543
transform 1 0 2692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9043
timestamp 1682952543
transform 1 0 2708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9044
timestamp 1682952543
transform 1 0 2716 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9045
timestamp 1682952543
transform 1 0 2740 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9123
timestamp 1682952543
transform 1 0 2756 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_9150
timestamp 1682952543
transform 1 0 2764 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_8937
timestamp 1682952543
transform 1 0 2780 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9215
timestamp 1682952543
transform 1 0 2772 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_8845
timestamp 1682952543
transform 1 0 2804 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9046
timestamp 1682952543
transform 1 0 2796 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9151
timestamp 1682952543
transform 1 0 2804 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_9037
timestamp 1682952543
transform 1 0 2836 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_8838
timestamp 1682952543
transform 1 0 2836 0 1 435
box -2 -2 2 2
use M3_M2  M3_M2_9097
timestamp 1682952543
transform 1 0 2844 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9019
timestamp 1682952543
transform 1 0 2916 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9038
timestamp 1682952543
transform 1 0 2916 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_8846
timestamp 1682952543
transform 1 0 2852 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_8938
timestamp 1682952543
transform 1 0 2844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8939
timestamp 1682952543
transform 1 0 2916 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9124
timestamp 1682952543
transform 1 0 2940 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9047
timestamp 1682952543
transform 1 0 2868 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9185
timestamp 1682952543
transform 1 0 2908 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9216
timestamp 1682952543
transform 1 0 2860 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9020
timestamp 1682952543
transform 1 0 2956 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9048
timestamp 1682952543
transform 1 0 2956 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9186
timestamp 1682952543
transform 1 0 2956 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9217
timestamp 1682952543
transform 1 0 2948 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_8940
timestamp 1682952543
transform 1 0 2964 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9039
timestamp 1682952543
transform 1 0 2996 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9098
timestamp 1682952543
transform 1 0 2980 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9040
timestamp 1682952543
transform 1 0 3012 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_8941
timestamp 1682952543
transform 1 0 2980 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8942
timestamp 1682952543
transform 1 0 3004 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9125
timestamp 1682952543
transform 1 0 3012 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9049
timestamp 1682952543
transform 1 0 2988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9050
timestamp 1682952543
transform 1 0 3004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9051
timestamp 1682952543
transform 1 0 3012 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9187
timestamp 1682952543
transform 1 0 2972 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9218
timestamp 1682952543
transform 1 0 2988 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9188
timestamp 1682952543
transform 1 0 3012 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9021
timestamp 1682952543
transform 1 0 3028 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9022
timestamp 1682952543
transform 1 0 3060 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9065
timestamp 1682952543
transform 1 0 3044 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9099
timestamp 1682952543
transform 1 0 3060 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8943
timestamp 1682952543
transform 1 0 3028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8944
timestamp 1682952543
transform 1 0 3044 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9126
timestamp 1682952543
transform 1 0 3052 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8945
timestamp 1682952543
transform 1 0 3060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9052
timestamp 1682952543
transform 1 0 3052 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9066
timestamp 1682952543
transform 1 0 3132 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9100
timestamp 1682952543
transform 1 0 3132 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8839
timestamp 1682952543
transform 1 0 3196 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_8847
timestamp 1682952543
transform 1 0 3188 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_8946
timestamp 1682952543
transform 1 0 3124 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9053
timestamp 1682952543
transform 1 0 3172 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9189
timestamp 1682952543
transform 1 0 3148 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9219
timestamp 1682952543
transform 1 0 3124 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9220
timestamp 1682952543
transform 1 0 3172 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9101
timestamp 1682952543
transform 1 0 3204 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8947
timestamp 1682952543
transform 1 0 3204 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9190
timestamp 1682952543
transform 1 0 3204 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9067
timestamp 1682952543
transform 1 0 3236 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8848
timestamp 1682952543
transform 1 0 3228 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_9023
timestamp 1682952543
transform 1 0 3268 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_9102
timestamp 1682952543
transform 1 0 3252 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9103
timestamp 1682952543
transform 1 0 3268 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8948
timestamp 1682952543
transform 1 0 3236 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9127
timestamp 1682952543
transform 1 0 3244 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8949
timestamp 1682952543
transform 1 0 3252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8950
timestamp 1682952543
transform 1 0 3268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8951
timestamp 1682952543
transform 1 0 3276 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9054
timestamp 1682952543
transform 1 0 3244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9055
timestamp 1682952543
transform 1 0 3268 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9191
timestamp 1682952543
transform 1 0 3268 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9041
timestamp 1682952543
transform 1 0 3316 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9042
timestamp 1682952543
transform 1 0 3348 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9068
timestamp 1682952543
transform 1 0 3324 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8952
timestamp 1682952543
transform 1 0 3324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8953
timestamp 1682952543
transform 1 0 3340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9056
timestamp 1682952543
transform 1 0 3308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9057
timestamp 1682952543
transform 1 0 3316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9058
timestamp 1682952543
transform 1 0 3332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9059
timestamp 1682952543
transform 1 0 3348 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9060
timestamp 1682952543
transform 1 0 3356 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9192
timestamp 1682952543
transform 1 0 3332 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_8954
timestamp 1682952543
transform 1 0 3364 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9128
timestamp 1682952543
transform 1 0 3388 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8955
timestamp 1682952543
transform 1 0 3396 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9152
timestamp 1682952543
transform 1 0 3380 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9061
timestamp 1682952543
transform 1 0 3388 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9062
timestamp 1682952543
transform 1 0 3404 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9193
timestamp 1682952543
transform 1 0 3388 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9008
timestamp 1682952543
transform 1 0 3460 0 1 465
box -3 -3 3 3
use M2_M1  M2_M1_8956
timestamp 1682952543
transform 1 0 3452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9063
timestamp 1682952543
transform 1 0 3428 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9194
timestamp 1682952543
transform 1 0 3452 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9195
timestamp 1682952543
transform 1 0 3492 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9221
timestamp 1682952543
transform 1 0 3428 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9129
timestamp 1682952543
transform 1 0 3524 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8957
timestamp 1682952543
transform 1 0 3532 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9130
timestamp 1682952543
transform 1 0 3556 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8958
timestamp 1682952543
transform 1 0 3580 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8959
timestamp 1682952543
transform 1 0 3636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9064
timestamp 1682952543
transform 1 0 3556 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9196
timestamp 1682952543
transform 1 0 3556 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9197
timestamp 1682952543
transform 1 0 3628 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9222
timestamp 1682952543
transform 1 0 3644 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9104
timestamp 1682952543
transform 1 0 3660 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_9105
timestamp 1682952543
transform 1 0 3684 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8960
timestamp 1682952543
transform 1 0 3668 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8961
timestamp 1682952543
transform 1 0 3684 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_9131
timestamp 1682952543
transform 1 0 3708 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_8962
timestamp 1682952543
transform 1 0 3732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9065
timestamp 1682952543
transform 1 0 3660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9066
timestamp 1682952543
transform 1 0 3676 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9067
timestamp 1682952543
transform 1 0 3692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9068
timestamp 1682952543
transform 1 0 3708 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9198
timestamp 1682952543
transform 1 0 3660 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9199
timestamp 1682952543
transform 1 0 3676 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9200
timestamp 1682952543
transform 1 0 3732 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9223
timestamp 1682952543
transform 1 0 3700 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9043
timestamp 1682952543
transform 1 0 3820 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_9069
timestamp 1682952543
transform 1 0 3844 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9106
timestamp 1682952543
transform 1 0 3812 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_8963
timestamp 1682952543
transform 1 0 3812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8964
timestamp 1682952543
transform 1 0 3828 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8965
timestamp 1682952543
transform 1 0 3844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8966
timestamp 1682952543
transform 1 0 3852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9069
timestamp 1682952543
transform 1 0 3820 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9070
timestamp 1682952543
transform 1 0 3836 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9153
timestamp 1682952543
transform 1 0 3844 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9071
timestamp 1682952543
transform 1 0 3852 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9201
timestamp 1682952543
transform 1 0 3836 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9070
timestamp 1682952543
transform 1 0 3916 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8967
timestamp 1682952543
transform 1 0 3908 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9072
timestamp 1682952543
transform 1 0 3956 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9202
timestamp 1682952543
transform 1 0 3908 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9224
timestamp 1682952543
transform 1 0 3892 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9225
timestamp 1682952543
transform 1 0 3924 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_9226
timestamp 1682952543
transform 1 0 3956 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9073
timestamp 1682952543
transform 1 0 3972 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9071
timestamp 1682952543
transform 1 0 3996 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_9072
timestamp 1682952543
transform 1 0 4012 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_8968
timestamp 1682952543
transform 1 0 3996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8969
timestamp 1682952543
transform 1 0 4020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9074
timestamp 1682952543
transform 1 0 4012 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9075
timestamp 1682952543
transform 1 0 4028 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9203
timestamp 1682952543
transform 1 0 4012 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9227
timestamp 1682952543
transform 1 0 4044 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_8970
timestamp 1682952543
transform 1 0 4084 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_8971
timestamp 1682952543
transform 1 0 4148 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9076
timestamp 1682952543
transform 1 0 4060 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_9204
timestamp 1682952543
transform 1 0 4084 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_9228
timestamp 1682952543
transform 1 0 4060 0 1 385
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_74
timestamp 1682952543
transform 1 0 48 0 1 370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_565
timestamp 1682952543
transform 1 0 72 0 1 370
box -8 -3 104 105
use INVX2  INVX2_643
timestamp 1682952543
transform -1 0 184 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_368
timestamp 1682952543
transform -1 0 224 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_9229
timestamp 1682952543
transform 1 0 284 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_566
timestamp 1682952543
transform 1 0 224 0 1 370
box -8 -3 104 105
use INVX2  INVX2_644
timestamp 1682952543
transform 1 0 320 0 1 370
box -9 -3 26 105
use INVX2  INVX2_645
timestamp 1682952543
transform 1 0 336 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_567
timestamp 1682952543
transform 1 0 352 0 1 370
box -8 -3 104 105
use INVX2  INVX2_646
timestamp 1682952543
transform -1 0 464 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_369
timestamp 1682952543
transform 1 0 464 0 1 370
box -8 -3 46 105
use INVX2  INVX2_647
timestamp 1682952543
transform -1 0 520 0 1 370
box -9 -3 26 105
use FILL  FILL_3866
timestamp 1682952543
transform 1 0 520 0 1 370
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1682952543
transform 1 0 528 0 1 370
box -8 -3 16 105
use INVX2  INVX2_648
timestamp 1682952543
transform 1 0 536 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_370
timestamp 1682952543
transform 1 0 552 0 1 370
box -8 -3 46 105
use INVX2  INVX2_649
timestamp 1682952543
transform 1 0 592 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_568
timestamp 1682952543
transform -1 0 704 0 1 370
box -8 -3 104 105
use NOR2X1  NOR2X1_107
timestamp 1682952543
transform 1 0 704 0 1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_164
timestamp 1682952543
transform -1 0 760 0 1 370
box -8 -3 34 105
use INVX2  INVX2_650
timestamp 1682952543
transform -1 0 776 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_371
timestamp 1682952543
transform 1 0 776 0 1 370
box -8 -3 46 105
use INVX2  INVX2_651
timestamp 1682952543
transform 1 0 816 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_372
timestamp 1682952543
transform 1 0 832 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_569
timestamp 1682952543
transform -1 0 968 0 1 370
box -8 -3 104 105
use INVX2  INVX2_652
timestamp 1682952543
transform 1 0 968 0 1 370
box -9 -3 26 105
use INVX2  INVX2_653
timestamp 1682952543
transform 1 0 984 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_9230
timestamp 1682952543
transform 1 0 1100 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_570
timestamp 1682952543
transform 1 0 1000 0 1 370
box -8 -3 104 105
use NOR2X1  NOR2X1_108
timestamp 1682952543
transform 1 0 1096 0 1 370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_571
timestamp 1682952543
transform 1 0 1120 0 1 370
box -8 -3 104 105
use INVX2  INVX2_654
timestamp 1682952543
transform 1 0 1216 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_572
timestamp 1682952543
transform 1 0 1232 0 1 370
box -8 -3 104 105
use INVX2  INVX2_655
timestamp 1682952543
transform 1 0 1328 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_9231
timestamp 1682952543
transform 1 0 1388 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_403
timestamp 1682952543
transform -1 0 1384 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_9232
timestamp 1682952543
transform 1 0 1404 0 1 375
box -3 -3 3 3
use INVX2  INVX2_656
timestamp 1682952543
transform 1 0 1384 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_9233
timestamp 1682952543
transform 1 0 1420 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_404
timestamp 1682952543
transform -1 0 1440 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_573
timestamp 1682952543
transform 1 0 1440 0 1 370
box -8 -3 104 105
use INVX2  INVX2_657
timestamp 1682952543
transform -1 0 1552 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_373
timestamp 1682952543
transform -1 0 1592 0 1 370
box -8 -3 46 105
use FILL  FILL_3868
timestamp 1682952543
transform 1 0 1592 0 1 370
box -8 -3 16 105
use INVX2  INVX2_658
timestamp 1682952543
transform 1 0 1600 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_374
timestamp 1682952543
transform 1 0 1616 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_574
timestamp 1682952543
transform -1 0 1752 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_575
timestamp 1682952543
transform 1 0 1752 0 1 370
box -8 -3 104 105
use INVX2  INVX2_659
timestamp 1682952543
transform -1 0 1864 0 1 370
box -9 -3 26 105
use FILL  FILL_3869
timestamp 1682952543
transform 1 0 1864 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_165
timestamp 1682952543
transform 1 0 1872 0 1 370
box -8 -3 34 105
use FILL  FILL_3870
timestamp 1682952543
transform 1 0 1904 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_109
timestamp 1682952543
transform 1 0 1912 0 1 370
box -8 -3 32 105
use FILL  FILL_3871
timestamp 1682952543
transform 1 0 1936 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_166
timestamp 1682952543
transform -1 0 1976 0 1 370
box -8 -3 34 105
use FILL  FILL_3872
timestamp 1682952543
transform 1 0 1976 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_576
timestamp 1682952543
transform 1 0 1984 0 1 370
box -8 -3 104 105
use INVX2  INVX2_660
timestamp 1682952543
transform 1 0 2080 0 1 370
box -9 -3 26 105
use FILL  FILL_3873
timestamp 1682952543
transform 1 0 2096 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_405
timestamp 1682952543
transform -1 0 2144 0 1 370
box -8 -3 46 105
use FILL  FILL_3874
timestamp 1682952543
transform 1 0 2144 0 1 370
box -8 -3 16 105
use BUFX2  BUFX2_113
timestamp 1682952543
transform 1 0 2152 0 1 370
box -5 -3 28 105
use BUFX2  BUFX2_114
timestamp 1682952543
transform 1 0 2176 0 1 370
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_577
timestamp 1682952543
transform 1 0 2200 0 1 370
box -8 -3 104 105
use M3_M2  M3_M2_9234
timestamp 1682952543
transform 1 0 2308 0 1 375
box -3 -3 3 3
use FILL  FILL_3875
timestamp 1682952543
transform 1 0 2296 0 1 370
box -8 -3 16 105
use INVX2  INVX2_661
timestamp 1682952543
transform 1 0 2304 0 1 370
box -9 -3 26 105
use FILL  FILL_3876
timestamp 1682952543
transform 1 0 2320 0 1 370
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1682952543
transform 1 0 2328 0 1 370
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1682952543
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1682952543
transform 1 0 2344 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_167
timestamp 1682952543
transform 1 0 2352 0 1 370
box -8 -3 34 105
use FILL  FILL_3880
timestamp 1682952543
transform 1 0 2384 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_375
timestamp 1682952543
transform 1 0 2392 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_578
timestamp 1682952543
transform -1 0 2528 0 1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_376
timestamp 1682952543
transform 1 0 2528 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_579
timestamp 1682952543
transform -1 0 2664 0 1 370
box -8 -3 104 105
use FILL  FILL_3881
timestamp 1682952543
transform 1 0 2664 0 1 370
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1682952543
transform 1 0 2672 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_377
timestamp 1682952543
transform 1 0 2680 0 1 370
box -8 -3 46 105
use INVX2  INVX2_662
timestamp 1682952543
transform 1 0 2720 0 1 370
box -9 -3 26 105
use BUFX2  BUFX2_115
timestamp 1682952543
transform -1 0 2760 0 1 370
box -5 -3 28 105
use FILL  FILL_3883
timestamp 1682952543
transform 1 0 2760 0 1 370
box -8 -3 16 105
use FILL  FILL_3884
timestamp 1682952543
transform 1 0 2768 0 1 370
box -8 -3 16 105
use BUFX2  BUFX2_116
timestamp 1682952543
transform 1 0 2776 0 1 370
box -5 -3 28 105
use FILL  FILL_3885
timestamp 1682952543
transform 1 0 2800 0 1 370
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1682952543
transform 1 0 2808 0 1 370
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1682952543
transform 1 0 2816 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_73
timestamp 1682952543
transform -1 0 2856 0 1 370
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_580
timestamp 1682952543
transform 1 0 2856 0 1 370
box -8 -3 104 105
use FILL  FILL_3888
timestamp 1682952543
transform 1 0 2952 0 1 370
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1682952543
transform 1 0 2960 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_9235
timestamp 1682952543
transform 1 0 3004 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_406
timestamp 1682952543
transform -1 0 3008 0 1 370
box -8 -3 46 105
use FILL  FILL_3890
timestamp 1682952543
transform 1 0 3008 0 1 370
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1682952543
transform 1 0 3016 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_9236
timestamp 1682952543
transform 1 0 3052 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_378
timestamp 1682952543
transform -1 0 3064 0 1 370
box -8 -3 46 105
use FILL  FILL_3892
timestamp 1682952543
transform 1 0 3064 0 1 370
box -8 -3 16 105
use INVX2  INVX2_663
timestamp 1682952543
transform -1 0 3088 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_581
timestamp 1682952543
transform -1 0 3184 0 1 370
box -8 -3 104 105
use NAND3X1  NAND3X1_74
timestamp 1682952543
transform -1 0 3216 0 1 370
box -8 -3 40 105
use FILL  FILL_3893
timestamp 1682952543
transform 1 0 3216 0 1 370
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1682952543
transform 1 0 3224 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_9237
timestamp 1682952543
transform 1 0 3260 0 1 375
box -3 -3 3 3
use AOI22X1  AOI22X1_379
timestamp 1682952543
transform 1 0 3232 0 1 370
box -8 -3 46 105
use INVX2  INVX2_664
timestamp 1682952543
transform -1 0 3288 0 1 370
box -9 -3 26 105
use FILL  FILL_3895
timestamp 1682952543
transform 1 0 3288 0 1 370
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1682952543
transform 1 0 3296 0 1 370
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1682952543
transform 1 0 3304 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_407
timestamp 1682952543
transform 1 0 3312 0 1 370
box -8 -3 46 105
use FILL  FILL_3898
timestamp 1682952543
transform 1 0 3352 0 1 370
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1682952543
transform 1 0 3360 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_421
timestamp 1682952543
transform 1 0 3368 0 1 370
box -8 -3 46 105
use FILL  FILL_3925
timestamp 1682952543
transform 1 0 3408 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_598
timestamp 1682952543
transform 1 0 3416 0 1 370
box -8 -3 104 105
use FILL  FILL_3926
timestamp 1682952543
transform 1 0 3512 0 1 370
box -8 -3 16 105
use INVX2  INVX2_676
timestamp 1682952543
transform 1 0 3520 0 1 370
box -9 -3 26 105
use FILL  FILL_3927
timestamp 1682952543
transform 1 0 3536 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_9238
timestamp 1682952543
transform 1 0 3564 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_9239
timestamp 1682952543
transform 1 0 3596 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_9240
timestamp 1682952543
transform 1 0 3612 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_9241
timestamp 1682952543
transform 1 0 3636 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_599
timestamp 1682952543
transform 1 0 3544 0 1 370
box -8 -3 104 105
use FILL  FILL_3928
timestamp 1682952543
transform 1 0 3640 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_9242
timestamp 1682952543
transform 1 0 3660 0 1 375
box -3 -3 3 3
use FILL  FILL_3929
timestamp 1682952543
transform 1 0 3648 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_422
timestamp 1682952543
transform 1 0 3656 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_601
timestamp 1682952543
transform 1 0 3696 0 1 370
box -8 -3 104 105
use FILL  FILL_3933
timestamp 1682952543
transform 1 0 3792 0 1 370
box -8 -3 16 105
use INVX2  INVX2_679
timestamp 1682952543
transform 1 0 3800 0 1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_425
timestamp 1682952543
transform -1 0 3856 0 1 370
box -8 -3 46 105
use FILL  FILL_3934
timestamp 1682952543
transform 1 0 3856 0 1 370
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1682952543
transform 1 0 3864 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_9243
timestamp 1682952543
transform 1 0 3932 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_9244
timestamp 1682952543
transform 1 0 3972 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_602
timestamp 1682952543
transform -1 0 3968 0 1 370
box -8 -3 104 105
use FILL  FILL_3936
timestamp 1682952543
transform 1 0 3968 0 1 370
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1682952543
transform 1 0 3976 0 1 370
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1682952543
transform 1 0 3984 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_426
timestamp 1682952543
transform 1 0 3992 0 1 370
box -8 -3 46 105
use FILL  FILL_3939
timestamp 1682952543
transform 1 0 4032 0 1 370
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1682952543
transform 1 0 4040 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_603
timestamp 1682952543
transform 1 0 4048 0 1 370
box -8 -3 104 105
use FILL  FILL_3941
timestamp 1682952543
transform 1 0 4144 0 1 370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_75
timestamp 1682952543
transform 1 0 4177 0 1 370
box -10 -3 10 3
use M2_M1  M2_M1_9208
timestamp 1682952543
transform 1 0 108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9085
timestamp 1682952543
transform 1 0 132 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9209
timestamp 1682952543
transform 1 0 132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9417
timestamp 1682952543
transform 1 0 156 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9386
timestamp 1682952543
transform 1 0 164 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9262
timestamp 1682952543
transform 1 0 196 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9086
timestamp 1682952543
transform 1 0 180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9087
timestamp 1682952543
transform 1 0 188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9210
timestamp 1682952543
transform 1 0 172 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9352
timestamp 1682952543
transform 1 0 204 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9088
timestamp 1682952543
transform 1 0 212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9089
timestamp 1682952543
transform 1 0 220 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9387
timestamp 1682952543
transform 1 0 188 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9211
timestamp 1682952543
transform 1 0 196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9212
timestamp 1682952543
transform 1 0 212 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9388
timestamp 1682952543
transform 1 0 220 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9418
timestamp 1682952543
transform 1 0 212 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9480
timestamp 1682952543
transform 1 0 212 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9353
timestamp 1682952543
transform 1 0 236 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9090
timestamp 1682952543
transform 1 0 244 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9354
timestamp 1682952543
transform 1 0 252 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9091
timestamp 1682952543
transform 1 0 260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9092
timestamp 1682952543
transform 1 0 268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9093
timestamp 1682952543
transform 1 0 284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9213
timestamp 1682952543
transform 1 0 236 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9389
timestamp 1682952543
transform 1 0 244 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9419
timestamp 1682952543
transform 1 0 228 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9355
timestamp 1682952543
transform 1 0 292 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9094
timestamp 1682952543
transform 1 0 300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9214
timestamp 1682952543
transform 1 0 276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9215
timestamp 1682952543
transform 1 0 292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9420
timestamp 1682952543
transform 1 0 284 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9446
timestamp 1682952543
transform 1 0 236 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9447
timestamp 1682952543
transform 1 0 260 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9448
timestamp 1682952543
transform 1 0 276 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9245
timestamp 1682952543
transform 1 0 364 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9263
timestamp 1682952543
transform 1 0 420 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9296
timestamp 1682952543
transform 1 0 332 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9297
timestamp 1682952543
transform 1 0 364 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9246
timestamp 1682952543
transform 1 0 468 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9264
timestamp 1682952543
transform 1 0 500 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9298
timestamp 1682952543
transform 1 0 452 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9265
timestamp 1682952543
transform 1 0 564 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9266
timestamp 1682952543
transform 1 0 596 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9299
timestamp 1682952543
transform 1 0 580 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9300
timestamp 1682952543
transform 1 0 620 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9095
timestamp 1682952543
transform 1 0 332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9096
timestamp 1682952543
transform 1 0 420 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9097
timestamp 1682952543
transform 1 0 428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9098
timestamp 1682952543
transform 1 0 452 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9099
timestamp 1682952543
transform 1 0 468 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9100
timestamp 1682952543
transform 1 0 556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9101
timestamp 1682952543
transform 1 0 580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9102
timestamp 1682952543
transform 1 0 596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9103
timestamp 1682952543
transform 1 0 604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9104
timestamp 1682952543
transform 1 0 620 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9247
timestamp 1682952543
transform 1 0 644 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9105
timestamp 1682952543
transform 1 0 644 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9248
timestamp 1682952543
transform 1 0 844 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9267
timestamp 1682952543
transform 1 0 828 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9268
timestamp 1682952543
transform 1 0 860 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9301
timestamp 1682952543
transform 1 0 740 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9302
timestamp 1682952543
transform 1 0 772 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9106
timestamp 1682952543
transform 1 0 740 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9303
timestamp 1682952543
transform 1 0 836 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9080
timestamp 1682952543
transform 1 0 924 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9107
timestamp 1682952543
transform 1 0 836 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9249
timestamp 1682952543
transform 1 0 972 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9250
timestamp 1682952543
transform 1 0 988 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9269
timestamp 1682952543
transform 1 0 956 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9304
timestamp 1682952543
transform 1 0 940 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9108
timestamp 1682952543
transform 1 0 932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9109
timestamp 1682952543
transform 1 0 948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9216
timestamp 1682952543
transform 1 0 356 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9217
timestamp 1682952543
transform 1 0 412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9218
timestamp 1682952543
transform 1 0 436 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9219
timestamp 1682952543
transform 1 0 452 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9220
timestamp 1682952543
transform 1 0 508 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9221
timestamp 1682952543
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9222
timestamp 1682952543
transform 1 0 556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9223
timestamp 1682952543
transform 1 0 572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9224
timestamp 1682952543
transform 1 0 588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9225
timestamp 1682952543
transform 1 0 612 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9226
timestamp 1682952543
transform 1 0 628 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9227
timestamp 1682952543
transform 1 0 668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9228
timestamp 1682952543
transform 1 0 724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9229
timestamp 1682952543
transform 1 0 764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9230
timestamp 1682952543
transform 1 0 820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9231
timestamp 1682952543
transform 1 0 860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9232
timestamp 1682952543
transform 1 0 916 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9449
timestamp 1682952543
transform 1 0 516 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9508
timestamp 1682952543
transform 1 0 492 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9421
timestamp 1682952543
transform 1 0 604 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9450
timestamp 1682952543
transform 1 0 596 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9509
timestamp 1682952543
transform 1 0 588 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9422
timestamp 1682952543
transform 1 0 676 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9423
timestamp 1682952543
transform 1 0 724 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9451
timestamp 1682952543
transform 1 0 628 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9452
timestamp 1682952543
transform 1 0 724 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9510
timestamp 1682952543
transform 1 0 788 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9453
timestamp 1682952543
transform 1 0 860 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9305
timestamp 1682952543
transform 1 0 972 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9251
timestamp 1682952543
transform 1 0 1020 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9270
timestamp 1682952543
transform 1 0 1004 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9081
timestamp 1682952543
transform 1 0 980 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9110
timestamp 1682952543
transform 1 0 972 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9111
timestamp 1682952543
transform 1 0 988 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9356
timestamp 1682952543
transform 1 0 996 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9306
timestamp 1682952543
transform 1 0 1036 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9112
timestamp 1682952543
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9113
timestamp 1682952543
transform 1 0 1036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9114
timestamp 1682952543
transform 1 0 1044 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9233
timestamp 1682952543
transform 1 0 940 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9234
timestamp 1682952543
transform 1 0 956 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9390
timestamp 1682952543
transform 1 0 980 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9357
timestamp 1682952543
transform 1 0 1060 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9252
timestamp 1682952543
transform 1 0 1076 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9307
timestamp 1682952543
transform 1 0 1076 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9308
timestamp 1682952543
transform 1 0 1092 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9115
timestamp 1682952543
transform 1 0 1068 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9235
timestamp 1682952543
transform 1 0 996 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9236
timestamp 1682952543
transform 1 0 1004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9237
timestamp 1682952543
transform 1 0 1020 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9238
timestamp 1682952543
transform 1 0 1036 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9239
timestamp 1682952543
transform 1 0 1052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9240
timestamp 1682952543
transform 1 0 1068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9343
timestamp 1682952543
transform 1 0 972 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9454
timestamp 1682952543
transform 1 0 956 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9481
timestamp 1682952543
transform 1 0 996 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9455
timestamp 1682952543
transform 1 0 1060 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9116
timestamp 1682952543
transform 1 0 1076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9344
timestamp 1682952543
transform 1 0 1076 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9456
timestamp 1682952543
transform 1 0 1076 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9253
timestamp 1682952543
transform 1 0 1124 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9117
timestamp 1682952543
transform 1 0 1116 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9309
timestamp 1682952543
transform 1 0 1132 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9118
timestamp 1682952543
transform 1 0 1148 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9241
timestamp 1682952543
transform 1 0 1108 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9391
timestamp 1682952543
transform 1 0 1116 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9358
timestamp 1682952543
transform 1 0 1156 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9119
timestamp 1682952543
transform 1 0 1180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9120
timestamp 1682952543
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9242
timestamp 1682952543
transform 1 0 1140 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9243
timestamp 1682952543
transform 1 0 1148 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9345
timestamp 1682952543
transform 1 0 1116 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9346
timestamp 1682952543
transform 1 0 1124 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9511
timestamp 1682952543
transform 1 0 1108 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9424
timestamp 1682952543
transform 1 0 1132 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9244
timestamp 1682952543
transform 1 0 1172 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9392
timestamp 1682952543
transform 1 0 1188 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9310
timestamp 1682952543
transform 1 0 1252 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9311
timestamp 1682952543
transform 1 0 1276 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9121
timestamp 1682952543
transform 1 0 1212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9122
timestamp 1682952543
transform 1 0 1228 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9359
timestamp 1682952543
transform 1 0 1268 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9360
timestamp 1682952543
transform 1 0 1292 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9245
timestamp 1682952543
transform 1 0 1204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9347
timestamp 1682952543
transform 1 0 1156 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9425
timestamp 1682952543
transform 1 0 1180 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9348
timestamp 1682952543
transform 1 0 1188 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9457
timestamp 1682952543
transform 1 0 1148 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9458
timestamp 1682952543
transform 1 0 1172 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9482
timestamp 1682952543
transform 1 0 1124 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9483
timestamp 1682952543
transform 1 0 1156 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9512
timestamp 1682952543
transform 1 0 1140 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9393
timestamp 1682952543
transform 1 0 1212 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9312
timestamp 1682952543
transform 1 0 1348 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9313
timestamp 1682952543
transform 1 0 1364 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9361
timestamp 1682952543
transform 1 0 1324 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9271
timestamp 1682952543
transform 1 0 1412 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9123
timestamp 1682952543
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9124
timestamp 1682952543
transform 1 0 1348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9125
timestamp 1682952543
transform 1 0 1364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9126
timestamp 1682952543
transform 1 0 1372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9246
timestamp 1682952543
transform 1 0 1276 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9459
timestamp 1682952543
transform 1 0 1204 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9484
timestamp 1682952543
transform 1 0 1188 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9513
timestamp 1682952543
transform 1 0 1172 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9394
timestamp 1682952543
transform 1 0 1316 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9485
timestamp 1682952543
transform 1 0 1252 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9247
timestamp 1682952543
transform 1 0 1324 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9248
timestamp 1682952543
transform 1 0 1340 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9249
timestamp 1682952543
transform 1 0 1356 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9460
timestamp 1682952543
transform 1 0 1356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9362
timestamp 1682952543
transform 1 0 1380 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9314
timestamp 1682952543
transform 1 0 1420 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9127
timestamp 1682952543
transform 1 0 1388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9128
timestamp 1682952543
transform 1 0 1412 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9315
timestamp 1682952543
transform 1 0 1516 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9129
timestamp 1682952543
transform 1 0 1436 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9254
timestamp 1682952543
transform 1 0 1604 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9316
timestamp 1682952543
transform 1 0 1580 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9130
timestamp 1682952543
transform 1 0 1548 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9131
timestamp 1682952543
transform 1 0 1556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9132
timestamp 1682952543
transform 1 0 1572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9133
timestamp 1682952543
transform 1 0 1580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9134
timestamp 1682952543
transform 1 0 1604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9250
timestamp 1682952543
transform 1 0 1380 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9251
timestamp 1682952543
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9252
timestamp 1682952543
transform 1 0 1412 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9253
timestamp 1682952543
transform 1 0 1420 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9254
timestamp 1682952543
transform 1 0 1484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9255
timestamp 1682952543
transform 1 0 1516 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9256
timestamp 1682952543
transform 1 0 1524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9257
timestamp 1682952543
transform 1 0 1532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9258
timestamp 1682952543
transform 1 0 1540 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9426
timestamp 1682952543
transform 1 0 1380 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9427
timestamp 1682952543
transform 1 0 1404 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9461
timestamp 1682952543
transform 1 0 1396 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9428
timestamp 1682952543
transform 1 0 1484 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9429
timestamp 1682952543
transform 1 0 1524 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9462
timestamp 1682952543
transform 1 0 1484 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9395
timestamp 1682952543
transform 1 0 1556 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9363
timestamp 1682952543
transform 1 0 1620 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9259
timestamp 1682952543
transform 1 0 1564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9260
timestamp 1682952543
transform 1 0 1580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9261
timestamp 1682952543
transform 1 0 1588 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9262
timestamp 1682952543
transform 1 0 1612 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9430
timestamp 1682952543
transform 1 0 1548 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9486
timestamp 1682952543
transform 1 0 1580 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9272
timestamp 1682952543
transform 1 0 1636 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9317
timestamp 1682952543
transform 1 0 1700 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9318
timestamp 1682952543
transform 1 0 1748 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9364
timestamp 1682952543
transform 1 0 1668 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9135
timestamp 1682952543
transform 1 0 1732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9136
timestamp 1682952543
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9263
timestamp 1682952543
transform 1 0 1652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9264
timestamp 1682952543
transform 1 0 1708 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9265
timestamp 1682952543
transform 1 0 1748 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9431
timestamp 1682952543
transform 1 0 1652 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9432
timestamp 1682952543
transform 1 0 1692 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9433
timestamp 1682952543
transform 1 0 1708 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9434
timestamp 1682952543
transform 1 0 1748 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9487
timestamp 1682952543
transform 1 0 1684 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9488
timestamp 1682952543
transform 1 0 1716 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9319
timestamp 1682952543
transform 1 0 1836 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9273
timestamp 1682952543
transform 1 0 1868 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9274
timestamp 1682952543
transform 1 0 1884 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9320
timestamp 1682952543
transform 1 0 1884 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9137
timestamp 1682952543
transform 1 0 1772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9138
timestamp 1682952543
transform 1 0 1860 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9139
timestamp 1682952543
transform 1 0 1884 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9140
timestamp 1682952543
transform 1 0 1900 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9396
timestamp 1682952543
transform 1 0 1804 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9266
timestamp 1682952543
transform 1 0 1820 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9397
timestamp 1682952543
transform 1 0 1844 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9267
timestamp 1682952543
transform 1 0 1852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9268
timestamp 1682952543
transform 1 0 1860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9269
timestamp 1682952543
transform 1 0 1876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9270
timestamp 1682952543
transform 1 0 1892 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9435
timestamp 1682952543
transform 1 0 1804 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9436
timestamp 1682952543
transform 1 0 1844 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9437
timestamp 1682952543
transform 1 0 1860 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9489
timestamp 1682952543
transform 1 0 1756 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9490
timestamp 1682952543
transform 1 0 1796 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9398
timestamp 1682952543
transform 1 0 1900 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9255
timestamp 1682952543
transform 1 0 1932 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9275
timestamp 1682952543
transform 1 0 1948 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9082
timestamp 1682952543
transform 1 0 1932 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_9321
timestamp 1682952543
transform 1 0 1972 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9256
timestamp 1682952543
transform 1 0 2020 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9276
timestamp 1682952543
transform 1 0 1996 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9322
timestamp 1682952543
transform 1 0 2004 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9141
timestamp 1682952543
transform 1 0 1932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9142
timestamp 1682952543
transform 1 0 1948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9143
timestamp 1682952543
transform 1 0 1956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9144
timestamp 1682952543
transform 1 0 1980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9271
timestamp 1682952543
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9491
timestamp 1682952543
transform 1 0 1892 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9399
timestamp 1682952543
transform 1 0 1924 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9272
timestamp 1682952543
transform 1 0 1948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9349
timestamp 1682952543
transform 1 0 1924 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9514
timestamp 1682952543
transform 1 0 1908 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9400
timestamp 1682952543
transform 1 0 1956 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9365
timestamp 1682952543
transform 1 0 1988 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9273
timestamp 1682952543
transform 1 0 1972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9274
timestamp 1682952543
transform 1 0 1980 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9350
timestamp 1682952543
transform 1 0 1956 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9438
timestamp 1682952543
transform 1 0 1964 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9277
timestamp 1682952543
transform 1 0 2052 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9278
timestamp 1682952543
transform 1 0 2092 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9279
timestamp 1682952543
transform 1 0 2140 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9323
timestamp 1682952543
transform 1 0 2076 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9145
timestamp 1682952543
transform 1 0 2012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9146
timestamp 1682952543
transform 1 0 2020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9147
timestamp 1682952543
transform 1 0 2036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9148
timestamp 1682952543
transform 1 0 2052 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9149
timestamp 1682952543
transform 1 0 2060 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9150
timestamp 1682952543
transform 1 0 2076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9275
timestamp 1682952543
transform 1 0 2004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9351
timestamp 1682952543
transform 1 0 1988 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9492
timestamp 1682952543
transform 1 0 1956 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9515
timestamp 1682952543
transform 1 0 1956 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9493
timestamp 1682952543
transform 1 0 1988 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9401
timestamp 1682952543
transform 1 0 2012 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9366
timestamp 1682952543
transform 1 0 2084 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9324
timestamp 1682952543
transform 1 0 2132 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9325
timestamp 1682952543
transform 1 0 2180 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9151
timestamp 1682952543
transform 1 0 2092 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9152
timestamp 1682952543
transform 1 0 2180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9276
timestamp 1682952543
transform 1 0 2028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9277
timestamp 1682952543
transform 1 0 2044 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9278
timestamp 1682952543
transform 1 0 2060 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9279
timestamp 1682952543
transform 1 0 2084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9280
timestamp 1682952543
transform 1 0 2100 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9281
timestamp 1682952543
transform 1 0 2132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9494
timestamp 1682952543
transform 1 0 2044 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9495
timestamp 1682952543
transform 1 0 2060 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9516
timestamp 1682952543
transform 1 0 2028 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9402
timestamp 1682952543
transform 1 0 2140 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9496
timestamp 1682952543
transform 1 0 2116 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9326
timestamp 1682952543
transform 1 0 2204 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9327
timestamp 1682952543
transform 1 0 2252 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9153
timestamp 1682952543
transform 1 0 2204 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9367
timestamp 1682952543
transform 1 0 2292 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9328
timestamp 1682952543
transform 1 0 2324 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9154
timestamp 1682952543
transform 1 0 2308 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9155
timestamp 1682952543
transform 1 0 2324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9282
timestamp 1682952543
transform 1 0 2252 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9368
timestamp 1682952543
transform 1 0 2332 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9156
timestamp 1682952543
transform 1 0 2340 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9403
timestamp 1682952543
transform 1 0 2300 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9283
timestamp 1682952543
transform 1 0 2308 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9284
timestamp 1682952543
transform 1 0 2316 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9404
timestamp 1682952543
transform 1 0 2324 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9157
timestamp 1682952543
transform 1 0 2372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9285
timestamp 1682952543
transform 1 0 2332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9286
timestamp 1682952543
transform 1 0 2348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9287
timestamp 1682952543
transform 1 0 2356 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9329
timestamp 1682952543
transform 1 0 2388 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9158
timestamp 1682952543
transform 1 0 2388 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9288
timestamp 1682952543
transform 1 0 2388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9289
timestamp 1682952543
transform 1 0 2404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9352
timestamp 1682952543
transform 1 0 2380 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9497
timestamp 1682952543
transform 1 0 2372 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9463
timestamp 1682952543
transform 1 0 2404 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9159
timestamp 1682952543
transform 1 0 2420 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9369
timestamp 1682952543
transform 1 0 2428 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9160
timestamp 1682952543
transform 1 0 2444 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9290
timestamp 1682952543
transform 1 0 2428 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9291
timestamp 1682952543
transform 1 0 2436 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9464
timestamp 1682952543
transform 1 0 2420 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9405
timestamp 1682952543
transform 1 0 2444 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9280
timestamp 1682952543
transform 1 0 2508 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9257
timestamp 1682952543
transform 1 0 2596 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9330
timestamp 1682952543
transform 1 0 2588 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9161
timestamp 1682952543
transform 1 0 2468 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9162
timestamp 1682952543
transform 1 0 2484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9163
timestamp 1682952543
transform 1 0 2572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9292
timestamp 1682952543
transform 1 0 2452 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9406
timestamp 1682952543
transform 1 0 2468 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9370
timestamp 1682952543
transform 1 0 2580 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9083
timestamp 1682952543
transform 1 0 2604 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9164
timestamp 1682952543
transform 1 0 2588 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9165
timestamp 1682952543
transform 1 0 2596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9166
timestamp 1682952543
transform 1 0 2604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9293
timestamp 1682952543
transform 1 0 2532 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9294
timestamp 1682952543
transform 1 0 2564 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9295
timestamp 1682952543
transform 1 0 2572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9353
timestamp 1682952543
transform 1 0 2468 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9465
timestamp 1682952543
transform 1 0 2452 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9466
timestamp 1682952543
transform 1 0 2532 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9467
timestamp 1682952543
transform 1 0 2572 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9498
timestamp 1682952543
transform 1 0 2468 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9499
timestamp 1682952543
transform 1 0 2484 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9500
timestamp 1682952543
transform 1 0 2548 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9371
timestamp 1682952543
transform 1 0 2612 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9167
timestamp 1682952543
transform 1 0 2628 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9372
timestamp 1682952543
transform 1 0 2636 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9281
timestamp 1682952543
transform 1 0 2668 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9331
timestamp 1682952543
transform 1 0 2692 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9332
timestamp 1682952543
transform 1 0 2716 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9168
timestamp 1682952543
transform 1 0 2644 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9169
timestamp 1682952543
transform 1 0 2652 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9170
timestamp 1682952543
transform 1 0 2668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9296
timestamp 1682952543
transform 1 0 2620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9297
timestamp 1682952543
transform 1 0 2636 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9468
timestamp 1682952543
transform 1 0 2620 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9373
timestamp 1682952543
transform 1 0 2676 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9282
timestamp 1682952543
transform 1 0 2748 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9283
timestamp 1682952543
transform 1 0 2852 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9084
timestamp 1682952543
transform 1 0 2748 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9171
timestamp 1682952543
transform 1 0 2692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9172
timestamp 1682952543
transform 1 0 2700 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9173
timestamp 1682952543
transform 1 0 2716 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9374
timestamp 1682952543
transform 1 0 2732 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9174
timestamp 1682952543
transform 1 0 2740 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9298
timestamp 1682952543
transform 1 0 2660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9299
timestamp 1682952543
transform 1 0 2676 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9300
timestamp 1682952543
transform 1 0 2684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9301
timestamp 1682952543
transform 1 0 2708 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9302
timestamp 1682952543
transform 1 0 2724 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9303
timestamp 1682952543
transform 1 0 2732 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9469
timestamp 1682952543
transform 1 0 2660 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9407
timestamp 1682952543
transform 1 0 2740 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9333
timestamp 1682952543
transform 1 0 2764 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9334
timestamp 1682952543
transform 1 0 2836 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9375
timestamp 1682952543
transform 1 0 2788 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9175
timestamp 1682952543
transform 1 0 2836 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9304
timestamp 1682952543
transform 1 0 2756 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9305
timestamp 1682952543
transform 1 0 2788 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9284
timestamp 1682952543
transform 1 0 2948 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9335
timestamp 1682952543
transform 1 0 2860 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9336
timestamp 1682952543
transform 1 0 2908 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9176
timestamp 1682952543
transform 1 0 2860 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9306
timestamp 1682952543
transform 1 0 2908 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9408
timestamp 1682952543
transform 1 0 2940 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9501
timestamp 1682952543
transform 1 0 2900 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9502
timestamp 1682952543
transform 1 0 2932 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9337
timestamp 1682952543
transform 1 0 2980 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9177
timestamp 1682952543
transform 1 0 2964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9178
timestamp 1682952543
transform 1 0 2980 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9376
timestamp 1682952543
transform 1 0 2988 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9285
timestamp 1682952543
transform 1 0 3020 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9338
timestamp 1682952543
transform 1 0 3028 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9179
timestamp 1682952543
transform 1 0 2996 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9180
timestamp 1682952543
transform 1 0 3004 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9181
timestamp 1682952543
transform 1 0 3020 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9182
timestamp 1682952543
transform 1 0 3036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9183
timestamp 1682952543
transform 1 0 3044 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9307
timestamp 1682952543
transform 1 0 2956 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9308
timestamp 1682952543
transform 1 0 2972 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9309
timestamp 1682952543
transform 1 0 2988 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9409
timestamp 1682952543
transform 1 0 3004 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9310
timestamp 1682952543
transform 1 0 3012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9311
timestamp 1682952543
transform 1 0 3028 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9470
timestamp 1682952543
transform 1 0 3036 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9339
timestamp 1682952543
transform 1 0 3076 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9184
timestamp 1682952543
transform 1 0 3076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9312
timestamp 1682952543
transform 1 0 3052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9313
timestamp 1682952543
transform 1 0 3068 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9314
timestamp 1682952543
transform 1 0 3084 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9471
timestamp 1682952543
transform 1 0 3068 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9286
timestamp 1682952543
transform 1 0 3156 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9287
timestamp 1682952543
transform 1 0 3220 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9288
timestamp 1682952543
transform 1 0 3260 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9185
timestamp 1682952543
transform 1 0 3204 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9315
timestamp 1682952543
transform 1 0 3156 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9340
timestamp 1682952543
transform 1 0 3228 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9341
timestamp 1682952543
transform 1 0 3252 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9342
timestamp 1682952543
transform 1 0 3276 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9289
timestamp 1682952543
transform 1 0 3324 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9290
timestamp 1682952543
transform 1 0 3348 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9186
timestamp 1682952543
transform 1 0 3228 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9377
timestamp 1682952543
transform 1 0 3316 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9343
timestamp 1682952543
transform 1 0 3340 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9187
timestamp 1682952543
transform 1 0 3324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9188
timestamp 1682952543
transform 1 0 3340 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9410
timestamp 1682952543
transform 1 0 3228 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_9411
timestamp 1682952543
transform 1 0 3260 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9316
timestamp 1682952543
transform 1 0 3276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9317
timestamp 1682952543
transform 1 0 3308 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9503
timestamp 1682952543
transform 1 0 3228 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9378
timestamp 1682952543
transform 1 0 3348 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9189
timestamp 1682952543
transform 1 0 3356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9318
timestamp 1682952543
transform 1 0 3332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9319
timestamp 1682952543
transform 1 0 3348 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9344
timestamp 1682952543
transform 1 0 3460 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9190
timestamp 1682952543
transform 1 0 3380 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9191
timestamp 1682952543
transform 1 0 3500 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9379
timestamp 1682952543
transform 1 0 3508 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9320
timestamp 1682952543
transform 1 0 3404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9321
timestamp 1682952543
transform 1 0 3460 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9322
timestamp 1682952543
transform 1 0 3484 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9323
timestamp 1682952543
transform 1 0 3500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9354
timestamp 1682952543
transform 1 0 3468 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9355
timestamp 1682952543
transform 1 0 3484 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9359
timestamp 1682952543
transform 1 0 3476 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_9504
timestamp 1682952543
transform 1 0 3460 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9505
timestamp 1682952543
transform 1 0 3500 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9356
timestamp 1682952543
transform 1 0 3516 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_9380
timestamp 1682952543
transform 1 0 3540 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9291
timestamp 1682952543
transform 1 0 3588 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9192
timestamp 1682952543
transform 1 0 3556 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9193
timestamp 1682952543
transform 1 0 3572 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9381
timestamp 1682952543
transform 1 0 3580 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9194
timestamp 1682952543
transform 1 0 3588 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9324
timestamp 1682952543
transform 1 0 3540 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9412
timestamp 1682952543
transform 1 0 3548 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9325
timestamp 1682952543
transform 1 0 3556 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9326
timestamp 1682952543
transform 1 0 3580 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9327
timestamp 1682952543
transform 1 0 3596 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9357
timestamp 1682952543
transform 1 0 3548 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9360
timestamp 1682952543
transform 1 0 3532 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_9472
timestamp 1682952543
transform 1 0 3548 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9473
timestamp 1682952543
transform 1 0 3580 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9506
timestamp 1682952543
transform 1 0 3556 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9517
timestamp 1682952543
transform 1 0 3532 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_9258
timestamp 1682952543
transform 1 0 3604 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9195
timestamp 1682952543
transform 1 0 3612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9328
timestamp 1682952543
transform 1 0 3604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9196
timestamp 1682952543
transform 1 0 3620 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9259
timestamp 1682952543
transform 1 0 3660 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9292
timestamp 1682952543
transform 1 0 3692 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9345
timestamp 1682952543
transform 1 0 3660 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9346
timestamp 1682952543
transform 1 0 3676 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9197
timestamp 1682952543
transform 1 0 3660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9198
timestamp 1682952543
transform 1 0 3676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9329
timestamp 1682952543
transform 1 0 3644 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9439
timestamp 1682952543
transform 1 0 3628 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9440
timestamp 1682952543
transform 1 0 3644 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9382
timestamp 1682952543
transform 1 0 3684 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9199
timestamp 1682952543
transform 1 0 3692 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9330
timestamp 1682952543
transform 1 0 3668 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9331
timestamp 1682952543
transform 1 0 3684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9358
timestamp 1682952543
transform 1 0 3652 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9361
timestamp 1682952543
transform 1 0 3636 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_9474
timestamp 1682952543
transform 1 0 3652 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9475
timestamp 1682952543
transform 1 0 3684 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9507
timestamp 1682952543
transform 1 0 3668 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_9260
timestamp 1682952543
transform 1 0 3748 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_9347
timestamp 1682952543
transform 1 0 3732 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9348
timestamp 1682952543
transform 1 0 3804 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9200
timestamp 1682952543
transform 1 0 3716 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9332
timestamp 1682952543
transform 1 0 3740 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9441
timestamp 1682952543
transform 1 0 3780 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9293
timestamp 1682952543
transform 1 0 3820 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9383
timestamp 1682952543
transform 1 0 3812 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9333
timestamp 1682952543
transform 1 0 3812 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9442
timestamp 1682952543
transform 1 0 3812 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9476
timestamp 1682952543
transform 1 0 3804 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9261
timestamp 1682952543
transform 1 0 3852 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9334
timestamp 1682952543
transform 1 0 3844 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9477
timestamp 1682952543
transform 1 0 3844 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9201
timestamp 1682952543
transform 1 0 3860 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9384
timestamp 1682952543
transform 1 0 3868 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_9413
timestamp 1682952543
transform 1 0 3860 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9335
timestamp 1682952543
transform 1 0 3868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9336
timestamp 1682952543
transform 1 0 3884 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9294
timestamp 1682952543
transform 1 0 3940 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9295
timestamp 1682952543
transform 1 0 4028 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_9349
timestamp 1682952543
transform 1 0 3908 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9350
timestamp 1682952543
transform 1 0 3924 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_9351
timestamp 1682952543
transform 1 0 3980 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9202
timestamp 1682952543
transform 1 0 3900 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9203
timestamp 1682952543
transform 1 0 3908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9204
timestamp 1682952543
transform 1 0 3924 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9205
timestamp 1682952543
transform 1 0 3940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9206
timestamp 1682952543
transform 1 0 3956 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_9414
timestamp 1682952543
transform 1 0 3900 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9337
timestamp 1682952543
transform 1 0 3916 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9415
timestamp 1682952543
transform 1 0 3924 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9338
timestamp 1682952543
transform 1 0 3932 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9443
timestamp 1682952543
transform 1 0 3932 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9478
timestamp 1682952543
transform 1 0 3908 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9385
timestamp 1682952543
transform 1 0 4036 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9339
timestamp 1682952543
transform 1 0 3980 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9416
timestamp 1682952543
transform 1 0 4044 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9207
timestamp 1682952543
transform 1 0 4068 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9340
timestamp 1682952543
transform 1 0 4052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9341
timestamp 1682952543
transform 1 0 4092 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9342
timestamp 1682952543
transform 1 0 4148 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_9444
timestamp 1682952543
transform 1 0 4028 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_9479
timestamp 1682952543
transform 1 0 3980 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_9445
timestamp 1682952543
transform 1 0 4092 0 1 315
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_76
timestamp 1682952543
transform 1 0 24 0 1 270
box -10 -3 10 3
use FILL  FILL_3900
timestamp 1682952543
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1682952543
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1682952543
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_3903
timestamp 1682952543
transform 1 0 96 0 -1 370
box -8 -3 16 105
use FILL  FILL_3904
timestamp 1682952543
transform 1 0 104 0 -1 370
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1682952543
transform 1 0 112 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_665
timestamp 1682952543
transform -1 0 136 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_666
timestamp 1682952543
transform -1 0 152 0 -1 370
box -9 -3 26 105
use FILL  FILL_3906
timestamp 1682952543
transform 1 0 152 0 -1 370
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1682952543
transform 1 0 160 0 -1 370
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1682952543
transform 1 0 168 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_380
timestamp 1682952543
transform -1 0 216 0 -1 370
box -8 -3 46 105
use FILL  FILL_3909
timestamp 1682952543
transform 1 0 216 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_408
timestamp 1682952543
transform -1 0 264 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_409
timestamp 1682952543
transform 1 0 264 0 -1 370
box -8 -3 46 105
use FILL  FILL_3910
timestamp 1682952543
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1682952543
transform 1 0 312 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_582
timestamp 1682952543
transform 1 0 320 0 -1 370
box -8 -3 104 105
use M3_M2  M3_M2_9518
timestamp 1682952543
transform 1 0 452 0 1 275
box -3 -3 3 3
use AOI22X1  AOI22X1_381
timestamp 1682952543
transform -1 0 456 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_583
timestamp 1682952543
transform 1 0 456 0 -1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_382
timestamp 1682952543
transform -1 0 592 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_383
timestamp 1682952543
transform -1 0 632 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_9519
timestamp 1682952543
transform 1 0 724 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_584
timestamp 1682952543
transform 1 0 632 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_585
timestamp 1682952543
transform 1 0 728 0 -1 370
box -8 -3 104 105
use M3_M2  M3_M2_9520
timestamp 1682952543
transform 1 0 916 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_586
timestamp 1682952543
transform 1 0 824 0 -1 370
box -8 -3 104 105
use NOR2X1  NOR2X1_110
timestamp 1682952543
transform 1 0 920 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_168
timestamp 1682952543
transform 1 0 944 0 -1 370
box -8 -3 34 105
use NOR2X1  NOR2X1_111
timestamp 1682952543
transform 1 0 976 0 -1 370
box -8 -3 32 105
use AOI22X1  AOI22X1_384
timestamp 1682952543
transform 1 0 1000 0 -1 370
box -8 -3 46 105
use OAI21X1  OAI21X1_169
timestamp 1682952543
transform 1 0 1040 0 -1 370
box -8 -3 34 105
use FILL  FILL_3912
timestamp 1682952543
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_170
timestamp 1682952543
transform 1 0 1080 0 -1 370
box -8 -3 34 105
use FILL  FILL_3913
timestamp 1682952543
transform 1 0 1112 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_171
timestamp 1682952543
transform -1 0 1152 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_172
timestamp 1682952543
transform -1 0 1184 0 -1 370
box -8 -3 34 105
use OAI21X1  OAI21X1_173
timestamp 1682952543
transform -1 0 1216 0 -1 370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_587
timestamp 1682952543
transform 1 0 1216 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_667
timestamp 1682952543
transform 1 0 1312 0 -1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_410
timestamp 1682952543
transform -1 0 1368 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_9521
timestamp 1682952543
transform 1 0 1396 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_411
timestamp 1682952543
transform -1 0 1408 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_668
timestamp 1682952543
transform 1 0 1408 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_588
timestamp 1682952543
transform 1 0 1424 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_669
timestamp 1682952543
transform -1 0 1536 0 -1 370
box -9 -3 26 105
use FILL  FILL_3914
timestamp 1682952543
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_9522
timestamp 1682952543
transform 1 0 1588 0 1 275
box -3 -3 3 3
use AOI22X1  AOI22X1_385
timestamp 1682952543
transform -1 0 1584 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_412
timestamp 1682952543
transform 1 0 1584 0 -1 370
box -8 -3 46 105
use FILL  FILL_3915
timestamp 1682952543
transform 1 0 1624 0 -1 370
box -8 -3 16 105
use FILL  FILL_3916
timestamp 1682952543
transform 1 0 1632 0 -1 370
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1682952543
transform 1 0 1640 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_9523
timestamp 1682952543
transform 1 0 1740 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_589
timestamp 1682952543
transform -1 0 1744 0 -1 370
box -8 -3 104 105
use M3_M2  M3_M2_9524
timestamp 1682952543
transform 1 0 1756 0 1 275
box -3 -3 3 3
use INVX2  INVX2_670
timestamp 1682952543
transform 1 0 1744 0 -1 370
box -9 -3 26 105
use M3_M2  M3_M2_9525
timestamp 1682952543
transform 1 0 1828 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_9526
timestamp 1682952543
transform 1 0 1844 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_590
timestamp 1682952543
transform 1 0 1760 0 -1 370
box -8 -3 104 105
use AOI22X1  AOI22X1_386
timestamp 1682952543
transform -1 0 1896 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_9527
timestamp 1682952543
transform 1 0 1916 0 1 275
box -3 -3 3 3
use OAI21X1  OAI21X1_174
timestamp 1682952543
transform 1 0 1896 0 -1 370
box -8 -3 34 105
use NOR2X1  NOR2X1_112
timestamp 1682952543
transform 1 0 1928 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_175
timestamp 1682952543
transform -1 0 1984 0 -1 370
box -8 -3 34 105
use M3_M2  M3_M2_9528
timestamp 1682952543
transform 1 0 2004 0 1 275
box -3 -3 3 3
use OAI21X1  OAI21X1_176
timestamp 1682952543
transform -1 0 2016 0 -1 370
box -8 -3 34 105
use M3_M2  M3_M2_9529
timestamp 1682952543
transform 1 0 2060 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_413
timestamp 1682952543
transform 1 0 2016 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_414
timestamp 1682952543
transform 1 0 2056 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_591
timestamp 1682952543
transform -1 0 2192 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_592
timestamp 1682952543
transform 1 0 2192 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_671
timestamp 1682952543
transform 1 0 2288 0 -1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_415
timestamp 1682952543
transform 1 0 2304 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_9530
timestamp 1682952543
transform 1 0 2356 0 1 275
box -3 -3 3 3
use OAI21X1  OAI21X1_177
timestamp 1682952543
transform 1 0 2344 0 -1 370
box -8 -3 34 105
use FILL  FILL_3918
timestamp 1682952543
transform 1 0 2376 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_178
timestamp 1682952543
transform -1 0 2416 0 -1 370
box -8 -3 34 105
use FILL  FILL_3919
timestamp 1682952543
transform 1 0 2416 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_672
timestamp 1682952543
transform 1 0 2424 0 -1 370
box -9 -3 26 105
use OAI21X1  OAI21X1_179
timestamp 1682952543
transform 1 0 2440 0 -1 370
box -8 -3 34 105
use M3_M2  M3_M2_9531
timestamp 1682952543
transform 1 0 2508 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_593
timestamp 1682952543
transform 1 0 2472 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_673
timestamp 1682952543
transform 1 0 2568 0 -1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_113
timestamp 1682952543
transform -1 0 2608 0 -1 370
box -8 -3 32 105
use OAI22X1  OAI22X1_416
timestamp 1682952543
transform -1 0 2648 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_417
timestamp 1682952543
transform -1 0 2688 0 -1 370
box -8 -3 46 105
use AOI22X1  AOI22X1_387
timestamp 1682952543
transform 1 0 2688 0 -1 370
box -8 -3 46 105
use NOR2X1  NOR2X1_114
timestamp 1682952543
transform -1 0 2752 0 -1 370
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_594
timestamp 1682952543
transform -1 0 2848 0 -1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_595
timestamp 1682952543
transform 1 0 2848 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_674
timestamp 1682952543
transform 1 0 2944 0 -1 370
box -9 -3 26 105
use OAI22X1  OAI22X1_418
timestamp 1682952543
transform -1 0 3000 0 -1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_419
timestamp 1682952543
transform 1 0 3000 0 -1 370
box -8 -3 46 105
use FILL  FILL_3920
timestamp 1682952543
transform 1 0 3040 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_388
timestamp 1682952543
transform -1 0 3088 0 -1 370
box -8 -3 46 105
use FILL  FILL_3921
timestamp 1682952543
transform 1 0 3088 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_675
timestamp 1682952543
transform -1 0 3112 0 -1 370
box -9 -3 26 105
use FILL  FILL_3922
timestamp 1682952543
transform 1 0 3112 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_9532
timestamp 1682952543
transform 1 0 3188 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_596
timestamp 1682952543
transform -1 0 3216 0 -1 370
box -8 -3 104 105
use M3_M2  M3_M2_9533
timestamp 1682952543
transform 1 0 3284 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_597
timestamp 1682952543
transform 1 0 3216 0 -1 370
box -8 -3 104 105
use FILL  FILL_3923
timestamp 1682952543
transform 1 0 3312 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_9534
timestamp 1682952543
transform 1 0 3356 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_420
timestamp 1682952543
transform -1 0 3360 0 -1 370
box -8 -3 46 105
use FILL  FILL_3924
timestamp 1682952543
transform 1 0 3360 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_600
timestamp 1682952543
transform 1 0 3368 0 -1 370
box -8 -3 104 105
use NAND3X1  NAND3X1_75
timestamp 1682952543
transform -1 0 3496 0 -1 370
box -8 -3 40 105
use INVX2  INVX2_677
timestamp 1682952543
transform 1 0 3496 0 -1 370
box -9 -3 26 105
use FILL  FILL_3930
timestamp 1682952543
transform 1 0 3512 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_76
timestamp 1682952543
transform -1 0 3552 0 -1 370
box -8 -3 40 105
use M3_M2  M3_M2_9535
timestamp 1682952543
transform 1 0 3564 0 1 275
box -3 -3 3 3
use OAI22X1  OAI22X1_423
timestamp 1682952543
transform 1 0 3552 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_678
timestamp 1682952543
transform -1 0 3608 0 -1 370
box -9 -3 26 105
use FILL  FILL_3931
timestamp 1682952543
transform 1 0 3608 0 -1 370
box -8 -3 16 105
use FILL  FILL_3932
timestamp 1682952543
transform 1 0 3616 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_77
timestamp 1682952543
transform -1 0 3656 0 -1 370
box -8 -3 40 105
use OAI22X1  OAI22X1_424
timestamp 1682952543
transform 1 0 3656 0 -1 370
box -8 -3 46 105
use FILL  FILL_3942
timestamp 1682952543
transform 1 0 3696 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_604
timestamp 1682952543
transform 1 0 3704 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_680
timestamp 1682952543
transform 1 0 3800 0 -1 370
box -9 -3 26 105
use FILL  FILL_3943
timestamp 1682952543
transform 1 0 3816 0 -1 370
box -8 -3 16 105
use FILL  FILL_3944
timestamp 1682952543
transform 1 0 3824 0 -1 370
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1682952543
transform 1 0 3832 0 -1 370
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1682952543
transform 1 0 3840 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_389
timestamp 1682952543
transform -1 0 3888 0 -1 370
box -8 -3 46 105
use M3_M2  M3_M2_9536
timestamp 1682952543
transform 1 0 3900 0 1 275
box -3 -3 3 3
use FILL  FILL_3947
timestamp 1682952543
transform 1 0 3888 0 -1 370
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1682952543
transform 1 0 3896 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_427
timestamp 1682952543
transform 1 0 3904 0 -1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_605
timestamp 1682952543
transform 1 0 3944 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_681
timestamp 1682952543
transform 1 0 4040 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_606
timestamp 1682952543
transform 1 0 4056 0 -1 370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_77
timestamp 1682952543
transform 1 0 4201 0 1 270
box -10 -3 10 3
use M2_M1  M2_M1_9370
timestamp 1682952543
transform 1 0 132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9371
timestamp 1682952543
transform 1 0 164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9372
timestamp 1682952543
transform 1 0 172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9553
timestamp 1682952543
transform 1 0 84 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9797
timestamp 1682952543
transform 1 0 76 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9537
timestamp 1682952543
transform 1 0 284 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9639
timestamp 1682952543
transform 1 0 252 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9373
timestamp 1682952543
transform 1 0 212 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9677
timestamp 1682952543
transform 1 0 220 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9374
timestamp 1682952543
transform 1 0 228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9375
timestamp 1682952543
transform 1 0 252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9376
timestamp 1682952543
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9554
timestamp 1682952543
transform 1 0 212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9555
timestamp 1682952543
transform 1 0 220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9556
timestamp 1682952543
transform 1 0 236 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9798
timestamp 1682952543
transform 1 0 236 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9678
timestamp 1682952543
transform 1 0 276 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9377
timestamp 1682952543
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9557
timestamp 1682952543
transform 1 0 260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9558
timestamp 1682952543
transform 1 0 276 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9640
timestamp 1682952543
transform 1 0 316 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9378
timestamp 1682952543
transform 1 0 316 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9379
timestamp 1682952543
transform 1 0 356 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9679
timestamp 1682952543
transform 1 0 364 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9566
timestamp 1682952543
transform 1 0 380 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9380
timestamp 1682952543
transform 1 0 380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9559
timestamp 1682952543
transform 1 0 348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9560
timestamp 1682952543
transform 1 0 364 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9561
timestamp 1682952543
transform 1 0 372 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9748
timestamp 1682952543
transform 1 0 348 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9749
timestamp 1682952543
transform 1 0 372 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9588
timestamp 1682952543
transform 1 0 412 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9604
timestamp 1682952543
transform 1 0 428 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9567
timestamp 1682952543
transform 1 0 452 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9641
timestamp 1682952543
transform 1 0 444 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9381
timestamp 1682952543
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9382
timestamp 1682952543
transform 1 0 428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9562
timestamp 1682952543
transform 1 0 420 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9721
timestamp 1682952543
transform 1 0 428 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9383
timestamp 1682952543
transform 1 0 444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9563
timestamp 1682952543
transform 1 0 436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9384
timestamp 1682952543
transform 1 0 468 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9680
timestamp 1682952543
transform 1 0 476 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9568
timestamp 1682952543
transform 1 0 524 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9589
timestamp 1682952543
transform 1 0 508 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9605
timestamp 1682952543
transform 1 0 532 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9385
timestamp 1682952543
transform 1 0 492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9386
timestamp 1682952543
transform 1 0 500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9387
timestamp 1682952543
transform 1 0 508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9388
timestamp 1682952543
transform 1 0 532 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9681
timestamp 1682952543
transform 1 0 540 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9564
timestamp 1682952543
transform 1 0 460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9565
timestamp 1682952543
transform 1 0 476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9566
timestamp 1682952543
transform 1 0 484 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9567
timestamp 1682952543
transform 1 0 508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9568
timestamp 1682952543
transform 1 0 524 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9750
timestamp 1682952543
transform 1 0 460 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9751
timestamp 1682952543
transform 1 0 508 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9752
timestamp 1682952543
transform 1 0 532 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9569
timestamp 1682952543
transform 1 0 548 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9642
timestamp 1682952543
transform 1 0 580 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9590
timestamp 1682952543
transform 1 0 636 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9606
timestamp 1682952543
transform 1 0 628 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9643
timestamp 1682952543
transform 1 0 612 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9389
timestamp 1682952543
transform 1 0 588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9390
timestamp 1682952543
transform 1 0 596 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9682
timestamp 1682952543
transform 1 0 604 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9644
timestamp 1682952543
transform 1 0 636 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9391
timestamp 1682952543
transform 1 0 612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9392
timestamp 1682952543
transform 1 0 628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9393
timestamp 1682952543
transform 1 0 636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9570
timestamp 1682952543
transform 1 0 580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9571
timestamp 1682952543
transform 1 0 604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9394
timestamp 1682952543
transform 1 0 668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9572
timestamp 1682952543
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9573
timestamp 1682952543
transform 1 0 660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9574
timestamp 1682952543
transform 1 0 676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9575
timestamp 1682952543
transform 1 0 684 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9395
timestamp 1682952543
transform 1 0 692 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9722
timestamp 1682952543
transform 1 0 700 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_9591
timestamp 1682952543
transform 1 0 772 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9607
timestamp 1682952543
transform 1 0 764 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9396
timestamp 1682952543
transform 1 0 716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9397
timestamp 1682952543
transform 1 0 724 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9683
timestamp 1682952543
transform 1 0 732 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9362
timestamp 1682952543
transform 1 0 788 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9398
timestamp 1682952543
transform 1 0 740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9399
timestamp 1682952543
transform 1 0 764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9400
timestamp 1682952543
transform 1 0 772 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9576
timestamp 1682952543
transform 1 0 708 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9753
timestamp 1682952543
transform 1 0 668 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9754
timestamp 1682952543
transform 1 0 684 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9735
timestamp 1682952543
transform 1 0 700 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_9799
timestamp 1682952543
transform 1 0 660 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9723
timestamp 1682952543
transform 1 0 716 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9577
timestamp 1682952543
transform 1 0 732 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9578
timestamp 1682952543
transform 1 0 748 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9755
timestamp 1682952543
transform 1 0 740 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9592
timestamp 1682952543
transform 1 0 852 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9608
timestamp 1682952543
transform 1 0 844 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9401
timestamp 1682952543
transform 1 0 796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9402
timestamp 1682952543
transform 1 0 804 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9724
timestamp 1682952543
transform 1 0 780 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9579
timestamp 1682952543
transform 1 0 788 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9684
timestamp 1682952543
transform 1 0 820 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9403
timestamp 1682952543
transform 1 0 828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9404
timestamp 1682952543
transform 1 0 844 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9405
timestamp 1682952543
transform 1 0 852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9580
timestamp 1682952543
transform 1 0 812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9581
timestamp 1682952543
transform 1 0 820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9582
timestamp 1682952543
transform 1 0 852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9363
timestamp 1682952543
transform 1 0 876 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_9725
timestamp 1682952543
transform 1 0 876 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_9569
timestamp 1682952543
transform 1 0 924 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9609
timestamp 1682952543
transform 1 0 908 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9593
timestamp 1682952543
transform 1 0 932 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9594
timestamp 1682952543
transform 1 0 964 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9610
timestamp 1682952543
transform 1 0 956 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9406
timestamp 1682952543
transform 1 0 900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9407
timestamp 1682952543
transform 1 0 908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9408
timestamp 1682952543
transform 1 0 916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9583
timestamp 1682952543
transform 1 0 884 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9584
timestamp 1682952543
transform 1 0 892 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9756
timestamp 1682952543
transform 1 0 868 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9685
timestamp 1682952543
transform 1 0 932 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9409
timestamp 1682952543
transform 1 0 940 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9410
timestamp 1682952543
transform 1 0 956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9585
timestamp 1682952543
transform 1 0 924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9586
timestamp 1682952543
transform 1 0 932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9587
timestamp 1682952543
transform 1 0 948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9588
timestamp 1682952543
transform 1 0 956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9736
timestamp 1682952543
transform 1 0 884 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_9757
timestamp 1682952543
transform 1 0 892 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9800
timestamp 1682952543
transform 1 0 884 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9686
timestamp 1682952543
transform 1 0 972 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9538
timestamp 1682952543
transform 1 0 1004 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9570
timestamp 1682952543
transform 1 0 1012 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9595
timestamp 1682952543
transform 1 0 1020 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9611
timestamp 1682952543
transform 1 0 1028 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9411
timestamp 1682952543
transform 1 0 1004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9412
timestamp 1682952543
transform 1 0 1012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9413
timestamp 1682952543
transform 1 0 1028 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9589
timestamp 1682952543
transform 1 0 996 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9758
timestamp 1682952543
transform 1 0 996 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9539
timestamp 1682952543
transform 1 0 1060 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9612
timestamp 1682952543
transform 1 0 1052 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9364
timestamp 1682952543
transform 1 0 1052 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_9687
timestamp 1682952543
transform 1 0 1052 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9590
timestamp 1682952543
transform 1 0 1020 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9591
timestamp 1682952543
transform 1 0 1044 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9592
timestamp 1682952543
transform 1 0 1052 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9759
timestamp 1682952543
transform 1 0 1028 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9613
timestamp 1682952543
transform 1 0 1092 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9614
timestamp 1682952543
transform 1 0 1116 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9365
timestamp 1682952543
transform 1 0 1068 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_9688
timestamp 1682952543
transform 1 0 1068 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9366
timestamp 1682952543
transform 1 0 1100 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9414
timestamp 1682952543
transform 1 0 1092 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9689
timestamp 1682952543
transform 1 0 1100 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9615
timestamp 1682952543
transform 1 0 1140 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9415
timestamp 1682952543
transform 1 0 1116 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9690
timestamp 1682952543
transform 1 0 1124 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9416
timestamp 1682952543
transform 1 0 1140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9593
timestamp 1682952543
transform 1 0 1092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9594
timestamp 1682952543
transform 1 0 1100 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9726
timestamp 1682952543
transform 1 0 1108 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9595
timestamp 1682952543
transform 1 0 1124 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9596
timestamp 1682952543
transform 1 0 1132 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9760
timestamp 1682952543
transform 1 0 1092 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9761
timestamp 1682952543
transform 1 0 1140 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9801
timestamp 1682952543
transform 1 0 1124 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9571
timestamp 1682952543
transform 1 0 1188 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9691
timestamp 1682952543
transform 1 0 1164 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9572
timestamp 1682952543
transform 1 0 1236 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9616
timestamp 1682952543
transform 1 0 1228 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9417
timestamp 1682952543
transform 1 0 1172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9418
timestamp 1682952543
transform 1 0 1196 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9692
timestamp 1682952543
transform 1 0 1204 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9419
timestamp 1682952543
transform 1 0 1212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9420
timestamp 1682952543
transform 1 0 1228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9421
timestamp 1682952543
transform 1 0 1244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9597
timestamp 1682952543
transform 1 0 1164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9598
timestamp 1682952543
transform 1 0 1180 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9599
timestamp 1682952543
transform 1 0 1196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9600
timestamp 1682952543
transform 1 0 1204 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9601
timestamp 1682952543
transform 1 0 1220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9602
timestamp 1682952543
transform 1 0 1236 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9762
timestamp 1682952543
transform 1 0 1172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9763
timestamp 1682952543
transform 1 0 1188 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9802
timestamp 1682952543
transform 1 0 1212 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9803
timestamp 1682952543
transform 1 0 1244 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9617
timestamp 1682952543
transform 1 0 1284 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9693
timestamp 1682952543
transform 1 0 1260 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9540
timestamp 1682952543
transform 1 0 1308 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9573
timestamp 1682952543
transform 1 0 1396 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9596
timestamp 1682952543
transform 1 0 1356 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9618
timestamp 1682952543
transform 1 0 1356 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9619
timestamp 1682952543
transform 1 0 1388 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9422
timestamp 1682952543
transform 1 0 1268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9423
timestamp 1682952543
transform 1 0 1284 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9694
timestamp 1682952543
transform 1 0 1292 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9424
timestamp 1682952543
transform 1 0 1356 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9603
timestamp 1682952543
transform 1 0 1252 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9604
timestamp 1682952543
transform 1 0 1260 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9605
timestamp 1682952543
transform 1 0 1276 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9727
timestamp 1682952543
transform 1 0 1284 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9606
timestamp 1682952543
transform 1 0 1292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9607
timestamp 1682952543
transform 1 0 1308 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9425
timestamp 1682952543
transform 1 0 1404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9426
timestamp 1682952543
transform 1 0 1412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9608
timestamp 1682952543
transform 1 0 1412 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9764
timestamp 1682952543
transform 1 0 1412 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9427
timestamp 1682952543
transform 1 0 1436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9428
timestamp 1682952543
transform 1 0 1444 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9728
timestamp 1682952543
transform 1 0 1436 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_9620
timestamp 1682952543
transform 1 0 1468 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9429
timestamp 1682952543
transform 1 0 1452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9430
timestamp 1682952543
transform 1 0 1476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9609
timestamp 1682952543
transform 1 0 1460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9610
timestamp 1682952543
transform 1 0 1468 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9765
timestamp 1682952543
transform 1 0 1484 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9611
timestamp 1682952543
transform 1 0 1500 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9766
timestamp 1682952543
transform 1 0 1500 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9574
timestamp 1682952543
transform 1 0 1532 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9541
timestamp 1682952543
transform 1 0 1548 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9575
timestamp 1682952543
transform 1 0 1588 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9621
timestamp 1682952543
transform 1 0 1564 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9645
timestamp 1682952543
transform 1 0 1580 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9542
timestamp 1682952543
transform 1 0 1612 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9622
timestamp 1682952543
transform 1 0 1604 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9431
timestamp 1682952543
transform 1 0 1532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9432
timestamp 1682952543
transform 1 0 1540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9433
timestamp 1682952543
transform 1 0 1548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9434
timestamp 1682952543
transform 1 0 1572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9435
timestamp 1682952543
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9436
timestamp 1682952543
transform 1 0 1596 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9612
timestamp 1682952543
transform 1 0 1556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9613
timestamp 1682952543
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9614
timestamp 1682952543
transform 1 0 1580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9615
timestamp 1682952543
transform 1 0 1588 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9767
timestamp 1682952543
transform 1 0 1588 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9804
timestamp 1682952543
transform 1 0 1580 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9623
timestamp 1682952543
transform 1 0 1644 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9624
timestamp 1682952543
transform 1 0 1684 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9437
timestamp 1682952543
transform 1 0 1628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9438
timestamp 1682952543
transform 1 0 1644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9439
timestamp 1682952543
transform 1 0 1660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9440
timestamp 1682952543
transform 1 0 1684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9441
timestamp 1682952543
transform 1 0 1700 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9695
timestamp 1682952543
transform 1 0 1708 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9442
timestamp 1682952543
transform 1 0 1716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9616
timestamp 1682952543
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9617
timestamp 1682952543
transform 1 0 1644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9618
timestamp 1682952543
transform 1 0 1668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9619
timestamp 1682952543
transform 1 0 1684 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9620
timestamp 1682952543
transform 1 0 1692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9621
timestamp 1682952543
transform 1 0 1708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9622
timestamp 1682952543
transform 1 0 1716 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9768
timestamp 1682952543
transform 1 0 1668 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9769
timestamp 1682952543
transform 1 0 1708 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9805
timestamp 1682952543
transform 1 0 1716 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9543
timestamp 1682952543
transform 1 0 1764 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9544
timestamp 1682952543
transform 1 0 1788 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9545
timestamp 1682952543
transform 1 0 1812 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9576
timestamp 1682952543
transform 1 0 1748 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9577
timestamp 1682952543
transform 1 0 1780 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9625
timestamp 1682952543
transform 1 0 1780 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9626
timestamp 1682952543
transform 1 0 1804 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9443
timestamp 1682952543
transform 1 0 1740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9444
timestamp 1682952543
transform 1 0 1764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9445
timestamp 1682952543
transform 1 0 1780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9446
timestamp 1682952543
transform 1 0 1796 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9696
timestamp 1682952543
transform 1 0 1804 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9546
timestamp 1682952543
transform 1 0 1868 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9447
timestamp 1682952543
transform 1 0 1812 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9448
timestamp 1682952543
transform 1 0 1820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9449
timestamp 1682952543
transform 1 0 1828 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9623
timestamp 1682952543
transform 1 0 1756 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9624
timestamp 1682952543
transform 1 0 1772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9625
timestamp 1682952543
transform 1 0 1804 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9770
timestamp 1682952543
transform 1 0 1740 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9771
timestamp 1682952543
transform 1 0 1772 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9806
timestamp 1682952543
transform 1 0 1796 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9697
timestamp 1682952543
transform 1 0 1844 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9547
timestamp 1682952543
transform 1 0 1908 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9450
timestamp 1682952543
transform 1 0 1852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9451
timestamp 1682952543
transform 1 0 1868 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9698
timestamp 1682952543
transform 1 0 1884 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9548
timestamp 1682952543
transform 1 0 1948 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9549
timestamp 1682952543
transform 1 0 1964 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9452
timestamp 1682952543
transform 1 0 1892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9453
timestamp 1682952543
transform 1 0 1908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9454
timestamp 1682952543
transform 1 0 1916 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9699
timestamp 1682952543
transform 1 0 1924 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9455
timestamp 1682952543
transform 1 0 1932 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9700
timestamp 1682952543
transform 1 0 1940 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9456
timestamp 1682952543
transform 1 0 1948 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9457
timestamp 1682952543
transform 1 0 1956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9626
timestamp 1682952543
transform 1 0 1836 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9627
timestamp 1682952543
transform 1 0 1844 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9628
timestamp 1682952543
transform 1 0 1860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9629
timestamp 1682952543
transform 1 0 1876 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9630
timestamp 1682952543
transform 1 0 1884 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9631
timestamp 1682952543
transform 1 0 1916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9632
timestamp 1682952543
transform 1 0 1924 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9633
timestamp 1682952543
transform 1 0 1940 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9634
timestamp 1682952543
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9807
timestamp 1682952543
transform 1 0 1836 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9772
timestamp 1682952543
transform 1 0 1916 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9773
timestamp 1682952543
transform 1 0 1948 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9808
timestamp 1682952543
transform 1 0 1932 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9367
timestamp 1682952543
transform 1 0 1980 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_9550
timestamp 1682952543
transform 1 0 2020 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9458
timestamp 1682952543
transform 1 0 2004 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9701
timestamp 1682952543
transform 1 0 2012 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9597
timestamp 1682952543
transform 1 0 2052 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9598
timestamp 1682952543
transform 1 0 2076 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9368
timestamp 1682952543
transform 1 0 2044 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_9646
timestamp 1682952543
transform 1 0 2068 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9459
timestamp 1682952543
transform 1 0 2020 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9702
timestamp 1682952543
transform 1 0 2044 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9460
timestamp 1682952543
transform 1 0 2060 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9703
timestamp 1682952543
transform 1 0 2076 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9635
timestamp 1682952543
transform 1 0 1988 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9636
timestamp 1682952543
transform 1 0 2004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9637
timestamp 1682952543
transform 1 0 2012 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9638
timestamp 1682952543
transform 1 0 2036 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9737
timestamp 1682952543
transform 1 0 1988 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_9774
timestamp 1682952543
transform 1 0 2036 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9809
timestamp 1682952543
transform 1 0 2020 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9551
timestamp 1682952543
transform 1 0 2092 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9647
timestamp 1682952543
transform 1 0 2116 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9552
timestamp 1682952543
transform 1 0 2148 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9553
timestamp 1682952543
transform 1 0 2188 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9648
timestamp 1682952543
transform 1 0 2156 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9461
timestamp 1682952543
transform 1 0 2092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9462
timestamp 1682952543
transform 1 0 2100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9463
timestamp 1682952543
transform 1 0 2116 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9464
timestamp 1682952543
transform 1 0 2140 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9465
timestamp 1682952543
transform 1 0 2156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9639
timestamp 1682952543
transform 1 0 2076 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9640
timestamp 1682952543
transform 1 0 2084 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9738
timestamp 1682952543
transform 1 0 2076 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_9810
timestamp 1682952543
transform 1 0 2052 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9704
timestamp 1682952543
transform 1 0 2172 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9466
timestamp 1682952543
transform 1 0 2180 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9554
timestamp 1682952543
transform 1 0 2292 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9555
timestamp 1682952543
transform 1 0 2316 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9649
timestamp 1682952543
transform 1 0 2308 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9467
timestamp 1682952543
transform 1 0 2228 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9705
timestamp 1682952543
transform 1 0 2292 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9468
timestamp 1682952543
transform 1 0 2300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9469
timestamp 1682952543
transform 1 0 2308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9470
timestamp 1682952543
transform 1 0 2332 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9471
timestamp 1682952543
transform 1 0 2348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9641
timestamp 1682952543
transform 1 0 2108 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9642
timestamp 1682952543
transform 1 0 2116 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9643
timestamp 1682952543
transform 1 0 2132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9644
timestamp 1682952543
transform 1 0 2148 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9645
timestamp 1682952543
transform 1 0 2156 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9646
timestamp 1682952543
transform 1 0 2172 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9647
timestamp 1682952543
transform 1 0 2188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9648
timestamp 1682952543
transform 1 0 2204 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9775
timestamp 1682952543
transform 1 0 2092 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9811
timestamp 1682952543
transform 1 0 2100 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9812
timestamp 1682952543
transform 1 0 2116 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9776
timestamp 1682952543
transform 1 0 2172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9813
timestamp 1682952543
transform 1 0 2148 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9777
timestamp 1682952543
transform 1 0 2228 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9814
timestamp 1682952543
transform 1 0 2204 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9729
timestamp 1682952543
transform 1 0 2300 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9649
timestamp 1682952543
transform 1 0 2308 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9730
timestamp 1682952543
transform 1 0 2316 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9650
timestamp 1682952543
transform 1 0 2324 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9731
timestamp 1682952543
transform 1 0 2332 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9651
timestamp 1682952543
transform 1 0 2340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9652
timestamp 1682952543
transform 1 0 2348 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9556
timestamp 1682952543
transform 1 0 2404 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9369
timestamp 1682952543
transform 1 0 2388 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_9650
timestamp 1682952543
transform 1 0 2396 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9472
timestamp 1682952543
transform 1 0 2372 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9651
timestamp 1682952543
transform 1 0 2452 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9652
timestamp 1682952543
transform 1 0 2476 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9473
timestamp 1682952543
transform 1 0 2396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9474
timestamp 1682952543
transform 1 0 2412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9653
timestamp 1682952543
transform 1 0 2388 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9706
timestamp 1682952543
transform 1 0 2420 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9475
timestamp 1682952543
transform 1 0 2428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9476
timestamp 1682952543
transform 1 0 2444 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9477
timestamp 1682952543
transform 1 0 2468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9478
timestamp 1682952543
transform 1 0 2492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9479
timestamp 1682952543
transform 1 0 2500 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9654
timestamp 1682952543
transform 1 0 2412 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9655
timestamp 1682952543
transform 1 0 2420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9656
timestamp 1682952543
transform 1 0 2436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9657
timestamp 1682952543
transform 1 0 2444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9658
timestamp 1682952543
transform 1 0 2460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9659
timestamp 1682952543
transform 1 0 2476 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9660
timestamp 1682952543
transform 1 0 2484 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9778
timestamp 1682952543
transform 1 0 2412 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9779
timestamp 1682952543
transform 1 0 2428 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9780
timestamp 1682952543
transform 1 0 2492 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9815
timestamp 1682952543
transform 1 0 2420 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9816
timestamp 1682952543
transform 1 0 2452 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9653
timestamp 1682952543
transform 1 0 2540 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9661
timestamp 1682952543
transform 1 0 2540 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9627
timestamp 1682952543
transform 1 0 2556 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9662
timestamp 1682952543
transform 1 0 2556 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9557
timestamp 1682952543
transform 1 0 2620 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9578
timestamp 1682952543
transform 1 0 2612 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9654
timestamp 1682952543
transform 1 0 2588 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9480
timestamp 1682952543
transform 1 0 2564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9481
timestamp 1682952543
transform 1 0 2572 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9707
timestamp 1682952543
transform 1 0 2580 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9628
timestamp 1682952543
transform 1 0 2636 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9655
timestamp 1682952543
transform 1 0 2644 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9482
timestamp 1682952543
transform 1 0 2588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9483
timestamp 1682952543
transform 1 0 2612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9484
timestamp 1682952543
transform 1 0 2628 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9663
timestamp 1682952543
transform 1 0 2596 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9664
timestamp 1682952543
transform 1 0 2612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9665
timestamp 1682952543
transform 1 0 2620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9666
timestamp 1682952543
transform 1 0 2636 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9667
timestamp 1682952543
transform 1 0 2644 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9629
timestamp 1682952543
transform 1 0 2660 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9485
timestamp 1682952543
transform 1 0 2660 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9781
timestamp 1682952543
transform 1 0 2660 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9630
timestamp 1682952543
transform 1 0 2684 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9486
timestamp 1682952543
transform 1 0 2684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9487
timestamp 1682952543
transform 1 0 2692 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9732
timestamp 1682952543
transform 1 0 2692 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_9656
timestamp 1682952543
transform 1 0 2724 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9708
timestamp 1682952543
transform 1 0 2708 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9657
timestamp 1682952543
transform 1 0 2756 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9658
timestamp 1682952543
transform 1 0 2796 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9488
timestamp 1682952543
transform 1 0 2716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9489
timestamp 1682952543
transform 1 0 2732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9668
timestamp 1682952543
transform 1 0 2700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9669
timestamp 1682952543
transform 1 0 2724 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9782
timestamp 1682952543
transform 1 0 2724 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9709
timestamp 1682952543
transform 1 0 2740 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9490
timestamp 1682952543
transform 1 0 2756 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9491
timestamp 1682952543
transform 1 0 2764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9492
timestamp 1682952543
transform 1 0 2796 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9670
timestamp 1682952543
transform 1 0 2740 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9733
timestamp 1682952543
transform 1 0 2812 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9671
timestamp 1682952543
transform 1 0 2844 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9783
timestamp 1682952543
transform 1 0 2756 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9659
timestamp 1682952543
transform 1 0 2876 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9493
timestamp 1682952543
transform 1 0 2876 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9494
timestamp 1682952543
transform 1 0 2892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9495
timestamp 1682952543
transform 1 0 2908 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9672
timestamp 1682952543
transform 1 0 2868 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9673
timestamp 1682952543
transform 1 0 2884 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9734
timestamp 1682952543
transform 1 0 2892 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9674
timestamp 1682952543
transform 1 0 2900 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9784
timestamp 1682952543
transform 1 0 2868 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9817
timestamp 1682952543
transform 1 0 2900 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9675
timestamp 1682952543
transform 1 0 2916 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9558
timestamp 1682952543
transform 1 0 2964 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9631
timestamp 1682952543
transform 1 0 2980 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9632
timestamp 1682952543
transform 1 0 3004 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9660
timestamp 1682952543
transform 1 0 2972 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9496
timestamp 1682952543
transform 1 0 2932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9497
timestamp 1682952543
transform 1 0 2948 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9498
timestamp 1682952543
transform 1 0 2964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9499
timestamp 1682952543
transform 1 0 2972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9500
timestamp 1682952543
transform 1 0 3004 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9633
timestamp 1682952543
transform 1 0 3020 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9501
timestamp 1682952543
transform 1 0 3020 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9676
timestamp 1682952543
transform 1 0 2972 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9677
timestamp 1682952543
transform 1 0 2980 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9678
timestamp 1682952543
transform 1 0 2996 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9679
timestamp 1682952543
transform 1 0 3012 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9680
timestamp 1682952543
transform 1 0 3020 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9785
timestamp 1682952543
transform 1 0 2988 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9710
timestamp 1682952543
transform 1 0 3028 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9786
timestamp 1682952543
transform 1 0 3020 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9818
timestamp 1682952543
transform 1 0 3012 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9579
timestamp 1682952543
transform 1 0 3068 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9711
timestamp 1682952543
transform 1 0 3052 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9502
timestamp 1682952543
transform 1 0 3060 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9559
timestamp 1682952543
transform 1 0 3084 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9503
timestamp 1682952543
transform 1 0 3076 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9681
timestamp 1682952543
transform 1 0 3052 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9682
timestamp 1682952543
transform 1 0 3068 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9787
timestamp 1682952543
transform 1 0 3052 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9504
timestamp 1682952543
transform 1 0 3116 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9712
timestamp 1682952543
transform 1 0 3132 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9683
timestamp 1682952543
transform 1 0 3164 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9788
timestamp 1682952543
transform 1 0 3116 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9789
timestamp 1682952543
transform 1 0 3148 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9819
timestamp 1682952543
transform 1 0 3132 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9820
timestamp 1682952543
transform 1 0 3164 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9661
timestamp 1682952543
transform 1 0 3180 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9505
timestamp 1682952543
transform 1 0 3180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9506
timestamp 1682952543
transform 1 0 3212 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9713
timestamp 1682952543
transform 1 0 3220 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9560
timestamp 1682952543
transform 1 0 3260 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9634
timestamp 1682952543
transform 1 0 3276 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9662
timestamp 1682952543
transform 1 0 3268 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9507
timestamp 1682952543
transform 1 0 3228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9508
timestamp 1682952543
transform 1 0 3244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9509
timestamp 1682952543
transform 1 0 3260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9684
timestamp 1682952543
transform 1 0 3188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9685
timestamp 1682952543
transform 1 0 3204 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9686
timestamp 1682952543
transform 1 0 3220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9687
timestamp 1682952543
transform 1 0 3228 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9790
timestamp 1682952543
transform 1 0 3204 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9821
timestamp 1682952543
transform 1 0 3196 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9822
timestamp 1682952543
transform 1 0 3220 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9580
timestamp 1682952543
transform 1 0 3308 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9663
timestamp 1682952543
transform 1 0 3300 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9510
timestamp 1682952543
transform 1 0 3276 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9511
timestamp 1682952543
transform 1 0 3300 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9635
timestamp 1682952543
transform 1 0 3324 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9664
timestamp 1682952543
transform 1 0 3316 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9688
timestamp 1682952543
transform 1 0 3268 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9689
timestamp 1682952543
transform 1 0 3276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9690
timestamp 1682952543
transform 1 0 3292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9691
timestamp 1682952543
transform 1 0 3308 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9512
timestamp 1682952543
transform 1 0 3324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9513
timestamp 1682952543
transform 1 0 3364 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9714
timestamp 1682952543
transform 1 0 3372 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9514
timestamp 1682952543
transform 1 0 3380 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9692
timestamp 1682952543
transform 1 0 3324 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9693
timestamp 1682952543
transform 1 0 3340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9694
timestamp 1682952543
transform 1 0 3356 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9735
timestamp 1682952543
transform 1 0 3364 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9695
timestamp 1682952543
transform 1 0 3372 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9696
timestamp 1682952543
transform 1 0 3380 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9823
timestamp 1682952543
transform 1 0 3332 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9824
timestamp 1682952543
transform 1 0 3348 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9561
timestamp 1682952543
transform 1 0 3412 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9515
timestamp 1682952543
transform 1 0 3412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9516
timestamp 1682952543
transform 1 0 3428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9697
timestamp 1682952543
transform 1 0 3404 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9698
timestamp 1682952543
transform 1 0 3420 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9825
timestamp 1682952543
transform 1 0 3380 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_9736
timestamp 1682952543
transform 1 0 3428 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_9791
timestamp 1682952543
transform 1 0 3420 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9699
timestamp 1682952543
transform 1 0 3444 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9581
timestamp 1682952543
transform 1 0 3460 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9517
timestamp 1682952543
transform 1 0 3460 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9599
timestamp 1682952543
transform 1 0 3476 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9636
timestamp 1682952543
transform 1 0 3492 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9518
timestamp 1682952543
transform 1 0 3484 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9715
timestamp 1682952543
transform 1 0 3500 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9737
timestamp 1682952543
transform 1 0 3484 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9700
timestamp 1682952543
transform 1 0 3492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9701
timestamp 1682952543
transform 1 0 3500 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9562
timestamp 1682952543
transform 1 0 3516 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9563
timestamp 1682952543
transform 1 0 3564 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9582
timestamp 1682952543
transform 1 0 3596 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9600
timestamp 1682952543
transform 1 0 3564 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9665
timestamp 1682952543
transform 1 0 3532 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9519
timestamp 1682952543
transform 1 0 3524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9520
timestamp 1682952543
transform 1 0 3532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9521
timestamp 1682952543
transform 1 0 3548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9702
timestamp 1682952543
transform 1 0 3516 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9792
timestamp 1682952543
transform 1 0 3508 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9716
timestamp 1682952543
transform 1 0 3556 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9522
timestamp 1682952543
transform 1 0 3564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9523
timestamp 1682952543
transform 1 0 3580 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9524
timestamp 1682952543
transform 1 0 3596 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9738
timestamp 1682952543
transform 1 0 3532 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9703
timestamp 1682952543
transform 1 0 3540 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9704
timestamp 1682952543
transform 1 0 3556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9705
timestamp 1682952543
transform 1 0 3564 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9666
timestamp 1682952543
transform 1 0 3612 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9525
timestamp 1682952543
transform 1 0 3612 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9526
timestamp 1682952543
transform 1 0 3636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9527
timestamp 1682952543
transform 1 0 3652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9706
timestamp 1682952543
transform 1 0 3604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9707
timestamp 1682952543
transform 1 0 3612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9708
timestamp 1682952543
transform 1 0 3628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9739
timestamp 1682952543
transform 1 0 3636 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9709
timestamp 1682952543
transform 1 0 3644 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9583
timestamp 1682952543
transform 1 0 3668 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9584
timestamp 1682952543
transform 1 0 3692 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9585
timestamp 1682952543
transform 1 0 3708 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9601
timestamp 1682952543
transform 1 0 3700 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9602
timestamp 1682952543
transform 1 0 3764 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9667
timestamp 1682952543
transform 1 0 3716 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9668
timestamp 1682952543
transform 1 0 3740 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9528
timestamp 1682952543
transform 1 0 3660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9529
timestamp 1682952543
transform 1 0 3668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9530
timestamp 1682952543
transform 1 0 3684 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9531
timestamp 1682952543
transform 1 0 3700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9532
timestamp 1682952543
transform 1 0 3716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9710
timestamp 1682952543
transform 1 0 3668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9711
timestamp 1682952543
transform 1 0 3676 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9740
timestamp 1682952543
transform 1 0 3692 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_9717
timestamp 1682952543
transform 1 0 3724 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9669
timestamp 1682952543
transform 1 0 3788 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9586
timestamp 1682952543
transform 1 0 3836 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9603
timestamp 1682952543
transform 1 0 3836 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_9637
timestamp 1682952543
transform 1 0 3820 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9670
timestamp 1682952543
transform 1 0 3828 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9533
timestamp 1682952543
transform 1 0 3732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9534
timestamp 1682952543
transform 1 0 3740 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9535
timestamp 1682952543
transform 1 0 3764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9536
timestamp 1682952543
transform 1 0 3780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9537
timestamp 1682952543
transform 1 0 3804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9538
timestamp 1682952543
transform 1 0 3820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9712
timestamp 1682952543
transform 1 0 3700 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9713
timestamp 1682952543
transform 1 0 3708 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9714
timestamp 1682952543
transform 1 0 3724 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9715
timestamp 1682952543
transform 1 0 3740 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9741
timestamp 1682952543
transform 1 0 3748 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9716
timestamp 1682952543
transform 1 0 3764 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9717
timestamp 1682952543
transform 1 0 3772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9718
timestamp 1682952543
transform 1 0 3788 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9793
timestamp 1682952543
transform 1 0 3772 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9718
timestamp 1682952543
transform 1 0 3828 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_9564
timestamp 1682952543
transform 1 0 3876 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9587
timestamp 1682952543
transform 1 0 3884 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_9671
timestamp 1682952543
transform 1 0 3852 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9539
timestamp 1682952543
transform 1 0 3836 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9540
timestamp 1682952543
transform 1 0 3852 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9541
timestamp 1682952543
transform 1 0 3868 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9542
timestamp 1682952543
transform 1 0 3884 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9565
timestamp 1682952543
transform 1 0 3908 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_9672
timestamp 1682952543
transform 1 0 3892 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9673
timestamp 1682952543
transform 1 0 3924 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_9638
timestamp 1682952543
transform 1 0 3964 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_9674
timestamp 1682952543
transform 1 0 3972 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9543
timestamp 1682952543
transform 1 0 3892 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9544
timestamp 1682952543
transform 1 0 3924 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9719
timestamp 1682952543
transform 1 0 3812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9720
timestamp 1682952543
transform 1 0 3828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9721
timestamp 1682952543
transform 1 0 3844 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9742
timestamp 1682952543
transform 1 0 3852 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9722
timestamp 1682952543
transform 1 0 3860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9723
timestamp 1682952543
transform 1 0 3876 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9743
timestamp 1682952543
transform 1 0 3884 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_9719
timestamp 1682952543
transform 1 0 3940 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9545
timestamp 1682952543
transform 1 0 3948 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9546
timestamp 1682952543
transform 1 0 3964 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9547
timestamp 1682952543
transform 1 0 3972 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9724
timestamp 1682952543
transform 1 0 3892 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9725
timestamp 1682952543
transform 1 0 3900 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9794
timestamp 1682952543
transform 1 0 3868 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9744
timestamp 1682952543
transform 1 0 3908 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9726
timestamp 1682952543
transform 1 0 3916 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9745
timestamp 1682952543
transform 1 0 3924 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9727
timestamp 1682952543
transform 1 0 3932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9728
timestamp 1682952543
transform 1 0 3956 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9729
timestamp 1682952543
transform 1 0 3972 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9795
timestamp 1682952543
transform 1 0 3900 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9826
timestamp 1682952543
transform 1 0 3972 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9548
timestamp 1682952543
transform 1 0 3996 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9675
timestamp 1682952543
transform 1 0 4036 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9549
timestamp 1682952543
transform 1 0 4036 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_9720
timestamp 1682952543
transform 1 0 4044 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9550
timestamp 1682952543
transform 1 0 4052 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9730
timestamp 1682952543
transform 1 0 4004 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9731
timestamp 1682952543
transform 1 0 4012 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9746
timestamp 1682952543
transform 1 0 4020 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9732
timestamp 1682952543
transform 1 0 4028 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9747
timestamp 1682952543
transform 1 0 4036 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9733
timestamp 1682952543
transform 1 0 4044 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_9796
timestamp 1682952543
transform 1 0 4012 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_9676
timestamp 1682952543
transform 1 0 4084 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9551
timestamp 1682952543
transform 1 0 4084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9734
timestamp 1682952543
transform 1 0 4084 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9552
timestamp 1682952543
transform 1 0 4148 0 1 215
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_78
timestamp 1682952543
transform 1 0 48 0 1 170
box -10 -3 10 3
use M3_M2  M3_M2_9827
timestamp 1682952543
transform 1 0 132 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_9828
timestamp 1682952543
transform 1 0 172 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_607
timestamp 1682952543
transform 1 0 72 0 1 170
box -8 -3 104 105
use INVX2  INVX2_682
timestamp 1682952543
transform -1 0 184 0 1 170
box -9 -3 26 105
use FILL  FILL_3949
timestamp 1682952543
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1682952543
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1682952543
transform 1 0 200 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_390
timestamp 1682952543
transform 1 0 208 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_391
timestamp 1682952543
transform -1 0 288 0 1 170
box -8 -3 46 105
use FILL  FILL_3952
timestamp 1682952543
transform 1 0 288 0 1 170
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1682952543
transform 1 0 296 0 1 170
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1682952543
transform 1 0 304 0 1 170
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1682952543
transform 1 0 312 0 1 170
box -8 -3 16 105
use FILL  FILL_3961
timestamp 1682952543
transform 1 0 320 0 1 170
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1682952543
transform 1 0 328 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_392
timestamp 1682952543
transform -1 0 376 0 1 170
box -8 -3 46 105
use FILL  FILL_3964
timestamp 1682952543
transform 1 0 376 0 1 170
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1682952543
transform 1 0 384 0 1 170
box -8 -3 16 105
use FILL  FILL_3966
timestamp 1682952543
transform 1 0 392 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_428
timestamp 1682952543
transform 1 0 400 0 1 170
box -8 -3 46 105
use FILL  FILL_3967
timestamp 1682952543
transform 1 0 440 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_393
timestamp 1682952543
transform -1 0 488 0 1 170
box -8 -3 46 105
use INVX2  INVX2_684
timestamp 1682952543
transform 1 0 488 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_429
timestamp 1682952543
transform 1 0 504 0 1 170
box -8 -3 46 105
use FILL  FILL_3968
timestamp 1682952543
transform 1 0 544 0 1 170
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1682952543
transform 1 0 552 0 1 170
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1682952543
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1682952543
transform 1 0 568 0 1 170
box -8 -3 16 105
use INVX2  INVX2_685
timestamp 1682952543
transform 1 0 576 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_394
timestamp 1682952543
transform 1 0 592 0 1 170
box -8 -3 46 105
use FILL  FILL_3972
timestamp 1682952543
transform 1 0 632 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9829
timestamp 1682952543
transform 1 0 668 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_430
timestamp 1682952543
transform 1 0 640 0 1 170
box -8 -3 46 105
use INVX2  INVX2_686
timestamp 1682952543
transform 1 0 680 0 1 170
box -9 -3 26 105
use NOR2X1  NOR2X1_115
timestamp 1682952543
transform 1 0 696 0 1 170
box -8 -3 32 105
use AOI22X1  AOI22X1_395
timestamp 1682952543
transform 1 0 720 0 1 170
box -8 -3 46 105
use OAI21X1  OAI21X1_180
timestamp 1682952543
transform 1 0 760 0 1 170
box -8 -3 34 105
use INVX2  INVX2_687
timestamp 1682952543
transform -1 0 808 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_396
timestamp 1682952543
transform 1 0 808 0 1 170
box -8 -3 46 105
use OAI21X1  OAI21X1_181
timestamp 1682952543
transform 1 0 848 0 1 170
box -8 -3 34 105
use NOR2X1  NOR2X1_116
timestamp 1682952543
transform 1 0 880 0 1 170
box -8 -3 32 105
use INVX2  INVX2_688
timestamp 1682952543
transform -1 0 920 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_397
timestamp 1682952543
transform 1 0 920 0 1 170
box -8 -3 46 105
use FILL  FILL_3973
timestamp 1682952543
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1682952543
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1682952543
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1682952543
transform 1 0 984 0 1 170
box -8 -3 16 105
use INVX2  INVX2_690
timestamp 1682952543
transform 1 0 992 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_398
timestamp 1682952543
transform 1 0 1008 0 1 170
box -8 -3 46 105
use FILL  FILL_3983
timestamp 1682952543
transform 1 0 1048 0 1 170
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1682952543
transform 1 0 1056 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_182
timestamp 1682952543
transform -1 0 1096 0 1 170
box -8 -3 34 105
use OAI21X1  OAI21X1_183
timestamp 1682952543
transform -1 0 1128 0 1 170
box -8 -3 34 105
use INVX2  INVX2_691
timestamp 1682952543
transform 1 0 1128 0 1 170
box -9 -3 26 105
use FILL  FILL_3985
timestamp 1682952543
transform 1 0 1144 0 1 170
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1682952543
transform 1 0 1152 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9830
timestamp 1682952543
transform 1 0 1172 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_431
timestamp 1682952543
transform -1 0 1200 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_432
timestamp 1682952543
transform -1 0 1240 0 1 170
box -8 -3 46 105
use INVX2  INVX2_692
timestamp 1682952543
transform -1 0 1256 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_433
timestamp 1682952543
transform -1 0 1296 0 1 170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_616
timestamp 1682952543
transform 1 0 1296 0 1 170
box -8 -3 104 105
use INVX2  INVX2_693
timestamp 1682952543
transform 1 0 1392 0 1 170
box -9 -3 26 105
use FILL  FILL_3987
timestamp 1682952543
transform 1 0 1408 0 1 170
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1682952543
transform 1 0 1416 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9831
timestamp 1682952543
transform 1 0 1452 0 1 175
box -3 -3 3 3
use INVX2  INVX2_694
timestamp 1682952543
transform 1 0 1424 0 1 170
box -9 -3 26 105
use INVX2  INVX2_695
timestamp 1682952543
transform -1 0 1456 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_399
timestamp 1682952543
transform 1 0 1456 0 1 170
box -8 -3 46 105
use FILL  FILL_3989
timestamp 1682952543
transform 1 0 1496 0 1 170
box -8 -3 16 105
use FILL  FILL_3990
timestamp 1682952543
transform 1 0 1504 0 1 170
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1682952543
transform 1 0 1512 0 1 170
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1682952543
transform 1 0 1520 0 1 170
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1682952543
transform 1 0 1528 0 1 170
box -8 -3 16 105
use INVX2  INVX2_696
timestamp 1682952543
transform -1 0 1552 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_400
timestamp 1682952543
transform 1 0 1552 0 1 170
box -8 -3 46 105
use FILL  FILL_3994
timestamp 1682952543
transform 1 0 1592 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9832
timestamp 1682952543
transform 1 0 1620 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_434
timestamp 1682952543
transform 1 0 1600 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_401
timestamp 1682952543
transform -1 0 1680 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_402
timestamp 1682952543
transform -1 0 1720 0 1 170
box -8 -3 46 105
use FILL  FILL_3995
timestamp 1682952543
transform 1 0 1720 0 1 170
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1682952543
transform 1 0 1728 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9833
timestamp 1682952543
transform 1 0 1756 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_435
timestamp 1682952543
transform 1 0 1736 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_403
timestamp 1682952543
transform -1 0 1816 0 1 170
box -8 -3 46 105
use INVX2  INVX2_697
timestamp 1682952543
transform -1 0 1832 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_404
timestamp 1682952543
transform 1 0 1832 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_405
timestamp 1682952543
transform 1 0 1872 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_406
timestamp 1682952543
transform 1 0 1912 0 1 170
box -8 -3 46 105
use OAI21X1  OAI21X1_184
timestamp 1682952543
transform 1 0 1952 0 1 170
box -8 -3 34 105
use NOR2X1  NOR2X1_117
timestamp 1682952543
transform 1 0 1984 0 1 170
box -8 -3 32 105
use OAI21X1  OAI21X1_185
timestamp 1682952543
transform 1 0 2008 0 1 170
box -8 -3 34 105
use M3_M2  M3_M2_9834
timestamp 1682952543
transform 1 0 2076 0 1 175
box -3 -3 3 3
use OAI21X1  OAI21X1_186
timestamp 1682952543
transform -1 0 2072 0 1 170
box -8 -3 34 105
use NOR2X1  NOR2X1_118
timestamp 1682952543
transform 1 0 2072 0 1 170
box -8 -3 32 105
use INVX2  INVX2_698
timestamp 1682952543
transform -1 0 2112 0 1 170
box -9 -3 26 105
use M3_M2  M3_M2_9835
timestamp 1682952543
transform 1 0 2140 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_436
timestamp 1682952543
transform 1 0 2112 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_437
timestamp 1682952543
transform 1 0 2152 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_9836
timestamp 1682952543
transform 1 0 2244 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_617
timestamp 1682952543
transform 1 0 2192 0 1 170
box -8 -3 104 105
use INVX2  INVX2_699
timestamp 1682952543
transform 1 0 2288 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_438
timestamp 1682952543
transform 1 0 2304 0 1 170
box -8 -3 46 105
use INVX2  INVX2_700
timestamp 1682952543
transform 1 0 2344 0 1 170
box -9 -3 26 105
use OAI21X1  OAI21X1_187
timestamp 1682952543
transform 1 0 2360 0 1 170
box -8 -3 34 105
use INVX2  INVX2_701
timestamp 1682952543
transform -1 0 2408 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_407
timestamp 1682952543
transform 1 0 2408 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_408
timestamp 1682952543
transform -1 0 2488 0 1 170
box -8 -3 46 105
use INVX2  INVX2_702
timestamp 1682952543
transform 1 0 2488 0 1 170
box -9 -3 26 105
use FILL  FILL_3997
timestamp 1682952543
transform 1 0 2504 0 1 170
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1682952543
transform 1 0 2512 0 1 170
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1682952543
transform 1 0 2520 0 1 170
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1682952543
transform 1 0 2528 0 1 170
box -8 -3 16 105
use INVX2  INVX2_703
timestamp 1682952543
transform 1 0 2536 0 1 170
box -9 -3 26 105
use FILL  FILL_4001
timestamp 1682952543
transform 1 0 2552 0 1 170
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1682952543
transform 1 0 2560 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_409
timestamp 1682952543
transform 1 0 2568 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_410
timestamp 1682952543
transform -1 0 2648 0 1 170
box -8 -3 46 105
use FILL  FILL_4003
timestamp 1682952543
transform 1 0 2648 0 1 170
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1682952543
transform 1 0 2656 0 1 170
box -8 -3 16 105
use INVX2  INVX2_704
timestamp 1682952543
transform 1 0 2664 0 1 170
box -9 -3 26 105
use FILL  FILL_4005
timestamp 1682952543
transform 1 0 2680 0 1 170
box -8 -3 16 105
use FILL  FILL_4006
timestamp 1682952543
transform 1 0 2688 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_411
timestamp 1682952543
transform 1 0 2696 0 1 170
box -8 -3 46 105
use FILL  FILL_4007
timestamp 1682952543
transform 1 0 2736 0 1 170
box -8 -3 16 105
use INVX2  INVX2_705
timestamp 1682952543
transform 1 0 2744 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_618
timestamp 1682952543
transform -1 0 2856 0 1 170
box -8 -3 104 105
use FILL  FILL_4008
timestamp 1682952543
transform 1 0 2856 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_439
timestamp 1682952543
transform 1 0 2864 0 1 170
box -8 -3 46 105
use INVX2  INVX2_706
timestamp 1682952543
transform -1 0 2920 0 1 170
box -9 -3 26 105
use FILL  FILL_4009
timestamp 1682952543
transform 1 0 2920 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9837
timestamp 1682952543
transform 1 0 2972 0 1 175
box -3 -3 3 3
use AOI22X1  AOI22X1_412
timestamp 1682952543
transform -1 0 2968 0 1 170
box -8 -3 46 105
use FILL  FILL_4010
timestamp 1682952543
transform 1 0 2968 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_440
timestamp 1682952543
transform 1 0 2976 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_9838
timestamp 1682952543
transform 1 0 3028 0 1 175
box -3 -3 3 3
use FILL  FILL_4011
timestamp 1682952543
transform 1 0 3016 0 1 170
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1682952543
transform 1 0 3024 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9839
timestamp 1682952543
transform 1 0 3068 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_441
timestamp 1682952543
transform 1 0 3032 0 1 170
box -8 -3 46 105
use FILL  FILL_4013
timestamp 1682952543
transform 1 0 3072 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_619
timestamp 1682952543
transform -1 0 3176 0 1 170
box -8 -3 104 105
use M3_M2  M3_M2_9840
timestamp 1682952543
transform 1 0 3188 0 1 175
box -3 -3 3 3
use FILL  FILL_4014
timestamp 1682952543
transform 1 0 3176 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_442
timestamp 1682952543
transform 1 0 3184 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_413
timestamp 1682952543
transform -1 0 3264 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_9841
timestamp 1682952543
transform 1 0 3276 0 1 175
box -3 -3 3 3
use FILL  FILL_4015
timestamp 1682952543
transform 1 0 3264 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_443
timestamp 1682952543
transform 1 0 3272 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_9842
timestamp 1682952543
transform 1 0 3324 0 1 175
box -3 -3 3 3
use FILL  FILL_4016
timestamp 1682952543
transform 1 0 3312 0 1 170
box -8 -3 16 105
use INVX2  INVX2_707
timestamp 1682952543
transform 1 0 3320 0 1 170
box -9 -3 26 105
use M3_M2  M3_M2_9843
timestamp 1682952543
transform 1 0 3372 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_444
timestamp 1682952543
transform 1 0 3336 0 1 170
box -8 -3 46 105
use FILL  FILL_4017
timestamp 1682952543
transform 1 0 3376 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_445
timestamp 1682952543
transform 1 0 3384 0 1 170
box -8 -3 46 105
use INVX2  INVX2_708
timestamp 1682952543
transform -1 0 3440 0 1 170
box -9 -3 26 105
use FILL  FILL_4018
timestamp 1682952543
transform 1 0 3440 0 1 170
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1682952543
transform 1 0 3448 0 1 170
box -8 -3 16 105
use FILL  FILL_4042
timestamp 1682952543
transform 1 0 3456 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_414
timestamp 1682952543
transform -1 0 3504 0 1 170
box -8 -3 46 105
use FILL  FILL_4043
timestamp 1682952543
transform 1 0 3504 0 1 170
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1682952543
transform 1 0 3512 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_9844
timestamp 1682952543
transform 1 0 3532 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_446
timestamp 1682952543
transform 1 0 3520 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_415
timestamp 1682952543
transform 1 0 3560 0 1 170
box -8 -3 46 105
use FILL  FILL_4045
timestamp 1682952543
transform 1 0 3600 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_447
timestamp 1682952543
transform 1 0 3608 0 1 170
box -8 -3 46 105
use INVX2  INVX2_721
timestamp 1682952543
transform -1 0 3664 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_416
timestamp 1682952543
transform -1 0 3704 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_448
timestamp 1682952543
transform -1 0 3744 0 1 170
box -8 -3 46 105
use INVX2  INVX2_722
timestamp 1682952543
transform -1 0 3760 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_417
timestamp 1682952543
transform 1 0 3760 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_418
timestamp 1682952543
transform -1 0 3840 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_449
timestamp 1682952543
transform 1 0 3840 0 1 170
box -8 -3 46 105
use INVX2  INVX2_723
timestamp 1682952543
transform -1 0 3896 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_450
timestamp 1682952543
transform 1 0 3896 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_451
timestamp 1682952543
transform -1 0 3976 0 1 170
box -8 -3 46 105
use INVX2  INVX2_724
timestamp 1682952543
transform -1 0 3992 0 1 170
box -9 -3 26 105
use FILL  FILL_4046
timestamp 1682952543
transform 1 0 3992 0 1 170
box -8 -3 16 105
use FILL  FILL_4047
timestamp 1682952543
transform 1 0 4000 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_452
timestamp 1682952543
transform 1 0 4008 0 1 170
box -8 -3 46 105
use FILL  FILL_4048
timestamp 1682952543
transform 1 0 4048 0 1 170
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1682952543
transform 1 0 4056 0 1 170
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1682952543
transform 1 0 4064 0 1 170
box -8 -3 16 105
use INVX2  INVX2_725
timestamp 1682952543
transform -1 0 4088 0 1 170
box -9 -3 26 105
use INVX2  INVX2_726
timestamp 1682952543
transform -1 0 4104 0 1 170
box -9 -3 26 105
use FILL  FILL_4051
timestamp 1682952543
transform 1 0 4104 0 1 170
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1682952543
transform 1 0 4112 0 1 170
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1682952543
transform 1 0 4120 0 1 170
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1682952543
transform 1 0 4128 0 1 170
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1682952543
transform 1 0 4136 0 1 170
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1682952543
transform 1 0 4144 0 1 170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_79
timestamp 1682952543
transform 1 0 4177 0 1 170
box -10 -3 10 3
use M3_M2  M3_M2_9878
timestamp 1682952543
transform 1 0 156 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9739
timestamp 1682952543
transform 1 0 156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9783
timestamp 1682952543
transform 1 0 76 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9784
timestamp 1682952543
transform 1 0 132 0 1 125
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_80
timestamp 1682952543
transform 1 0 24 0 1 70
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_608
timestamp 1682952543
transform -1 0 168 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9879
timestamp 1682952543
transform 1 0 180 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_9880
timestamp 1682952543
transform 1 0 204 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9740
timestamp 1682952543
transform 1 0 180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9741
timestamp 1682952543
transform 1 0 268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9785
timestamp 1682952543
transform 1 0 228 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9786
timestamp 1682952543
transform 1 0 260 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9787
timestamp 1682952543
transform 1 0 268 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9925
timestamp 1682952543
transform 1 0 228 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9926
timestamp 1682952543
transform 1 0 268 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_609
timestamp 1682952543
transform 1 0 168 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_683
timestamp 1682952543
transform 1 0 264 0 -1 170
box -9 -3 26 105
use FILL  FILL_3953
timestamp 1682952543
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1682952543
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1682952543
transform 1 0 296 0 -1 170
box -8 -3 16 105
use FILL  FILL_3958
timestamp 1682952543
transform 1 0 304 0 -1 170
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1682952543
transform 1 0 312 0 -1 170
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1682952543
transform 1 0 320 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9742
timestamp 1682952543
transform 1 0 340 0 1 135
box -2 -2 2 2
use FILL  FILL_3974
timestamp 1682952543
transform 1 0 328 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9881
timestamp 1682952543
transform 1 0 436 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9743
timestamp 1682952543
transform 1 0 436 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9788
timestamp 1682952543
transform 1 0 348 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9789
timestamp 1682952543
transform 1 0 356 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9790
timestamp 1682952543
transform 1 0 388 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9927
timestamp 1682952543
transform 1 0 348 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9928
timestamp 1682952543
transform 1 0 388 0 1 115
box -3 -3 3 3
use INVX2  INVX2_689
timestamp 1682952543
transform 1 0 336 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_610
timestamp 1682952543
transform -1 0 448 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9882
timestamp 1682952543
transform 1 0 540 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9744
timestamp 1682952543
transform 1 0 540 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9791
timestamp 1682952543
transform 1 0 460 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9792
timestamp 1682952543
transform 1 0 500 0 1 125
box -2 -2 2 2
use FILL  FILL_3975
timestamp 1682952543
transform 1 0 448 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9929
timestamp 1682952543
transform 1 0 516 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_611
timestamp 1682952543
transform -1 0 552 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9845
timestamp 1682952543
transform 1 0 596 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9883
timestamp 1682952543
transform 1 0 564 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9745
timestamp 1682952543
transform 1 0 564 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9793
timestamp 1682952543
transform 1 0 588 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9794
timestamp 1682952543
transform 1 0 644 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_612
timestamp 1682952543
transform 1 0 552 0 -1 170
box -8 -3 104 105
use FILL  FILL_3976
timestamp 1682952543
transform 1 0 648 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9884
timestamp 1682952543
transform 1 0 668 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9746
timestamp 1682952543
transform 1 0 668 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9795
timestamp 1682952543
transform 1 0 692 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9796
timestamp 1682952543
transform 1 0 748 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_613
timestamp 1682952543
transform 1 0 656 0 -1 170
box -8 -3 104 105
use FILL  FILL_3977
timestamp 1682952543
transform 1 0 752 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9846
timestamp 1682952543
transform 1 0 804 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9885
timestamp 1682952543
transform 1 0 772 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_9886
timestamp 1682952543
transform 1 0 836 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9747
timestamp 1682952543
transform 1 0 772 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9899
timestamp 1682952543
transform 1 0 804 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9797
timestamp 1682952543
transform 1 0 796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9798
timestamp 1682952543
transform 1 0 852 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_614
timestamp 1682952543
transform 1 0 760 0 -1 170
box -8 -3 104 105
use FILL  FILL_3978
timestamp 1682952543
transform 1 0 856 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9887
timestamp 1682952543
transform 1 0 876 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9748
timestamp 1682952543
transform 1 0 876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9799
timestamp 1682952543
transform 1 0 908 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9800
timestamp 1682952543
transform 1 0 956 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_615
timestamp 1682952543
transform 1 0 864 0 -1 170
box -8 -3 104 105
use FILL  FILL_3979
timestamp 1682952543
transform 1 0 960 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9888
timestamp 1682952543
transform 1 0 980 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9749
timestamp 1682952543
transform 1 0 980 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9801
timestamp 1682952543
transform 1 0 1004 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9802
timestamp 1682952543
transform 1 0 1060 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_620
timestamp 1682952543
transform 1 0 968 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9847
timestamp 1682952543
transform 1 0 1076 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9848
timestamp 1682952543
transform 1 0 1132 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9867
timestamp 1682952543
transform 1 0 1132 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_9889
timestamp 1682952543
transform 1 0 1156 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9750
timestamp 1682952543
transform 1 0 1156 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9803
timestamp 1682952543
transform 1 0 1076 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9804
timestamp 1682952543
transform 1 0 1132 0 1 125
box -2 -2 2 2
use FILL  FILL_4019
timestamp 1682952543
transform 1 0 1064 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9868
timestamp 1682952543
transform 1 0 1180 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_9900
timestamp 1682952543
transform 1 0 1172 0 1 135
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_621
timestamp 1682952543
transform -1 0 1168 0 -1 170
box -8 -3 104 105
use FILL  FILL_4020
timestamp 1682952543
transform 1 0 1168 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9869
timestamp 1682952543
transform 1 0 1268 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_9890
timestamp 1682952543
transform 1 0 1188 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_9891
timestamp 1682952543
transform 1 0 1204 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9751
timestamp 1682952543
transform 1 0 1188 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9901
timestamp 1682952543
transform 1 0 1276 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9805
timestamp 1682952543
transform 1 0 1220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9806
timestamp 1682952543
transform 1 0 1268 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_622
timestamp 1682952543
transform 1 0 1176 0 -1 170
box -8 -3 104 105
use FILL  FILL_4021
timestamp 1682952543
transform 1 0 1272 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9752
timestamp 1682952543
transform 1 0 1292 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9902
timestamp 1682952543
transform 1 0 1316 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_9916
timestamp 1682952543
transform 1 0 1292 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9807
timestamp 1682952543
transform 1 0 1316 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_623
timestamp 1682952543
transform 1 0 1280 0 -1 170
box -8 -3 104 105
use FILL  FILL_4022
timestamp 1682952543
transform 1 0 1376 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9870
timestamp 1682952543
transform 1 0 1396 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9808
timestamp 1682952543
transform 1 0 1396 0 1 125
box -2 -2 2 2
use INVX2  INVX2_709
timestamp 1682952543
transform 1 0 1384 0 -1 170
box -9 -3 26 105
use FILL  FILL_4023
timestamp 1682952543
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9753
timestamp 1682952543
transform 1 0 1420 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9917
timestamp 1682952543
transform 1 0 1420 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9754
timestamp 1682952543
transform 1 0 1516 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9809
timestamp 1682952543
transform 1 0 1444 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9810
timestamp 1682952543
transform 1 0 1500 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9944
timestamp 1682952543
transform 1 0 1452 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_624
timestamp 1682952543
transform 1 0 1408 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9918
timestamp 1682952543
transform 1 0 1516 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9811
timestamp 1682952543
transform 1 0 1540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9812
timestamp 1682952543
transform 1 0 1596 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_625
timestamp 1682952543
transform 1 0 1504 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9849
timestamp 1682952543
transform 1 0 1612 0 1 165
box -3 -3 3 3
use FILL  FILL_4024
timestamp 1682952543
transform 1 0 1600 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9850
timestamp 1682952543
transform 1 0 1628 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9871
timestamp 1682952543
transform 1 0 1620 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_9851
timestamp 1682952543
transform 1 0 1660 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9755
timestamp 1682952543
transform 1 0 1628 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9930
timestamp 1682952543
transform 1 0 1620 0 1 115
box -3 -3 3 3
use FILL  FILL_4025
timestamp 1682952543
transform 1 0 1608 0 -1 170
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1682952543
transform 1 0 1616 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9903
timestamp 1682952543
transform 1 0 1636 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_9904
timestamp 1682952543
transform 1 0 1684 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9756
timestamp 1682952543
transform 1 0 1724 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9905
timestamp 1682952543
transform 1 0 1788 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9757
timestamp 1682952543
transform 1 0 1820 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9758
timestamp 1682952543
transform 1 0 1836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9813
timestamp 1682952543
transform 1 0 1636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9814
timestamp 1682952543
transform 1 0 1644 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9815
timestamp 1682952543
transform 1 0 1676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9816
timestamp 1682952543
transform 1 0 1740 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9817
timestamp 1682952543
transform 1 0 1796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9818
timestamp 1682952543
transform 1 0 1836 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9931
timestamp 1682952543
transform 1 0 1636 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9932
timestamp 1682952543
transform 1 0 1676 0 1 115
box -3 -3 3 3
use INVX2  INVX2_710
timestamp 1682952543
transform 1 0 1624 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_9945
timestamp 1682952543
transform 1 0 1684 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_9946
timestamp 1682952543
transform 1 0 1724 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_626
timestamp 1682952543
transform -1 0 1736 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9933
timestamp 1682952543
transform 1 0 1796 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9934
timestamp 1682952543
transform 1 0 1836 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9947
timestamp 1682952543
transform 1 0 1820 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_627
timestamp 1682952543
transform -1 0 1832 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_711
timestamp 1682952543
transform 1 0 1832 0 -1 170
box -9 -3 26 105
use FILL  FILL_4027
timestamp 1682952543
transform 1 0 1848 0 -1 170
box -8 -3 16 105
use FILL  FILL_4028
timestamp 1682952543
transform 1 0 1856 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9906
timestamp 1682952543
transform 1 0 1876 0 1 135
box -3 -3 3 3
use FILL  FILL_4029
timestamp 1682952543
transform 1 0 1864 0 -1 170
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1682952543
transform 1 0 1872 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9759
timestamp 1682952543
transform 1 0 1892 0 1 135
box -2 -2 2 2
use FILL  FILL_4031
timestamp 1682952543
transform 1 0 1880 0 -1 170
box -8 -3 16 105
use FILL  FILL_4032
timestamp 1682952543
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1682952543
transform 1 0 1896 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9852
timestamp 1682952543
transform 1 0 1988 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9853
timestamp 1682952543
transform 1 0 2004 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9760
timestamp 1682952543
transform 1 0 2004 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9819
timestamp 1682952543
transform 1 0 1916 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9820
timestamp 1682952543
transform 1 0 1924 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9821
timestamp 1682952543
transform 1 0 1956 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9935
timestamp 1682952543
transform 1 0 1916 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9936
timestamp 1682952543
transform 1 0 1956 0 1 115
box -3 -3 3 3
use INVX2  INVX2_712
timestamp 1682952543
transform 1 0 1904 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_9761
timestamp 1682952543
transform 1 0 2020 0 1 135
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_628
timestamp 1682952543
transform -1 0 2016 0 -1 170
box -8 -3 104 105
use FILL  FILL_4034
timestamp 1682952543
transform 1 0 2016 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9854
timestamp 1682952543
transform 1 0 2116 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9855
timestamp 1682952543
transform 1 0 2132 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9856
timestamp 1682952543
transform 1 0 2172 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9857
timestamp 1682952543
transform 1 0 2204 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9907
timestamp 1682952543
transform 1 0 2100 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9762
timestamp 1682952543
transform 1 0 2124 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9822
timestamp 1682952543
transform 1 0 2036 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9823
timestamp 1682952543
transform 1 0 2044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9824
timestamp 1682952543
transform 1 0 2076 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9937
timestamp 1682952543
transform 1 0 2036 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9938
timestamp 1682952543
transform 1 0 2076 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9939
timestamp 1682952543
transform 1 0 2124 0 1 115
box -3 -3 3 3
use INVX2  INVX2_713
timestamp 1682952543
transform 1 0 2024 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_629
timestamp 1682952543
transform -1 0 2136 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9892
timestamp 1682952543
transform 1 0 2164 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9763
timestamp 1682952543
transform 1 0 2148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9825
timestamp 1682952543
transform 1 0 2172 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_630
timestamp 1682952543
transform 1 0 2136 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9858
timestamp 1682952543
transform 1 0 2260 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9764
timestamp 1682952543
transform 1 0 2260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9765
timestamp 1682952543
transform 1 0 2356 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9859
timestamp 1682952543
transform 1 0 2524 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9766
timestamp 1682952543
transform 1 0 2524 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9826
timestamp 1682952543
transform 1 0 2244 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9827
timestamp 1682952543
transform 1 0 2308 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9828
timestamp 1682952543
transform 1 0 2340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9829
timestamp 1682952543
transform 1 0 2396 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9830
timestamp 1682952543
transform 1 0 2436 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9831
timestamp 1682952543
transform 1 0 2444 0 1 125
box -2 -2 2 2
use INVX2  INVX2_714
timestamp 1682952543
transform 1 0 2232 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_9948
timestamp 1682952543
transform 1 0 2300 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_631
timestamp 1682952543
transform 1 0 2248 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9940
timestamp 1682952543
transform 1 0 2356 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_632
timestamp 1682952543
transform 1 0 2344 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9919
timestamp 1682952543
transform 1 0 2492 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9832
timestamp 1682952543
transform 1 0 2500 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9941
timestamp 1682952543
transform 1 0 2524 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_633
timestamp 1682952543
transform -1 0 2536 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_9767
timestamp 1682952543
transform 1 0 2548 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9920
timestamp 1682952543
transform 1 0 2548 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_9872
timestamp 1682952543
transform 1 0 2676 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9768
timestamp 1682952543
transform 1 0 2716 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9833
timestamp 1682952543
transform 1 0 2572 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9834
timestamp 1682952543
transform 1 0 2628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9835
timestamp 1682952543
transform 1 0 2636 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9836
timestamp 1682952543
transform 1 0 2684 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9950
timestamp 1682952543
transform 1 0 2548 0 1 95
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_634
timestamp 1682952543
transform 1 0 2536 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9921
timestamp 1682952543
transform 1 0 2716 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9769
timestamp 1682952543
transform 1 0 2732 0 1 135
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_635
timestamp 1682952543
transform -1 0 2728 0 -1 170
box -8 -3 104 105
use FILL  FILL_4035
timestamp 1682952543
transform 1 0 2728 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9770
timestamp 1682952543
transform 1 0 2836 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9837
timestamp 1682952543
transform 1 0 2748 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9838
timestamp 1682952543
transform 1 0 2756 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9839
timestamp 1682952543
transform 1 0 2788 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9942
timestamp 1682952543
transform 1 0 2748 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_9943
timestamp 1682952543
transform 1 0 2788 0 1 115
box -3 -3 3 3
use INVX2  INVX2_715
timestamp 1682952543
transform 1 0 2736 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_636
timestamp 1682952543
transform -1 0 2848 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9860
timestamp 1682952543
transform 1 0 2860 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9861
timestamp 1682952543
transform 1 0 2916 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9862
timestamp 1682952543
transform 1 0 2940 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9771
timestamp 1682952543
transform 1 0 2860 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9922
timestamp 1682952543
transform 1 0 2860 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9840
timestamp 1682952543
transform 1 0 2884 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9841
timestamp 1682952543
transform 1 0 2940 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_637
timestamp 1682952543
transform 1 0 2848 0 -1 170
box -8 -3 104 105
use FILL  FILL_4036
timestamp 1682952543
transform 1 0 2944 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9863
timestamp 1682952543
transform 1 0 3004 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9864
timestamp 1682952543
transform 1 0 3044 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9772
timestamp 1682952543
transform 1 0 2964 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9923
timestamp 1682952543
transform 1 0 2964 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9842
timestamp 1682952543
transform 1 0 2996 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_638
timestamp 1682952543
transform 1 0 2952 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9865
timestamp 1682952543
transform 1 0 3060 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_9843
timestamp 1682952543
transform 1 0 3060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9844
timestamp 1682952543
transform 1 0 3068 0 1 125
box -2 -2 2 2
use INVX2  INVX2_716
timestamp 1682952543
transform 1 0 3048 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_9773
timestamp 1682952543
transform 1 0 3076 0 1 135
box -2 -2 2 2
use INVX2  INVX2_717
timestamp 1682952543
transform -1 0 3080 0 -1 170
box -9 -3 26 105
use FILL  FILL_4037
timestamp 1682952543
transform 1 0 3080 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9774
timestamp 1682952543
transform 1 0 3100 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9924
timestamp 1682952543
transform 1 0 3100 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9845
timestamp 1682952543
transform 1 0 3148 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_639
timestamp 1682952543
transform 1 0 3088 0 -1 170
box -8 -3 104 105
use FILL  FILL_4038
timestamp 1682952543
transform 1 0 3184 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9775
timestamp 1682952543
transform 1 0 3220 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9908
timestamp 1682952543
transform 1 0 3268 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_9909
timestamp 1682952543
transform 1 0 3292 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9846
timestamp 1682952543
transform 1 0 3204 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9847
timestamp 1682952543
transform 1 0 3268 0 1 125
box -2 -2 2 2
use INVX2  INVX2_718
timestamp 1682952543
transform 1 0 3192 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_640
timestamp 1682952543
transform 1 0 3208 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_9866
timestamp 1682952543
transform 1 0 3340 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_9873
timestamp 1682952543
transform 1 0 3332 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9776
timestamp 1682952543
transform 1 0 3332 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9848
timestamp 1682952543
transform 1 0 3316 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9849
timestamp 1682952543
transform 1 0 3356 0 1 125
box -2 -2 2 2
use INVX2  INVX2_719
timestamp 1682952543
transform 1 0 3304 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_641
timestamp 1682952543
transform 1 0 3320 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_9850
timestamp 1682952543
transform 1 0 3428 0 1 125
box -2 -2 2 2
use INVX2  INVX2_720
timestamp 1682952543
transform 1 0 3416 0 -1 170
box -9 -3 26 105
use FILL  FILL_4039
timestamp 1682952543
transform 1 0 3432 0 -1 170
box -8 -3 16 105
use FILL  FILL_4040
timestamp 1682952543
transform 1 0 3440 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9874
timestamp 1682952543
transform 1 0 3460 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_9893
timestamp 1682952543
transform 1 0 3500 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9777
timestamp 1682952543
transform 1 0 3460 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9910
timestamp 1682952543
transform 1 0 3508 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_9911
timestamp 1682952543
transform 1 0 3540 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9851
timestamp 1682952543
transform 1 0 3508 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_642
timestamp 1682952543
transform 1 0 3448 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_9852
timestamp 1682952543
transform 1 0 3556 0 1 125
box -2 -2 2 2
use INVX2  INVX2_727
timestamp 1682952543
transform 1 0 3544 0 -1 170
box -9 -3 26 105
use FILL  FILL_4054
timestamp 1682952543
transform 1 0 3560 0 -1 170
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1682952543
transform 1 0 3568 0 -1 170
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1682952543
transform 1 0 3576 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9875
timestamp 1682952543
transform 1 0 3596 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9778
timestamp 1682952543
transform 1 0 3596 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9853
timestamp 1682952543
transform 1 0 3628 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9854
timestamp 1682952543
transform 1 0 3676 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_9949
timestamp 1682952543
transform 1 0 3620 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_643
timestamp 1682952543
transform 1 0 3584 0 -1 170
box -8 -3 104 105
use FILL  FILL_4057
timestamp 1682952543
transform 1 0 3680 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9894
timestamp 1682952543
transform 1 0 3700 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9779
timestamp 1682952543
transform 1 0 3700 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9855
timestamp 1682952543
transform 1 0 3724 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9856
timestamp 1682952543
transform 1 0 3780 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_644
timestamp 1682952543
transform 1 0 3688 0 -1 170
box -8 -3 104 105
use FILL  FILL_4058
timestamp 1682952543
transform 1 0 3784 0 -1 170
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1682952543
transform 1 0 3792 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9895
timestamp 1682952543
transform 1 0 3812 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9780
timestamp 1682952543
transform 1 0 3812 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9857
timestamp 1682952543
transform 1 0 3860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9858
timestamp 1682952543
transform 1 0 3892 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_645
timestamp 1682952543
transform 1 0 3800 0 -1 170
box -8 -3 104 105
use FILL  FILL_4060
timestamp 1682952543
transform 1 0 3896 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9876
timestamp 1682952543
transform 1 0 3916 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_9877
timestamp 1682952543
transform 1 0 3948 0 1 155
box -3 -3 3 3
use FILL  FILL_4061
timestamp 1682952543
transform 1 0 3904 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9896
timestamp 1682952543
transform 1 0 3924 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_9897
timestamp 1682952543
transform 1 0 3988 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9781
timestamp 1682952543
transform 1 0 3924 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9912
timestamp 1682952543
transform 1 0 3956 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9859
timestamp 1682952543
transform 1 0 3948 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9860
timestamp 1682952543
transform 1 0 4004 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_646
timestamp 1682952543
transform 1 0 3912 0 -1 170
box -8 -3 104 105
use FILL  FILL_4062
timestamp 1682952543
transform 1 0 4008 0 -1 170
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1682952543
transform 1 0 4016 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_9898
timestamp 1682952543
transform 1 0 4036 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9782
timestamp 1682952543
transform 1 0 4036 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_9913
timestamp 1682952543
transform 1 0 4060 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_9914
timestamp 1682952543
transform 1 0 4084 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_9915
timestamp 1682952543
transform 1 0 4116 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9861
timestamp 1682952543
transform 1 0 4060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9862
timestamp 1682952543
transform 1 0 4116 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_647
timestamp 1682952543
transform 1 0 4024 0 -1 170
box -8 -3 104 105
use FILL  FILL_4064
timestamp 1682952543
transform 1 0 4120 0 -1 170
box -8 -3 16 105
use FILL  FILL_4066
timestamp 1682952543
transform 1 0 4128 0 -1 170
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1682952543
transform 1 0 4136 0 -1 170
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1682952543
transform 1 0 4144 0 -1 170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_81
timestamp 1682952543
transform 1 0 4201 0 1 70
box -10 -3 10 3
use M3_M2  M3_M2_9951
timestamp 1682952543
transform 1 0 2404 0 1 65
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_4
timestamp 1682952543
transform 1 0 48 0 1 47
box -10 -10 10 10
use M3_M2  M3_M2_9952
timestamp 1682952543
transform 1 0 292 0 1 55
box -3 -3 3 3
use M3_M2  M3_M2_9953
timestamp 1682952543
transform 1 0 1604 0 1 45
box -3 -3 3 3
use M3_M2  M3_M2_9954
timestamp 1682952543
transform 1 0 2692 0 1 45
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_5
timestamp 1682952543
transform 1 0 4177 0 1 47
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_6
timestamp 1682952543
transform 1 0 24 0 1 23
box -10 -10 10 10
use M3_M2  M3_M2_9955
timestamp 1682952543
transform 1 0 1748 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_9956
timestamp 1682952543
transform 1 0 2740 0 1 25
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_7
timestamp 1682952543
transform 1 0 4201 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal2 2740 4138 2740 4138 6 clka
rlabel metal3 2 2325 2 2325 6 clkb
rlabel metal2 2756 4138 2756 4138 6 reset
rlabel metal2 2100 4138 2100 4138 6 we_ins
rlabel metal2 2052 4138 2052 4138 6 load[15]
rlabel metal2 1876 4138 1876 4138 6 load[14]
rlabel metal2 1916 4138 1916 4138 6 load[13]
rlabel metal2 1900 4138 1900 4138 6 load[12]
rlabel metal2 2020 4138 2020 4138 6 load[11]
rlabel metal2 1988 4138 1988 4138 6 load[10]
rlabel metal2 1932 4138 1932 4138 6 load[9]
rlabel metal2 1844 4138 1844 4138 6 load[8]
rlabel metal2 1948 4138 1948 4138 6 load[7]
rlabel metal2 2036 4138 2036 4138 6 load[6]
rlabel metal2 2004 4138 2004 4138 6 load[5]
rlabel metal2 2116 4138 2116 4138 6 load[4]
rlabel metal2 1972 4138 1972 4138 6 load[3]
rlabel metal2 2068 4138 2068 4138 6 load[2]
rlabel metal2 2084 4138 2084 4138 6 load[1]
rlabel metal2 1860 4138 1860 4138 6 load[0]
rlabel metal2 2684 4138 2684 4138 6 reg_0_out[7]
rlabel metal2 3116 4138 3116 4138 6 reg_0_out[6]
rlabel metal3 4224 3335 4224 3335 6 reg_0_out[5]
rlabel metal3 4224 3315 4224 3315 6 reg_0_out[4]
rlabel metal3 4224 3365 4224 3365 6 reg_0_out[3]
rlabel metal2 3308 4138 3308 4138 6 reg_0_out[2]
rlabel metal2 2820 4138 2820 4138 6 reg_0_out[1]
rlabel metal2 2948 4138 2948 4138 6 reg_0_out[0]
rlabel metal1 38 167 38 167 6 gnd
rlabel metal1 14 67 14 67 6 vdd
<< end >>

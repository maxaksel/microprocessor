magic
tech scmos
timestamp 1682952861
use with_frame_and_fill  with_frame_and_fill_0
timestamp 1682952543
transform 1 0 0 0 1 0
box -2500 -2400 4300 4400
<< end >>

magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -5 48 126 105
rect 23 46 100 48
rect 65 39 100 46
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
rect 23 6 25 26
rect 31 6 33 26
rect 36 6 38 26
rect 44 6 46 26
rect 52 6 54 26
rect 60 6 62 26
rect 68 6 70 26
rect 77 6 79 26
rect 82 6 84 26
rect 87 6 89 26
rect 95 6 97 16
rect 111 6 113 16
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
rect 31 54 33 94
rect 36 54 38 94
rect 44 54 46 94
rect 52 58 54 94
rect 60 58 62 94
rect 68 58 70 94
rect 77 46 79 94
rect 82 46 84 94
rect 87 46 89 94
rect 95 74 97 94
rect 111 74 113 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 6 15 26
rect 17 6 23 26
rect 25 6 31 26
rect 33 6 36 26
rect 38 6 44 26
rect 46 6 52 26
rect 54 6 60 26
rect 62 6 68 26
rect 70 6 77 26
rect 79 6 82 26
rect 84 6 87 26
rect 89 16 94 26
rect 89 6 95 16
rect 97 6 102 16
rect 106 6 111 16
rect 113 6 118 16
<< pdiffusion >>
rect 2 54 7 94
rect 9 54 15 94
rect 17 54 23 94
rect 25 54 31 94
rect 33 54 36 94
rect 38 54 44 94
rect 46 58 52 94
rect 54 58 60 94
rect 62 58 68 94
rect 70 58 77 94
rect 46 54 51 58
rect 71 51 77 58
rect 72 47 77 51
rect 74 46 77 47
rect 79 46 82 94
rect 84 46 87 94
rect 89 74 95 94
rect 97 74 102 94
rect 106 74 111 94
rect 113 74 118 94
rect 89 46 94 74
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
rect 46 -2 50 2
rect 62 -2 66 2
rect 78 -2 82 2
rect 94 -2 98 2
rect 110 -2 114 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
rect 46 98 50 102
rect 62 98 66 102
rect 78 98 82 102
rect 94 98 98 102
rect 110 98 114 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 36 94 38 96
rect 44 94 46 96
rect 52 94 54 96
rect 60 94 62 96
rect 68 94 70 96
rect 77 94 79 96
rect 82 94 84 96
rect 87 94 89 96
rect 95 94 97 96
rect 111 94 113 96
rect 7 33 9 54
rect 15 39 17 54
rect 23 47 25 54
rect 22 43 26 47
rect 14 35 18 39
rect 6 29 10 33
rect 7 26 9 29
rect 15 26 17 35
rect 23 26 25 43
rect 31 39 33 54
rect 36 53 38 54
rect 44 53 46 54
rect 52 53 54 58
rect 60 57 62 58
rect 68 57 70 58
rect 36 51 46 53
rect 49 51 54 53
rect 57 55 62 57
rect 66 55 70 57
rect 29 35 33 39
rect 31 26 33 35
rect 37 32 39 51
rect 49 38 51 51
rect 57 45 59 55
rect 66 51 68 55
rect 64 47 68 51
rect 55 41 59 45
rect 47 36 51 38
rect 47 34 54 36
rect 37 29 41 32
rect 36 27 46 29
rect 36 26 38 27
rect 44 26 46 27
rect 52 26 54 34
rect 57 29 59 41
rect 66 29 68 47
rect 95 73 97 74
rect 95 71 99 73
rect 77 44 79 46
rect 72 42 79 44
rect 72 40 76 42
rect 74 29 76 40
rect 82 38 84 46
rect 87 44 89 46
rect 87 42 91 44
rect 80 34 84 38
rect 57 27 62 29
rect 66 27 70 29
rect 74 27 79 29
rect 60 26 62 27
rect 68 26 70 27
rect 77 26 79 27
rect 82 26 84 34
rect 89 38 91 42
rect 97 39 99 71
rect 111 57 113 74
rect 108 53 113 57
rect 89 34 93 38
rect 97 35 101 39
rect 89 30 91 34
rect 87 28 91 30
rect 87 26 89 28
rect 97 25 99 35
rect 95 23 99 25
rect 95 16 97 23
rect 111 16 113 53
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
rect 31 4 33 6
rect 36 4 38 6
rect 44 4 46 6
rect 52 4 54 6
rect 60 4 62 6
rect 68 4 70 6
rect 77 4 79 6
rect 82 4 84 6
rect 87 4 89 6
rect 95 4 97 6
rect 111 4 113 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 31 99 33 101
rect 47 99 49 101
rect 63 99 65 101
rect 79 99 81 101
rect 95 99 97 101
rect 111 99 113 101
rect 3 90 5 92
rect 11 91 13 93
rect 19 90 21 92
rect 27 90 29 92
rect 40 90 42 92
rect 48 90 50 92
rect 56 90 58 92
rect 64 90 66 92
rect 72 89 74 91
rect 91 89 93 91
rect 99 90 101 92
rect 107 90 109 92
rect 115 90 117 92
rect 3 85 5 87
rect 11 86 13 88
rect 19 85 21 87
rect 27 85 29 87
rect 40 85 42 87
rect 48 85 50 87
rect 56 85 58 87
rect 64 85 66 87
rect 72 84 74 86
rect 91 84 93 86
rect 99 85 101 87
rect 107 85 109 87
rect 115 85 117 87
rect 3 80 5 82
rect 11 81 13 83
rect 19 80 21 82
rect 27 80 29 82
rect 40 80 42 82
rect 48 80 50 82
rect 56 80 58 82
rect 64 80 66 82
rect 72 79 74 81
rect 91 79 93 81
rect 99 80 101 82
rect 107 80 109 82
rect 115 80 117 82
rect 3 75 5 77
rect 11 76 13 78
rect 19 75 21 77
rect 27 75 29 77
rect 40 75 42 77
rect 48 75 50 77
rect 56 75 58 77
rect 64 75 66 77
rect 72 74 74 76
rect 91 74 93 76
rect 99 75 101 77
rect 107 75 109 77
rect 115 75 117 77
rect 3 70 5 72
rect 11 71 13 73
rect 19 70 21 72
rect 27 70 29 72
rect 40 70 42 72
rect 48 70 50 72
rect 56 70 58 72
rect 64 70 66 72
rect 72 69 74 71
rect 91 69 93 71
rect 3 65 5 67
rect 11 66 13 68
rect 19 65 21 67
rect 27 65 29 67
rect 40 65 42 67
rect 48 65 50 67
rect 56 65 58 67
rect 64 65 66 67
rect 72 64 74 66
rect 91 64 93 66
rect 3 60 5 62
rect 11 61 13 63
rect 19 60 21 62
rect 27 60 29 62
rect 40 60 42 62
rect 48 60 50 62
rect 64 60 66 62
rect 72 59 74 61
rect 91 59 93 61
rect 3 55 5 57
rect 19 55 21 57
rect 40 55 42 57
rect 48 55 50 57
rect 72 54 74 56
rect 91 54 93 56
rect 109 54 111 56
rect 65 48 67 50
rect 91 49 93 51
rect 23 44 25 46
rect 56 42 58 44
rect 73 41 75 43
rect 15 36 17 38
rect 30 36 32 38
rect 48 35 50 37
rect 81 35 83 37
rect 90 35 92 37
rect 98 36 100 38
rect 7 30 9 32
rect 38 29 40 31
rect 3 22 5 24
rect 19 22 21 24
rect 48 22 50 24
rect 64 22 66 24
rect 91 22 93 24
rect 3 17 5 19
rect 11 17 13 19
rect 19 17 21 19
rect 27 18 29 20
rect 40 19 42 21
rect 48 17 50 19
rect 64 17 66 19
rect 72 17 74 19
rect 91 17 93 19
rect 3 12 5 14
rect 11 12 13 14
rect 19 12 21 14
rect 27 13 29 15
rect 40 14 42 16
rect 56 14 58 16
rect 48 12 50 14
rect 64 12 66 14
rect 72 12 74 14
rect 91 12 93 14
rect 99 12 101 14
rect 107 12 109 14
rect 115 12 117 14
rect 3 7 5 9
rect 11 7 13 9
rect 19 7 21 9
rect 27 8 29 10
rect 40 9 42 11
rect 56 9 58 11
rect 48 7 50 9
rect 64 7 66 9
rect 72 7 74 9
rect 91 7 93 9
rect 99 7 101 9
rect 107 7 109 9
rect 115 7 117 9
rect -1 -1 1 1
rect 15 -1 17 1
rect 31 -1 33 1
rect 47 -1 49 1
rect 63 -1 65 1
rect 79 -1 81 1
rect 95 -1 97 1
rect 111 -1 113 1
<< metal1 >>
rect -2 97 122 103
rect 2 57 6 94
rect 10 60 14 97
rect 18 57 22 94
rect 2 54 22 57
rect 26 54 30 94
rect 39 54 43 97
rect 47 61 51 94
rect 55 64 59 97
rect 63 61 67 94
rect 47 58 67 61
rect 47 54 51 58
rect 60 51 64 52
rect 71 51 76 94
rect 60 48 68 51
rect 64 47 68 48
rect 72 47 76 51
rect 10 43 14 47
rect 18 46 26 47
rect 90 46 94 97
rect 98 77 102 94
rect 97 74 102 77
rect 106 74 110 97
rect 114 74 118 94
rect 97 49 100 74
rect 104 53 112 57
rect 97 46 107 49
rect 18 45 55 46
rect 18 44 59 45
rect 18 43 76 44
rect 11 39 14 43
rect 52 41 76 43
rect 72 40 76 41
rect 11 38 18 39
rect 29 38 33 39
rect 11 37 51 38
rect 80 37 84 38
rect 2 33 6 37
rect 11 36 84 37
rect 14 35 84 36
rect 47 34 84 35
rect 89 34 93 38
rect 97 35 101 43
rect 3 32 10 33
rect 3 31 41 32
rect 89 31 92 34
rect 3 30 92 31
rect 6 29 92 30
rect 37 28 92 29
rect 104 27 107 46
rect 115 37 118 74
rect 114 33 118 37
rect 2 23 22 26
rect 2 6 6 23
rect 10 3 14 20
rect 18 6 22 23
rect 26 6 30 26
rect 39 3 43 24
rect 47 22 67 25
rect 47 6 51 22
rect 55 3 59 19
rect 63 6 67 22
rect 72 21 76 25
rect 71 6 76 21
rect 90 3 94 25
rect 104 23 110 27
rect 104 22 107 23
rect 99 19 107 22
rect 99 16 102 19
rect 115 16 118 33
rect 98 6 102 16
rect 106 3 110 16
rect 114 6 118 16
rect -2 -3 122 3
<< metal2 >>
rect 26 57 30 58
rect 26 54 108 57
rect 27 26 30 54
rect 60 48 64 54
rect 104 53 108 54
rect 72 47 76 51
rect 26 22 30 26
rect 73 42 76 47
rect 97 42 101 43
rect 73 39 101 42
rect 73 25 76 39
rect 72 21 76 25
<< gv1 >>
rect 27 55 29 57
rect 105 54 107 56
rect 61 49 63 51
rect 73 48 75 50
rect 98 40 100 42
rect 27 23 29 25
rect 73 22 75 24
<< m1p >>
rect 10 43 14 47
rect 18 43 22 47
rect 2 33 6 37
rect 114 33 118 37
rect 106 23 110 27
<< labels >>
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 35 4 35 6 A
rlabel metal1 12 45 12 45 6 B
rlabel metal1 20 45 20 45 6 C
rlabel metal1 116 35 116 35 6 YC
rlabel metal1 108 25 108 25 6 YS
<< end >>

magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 40 105
<< ntransistor >>
rect 7 6 9 26
rect 12 6 14 26
rect 20 6 22 16
<< ptransistor >>
rect 7 74 9 94
rect 15 74 17 94
rect 23 74 25 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 6 12 26
rect 14 16 19 26
rect 14 6 20 16
rect 22 6 27 16
<< pdiffusion >>
rect 2 74 7 94
rect 9 74 15 94
rect 17 74 23 94
rect 25 74 30 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 7 41 9 74
rect 15 53 17 74
rect 13 49 17 53
rect 2 37 9 41
rect 15 39 17 49
rect 7 26 9 37
rect 12 37 17 39
rect 12 26 14 37
rect 23 33 25 74
rect 20 30 25 33
rect 20 29 24 30
rect 20 16 22 29
rect 7 4 9 6
rect 12 4 14 6
rect 20 4 22 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 3 90 5 92
rect 11 90 13 92
rect 19 90 21 92
rect 27 90 29 92
rect 3 85 5 87
rect 11 85 13 87
rect 19 85 21 87
rect 27 85 29 87
rect 3 80 5 82
rect 11 80 13 82
rect 19 80 21 82
rect 27 80 29 82
rect 3 75 5 77
rect 11 75 13 77
rect 19 75 21 77
rect 27 75 29 77
rect 14 50 16 52
rect 3 38 5 40
rect 21 30 23 32
rect 3 22 5 24
rect 16 22 18 24
rect 3 17 5 19
rect 16 17 18 19
rect 3 12 5 14
rect 16 12 18 14
rect 24 12 26 14
rect 3 7 5 9
rect 16 7 18 9
rect 24 7 26 9
rect -1 -1 1 1
rect 15 -1 17 1
<< metal1 >>
rect -2 97 34 103
rect 2 74 6 97
rect 10 74 14 94
rect 18 74 22 97
rect 26 74 30 94
rect 11 71 14 74
rect 11 68 23 71
rect 10 53 17 57
rect 13 49 17 53
rect 2 33 6 41
rect 20 33 23 68
rect 27 67 30 74
rect 26 63 30 67
rect 9 30 24 33
rect 9 29 12 30
rect 20 29 24 30
rect 3 26 12 29
rect 2 6 6 26
rect 15 3 19 26
rect 27 19 30 63
rect 23 16 30 19
rect 23 6 27 16
rect -2 -3 34 3
<< m1p >>
rect 26 63 30 67
rect 10 53 14 57
rect 2 33 6 37
<< labels >>
rlabel metal1 28 65 28 65 6 Y
rlabel metal1 12 55 12 55 6 B
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 35 4 35 6 A
<< end >>

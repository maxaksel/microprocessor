magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 46 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
rect 23 6 25 26
rect 31 6 33 26
<< ptransistor >>
rect 7 54 9 94
rect 12 54 14 94
rect 26 54 28 94
rect 31 54 33 94
<< ndiffusion >>
rect 2 6 7 26
rect 9 6 15 26
rect 17 6 23 26
rect 25 6 31 26
rect 33 6 38 26
<< pdiffusion >>
rect 2 54 7 94
rect 9 54 12 94
rect 14 54 26 94
rect 28 54 31 94
rect 33 54 38 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
<< polysilicon >>
rect 7 94 9 96
rect 12 94 14 96
rect 26 94 28 96
rect 31 94 33 96
rect 7 49 9 54
rect 12 53 14 54
rect 26 53 28 54
rect 12 51 17 53
rect 4 47 9 49
rect 4 35 6 47
rect 15 43 17 51
rect 10 39 17 43
rect 4 33 10 35
rect 6 31 10 33
rect 7 26 9 31
rect 15 26 17 39
rect 25 51 28 53
rect 31 53 33 54
rect 31 51 37 53
rect 25 43 27 51
rect 25 39 30 43
rect 35 41 37 51
rect 25 31 27 39
rect 34 37 38 41
rect 23 29 27 31
rect 35 30 37 37
rect 23 26 25 29
rect 31 28 37 30
rect 31 26 33 28
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
rect 31 4 33 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 31 99 33 101
rect 3 90 5 92
rect 16 90 18 92
rect 21 90 23 92
rect 35 90 37 92
rect 3 85 5 87
rect 16 85 18 87
rect 21 85 23 87
rect 35 85 37 87
rect 3 80 5 82
rect 16 80 18 82
rect 21 80 23 82
rect 35 80 37 82
rect 3 75 5 77
rect 16 75 18 77
rect 21 75 23 77
rect 35 75 37 77
rect 3 70 5 72
rect 16 70 18 72
rect 21 70 23 72
rect 35 70 37 72
rect 3 65 5 67
rect 16 65 18 67
rect 21 65 23 67
rect 35 65 37 67
rect 3 60 5 62
rect 16 60 18 62
rect 21 60 23 62
rect 35 60 37 62
rect 3 55 5 57
rect 16 55 18 57
rect 21 55 23 57
rect 35 55 37 57
rect 11 40 13 42
rect 27 40 29 42
rect 35 38 37 40
rect 7 32 9 34
rect 3 22 5 24
rect 19 22 21 24
rect 27 23 29 25
rect 35 22 37 24
rect 3 17 5 19
rect 11 18 13 20
rect 19 17 21 19
rect 27 18 29 20
rect 35 17 37 19
rect 3 12 5 14
rect 11 13 13 15
rect 19 12 21 14
rect 27 13 29 15
rect 35 12 37 14
rect 3 7 5 9
rect 11 8 13 10
rect 19 7 21 9
rect 35 7 37 9
rect -1 -1 1 1
rect 15 -1 17 1
rect 31 -1 33 1
<< metal1 >>
rect -2 97 42 103
rect 2 54 6 97
rect 15 54 25 94
rect 34 54 38 97
rect 10 39 14 47
rect 18 37 21 54
rect 26 39 30 47
rect 2 36 6 37
rect 18 36 22 37
rect 2 33 10 36
rect 18 33 30 36
rect 34 33 38 41
rect 6 31 10 33
rect 3 26 21 28
rect 27 26 30 33
rect 2 25 22 26
rect 2 6 6 25
rect 10 3 14 22
rect 18 9 22 25
rect 26 12 30 26
rect 34 9 38 26
rect 18 6 38 9
rect -2 -3 42 3
<< m1p >>
rect 10 43 14 47
rect 26 43 30 47
rect 2 33 6 37
rect 18 33 22 37
rect 34 33 38 37
<< labels >>
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 28 45 28 45 6 D
rlabel metal1 36 35 36 35 6 C
rlabel metal1 4 35 4 35 6 A
rlabel metal1 12 45 12 45 6 B
rlabel metal1 20 35 20 35 6 Y
<< end >>

magic
tech scmos
timestamp 1677622389
<< m2contact >>
rect -2 -2 2 2
<< end >>

magic
tech scmos
timestamp 1677677812
<< metal1 >>
rect 14 4707 4853 4727
rect 38 4683 4829 4703
rect 14 4667 4853 4673
rect 2812 4623 2829 4626
rect 116 4613 125 4616
rect 172 4613 181 4616
rect 314 4613 324 4616
rect 484 4613 493 4616
rect 586 4613 612 4616
rect 836 4613 861 4616
rect 892 4613 941 4616
rect 1066 4613 1092 4616
rect 1162 4613 1180 4616
rect 1226 4613 1236 4616
rect 1418 4613 1452 4616
rect 1612 4613 1621 4616
rect 1668 4613 1677 4616
rect 2012 4613 2037 4616
rect 2132 4613 2141 4616
rect 2338 4613 2356 4616
rect 2410 4613 2420 4616
rect 2466 4613 2476 4616
rect 2660 4613 2677 4616
rect 2772 4613 2781 4616
rect 2844 4613 2853 4616
rect 2890 4613 2916 4616
rect 3012 4613 3037 4616
rect 3068 4613 3085 4616
rect 3164 4613 3173 4616
rect 3220 4613 3237 4616
rect 3370 4613 3380 4616
rect 3508 4613 3533 4616
rect 3564 4613 3573 4616
rect 3580 4613 3621 4616
rect 3708 4613 3733 4616
rect 3764 4613 3773 4616
rect 3930 4613 3940 4616
rect 3946 4613 3972 4616
rect 4002 4613 4028 4616
rect 4476 4613 4501 4616
rect 4532 4613 4541 4616
rect 4764 4613 4773 4616
rect 178 4603 181 4613
rect 2778 4606 2781 4613
rect 650 4603 684 4606
rect 2778 4603 2788 4606
rect 2818 4603 2836 4606
rect 3082 4605 3085 4613
rect 3234 4605 3237 4613
rect 3570 4605 3573 4613
rect 3586 4603 3620 4606
rect 3770 4605 3773 4613
rect 3946 4605 3949 4613
rect 4538 4605 4541 4613
rect 4770 4605 4773 4613
rect 38 4567 4829 4573
rect 946 4543 972 4546
rect 2754 4543 2772 4546
rect 3362 4536 3365 4546
rect 148 4533 173 4536
rect 196 4533 276 4536
rect 298 4533 308 4536
rect 556 4533 628 4536
rect 644 4533 685 4536
rect 892 4533 909 4536
rect 932 4533 941 4536
rect 962 4533 980 4536
rect 986 4533 1020 4536
rect 1036 4533 1053 4536
rect 1090 4533 1132 4536
rect 1148 4533 1164 4536
rect 1210 4533 1244 4536
rect 1274 4533 1284 4536
rect 1314 4533 1348 4536
rect 1396 4533 1421 4536
rect 1460 4533 1493 4536
rect 1050 4526 1053 4533
rect 1530 4526 1533 4535
rect 1538 4533 1588 4536
rect 1636 4533 1653 4536
rect 1796 4533 1821 4536
rect 1852 4533 1885 4536
rect 1906 4533 1924 4536
rect 1962 4533 2020 4536
rect 2066 4533 2124 4536
rect 2180 4533 2229 4536
rect 2234 4533 2244 4536
rect 2276 4533 2300 4536
rect 2322 4533 2332 4536
rect 2354 4533 2364 4536
rect 2396 4533 2412 4536
rect 2434 4533 2444 4536
rect 2540 4533 2573 4536
rect 2602 4533 2644 4536
rect 2660 4533 2677 4536
rect 2714 4533 2724 4536
rect 2740 4533 2765 4536
rect 2786 4533 2812 4536
rect 2836 4533 2845 4536
rect 2858 4533 2892 4536
rect 2922 4533 2940 4536
rect 2964 4533 2973 4536
rect 3010 4533 3044 4536
rect 3068 4533 3077 4536
rect 3116 4533 3133 4536
rect 3188 4533 3252 4536
rect 3300 4533 3365 4536
rect 3442 4533 3500 4536
rect 3538 4533 3580 4536
rect 3596 4533 3605 4536
rect 3642 4533 3660 4536
rect 3676 4533 3733 4536
rect 3828 4533 3853 4536
rect 3884 4533 3901 4536
rect 3962 4533 4004 4536
rect 4036 4533 4068 4536
rect 4148 4533 4181 4536
rect 4194 4533 4220 4536
rect 4252 4533 4269 4536
rect 4292 4533 4301 4536
rect 4306 4533 4316 4536
rect 4362 4533 4388 4536
rect 4418 4533 4428 4536
rect 4458 4533 4516 4536
rect 4580 4533 4605 4536
rect 4610 4533 4668 4536
rect 4740 4533 4773 4536
rect 122 4523 140 4526
rect 204 4523 221 4526
rect 234 4523 268 4526
rect 420 4523 453 4526
rect 484 4523 493 4526
rect 506 4523 532 4526
rect 564 4523 589 4526
rect 610 4523 620 4526
rect 764 4523 781 4526
rect 890 4523 908 4526
rect 988 4523 1005 4526
rect 1050 4523 1061 4526
rect 1082 4523 1124 4526
rect 1162 4523 1172 4526
rect 1204 4523 1229 4526
rect 1260 4523 1285 4526
rect 1306 4523 1356 4526
rect 1362 4523 1388 4526
rect 1452 4523 1485 4526
rect 1530 4523 1596 4526
rect 1658 4523 1668 4526
rect 1716 4523 1741 4526
rect 1778 4523 1788 4526
rect 1794 4523 1828 4526
rect 1866 4523 1900 4526
rect 1906 4523 1932 4526
rect 1948 4523 1957 4526
rect 1970 4523 2012 4526
rect 2060 4523 2077 4526
rect 2082 4523 2116 4526
rect 2188 4523 2213 4526
rect 2242 4523 2252 4526
rect 2282 4523 2292 4526
rect 2346 4523 2372 4526
rect 2452 4523 2469 4526
rect 2474 4523 2516 4526
rect 2548 4523 2588 4526
rect 2594 4523 2636 4526
rect 2788 4523 2805 4526
rect 2810 4523 2820 4526
rect 2866 4523 2900 4526
rect 2922 4516 2925 4533
rect 2956 4523 2981 4526
rect 2996 4523 3045 4526
rect 3108 4523 3164 4526
rect 3282 4523 3292 4526
rect 3380 4523 3405 4526
rect 3604 4523 3645 4526
rect 3722 4523 3748 4526
rect 3786 4523 3804 4526
rect 3834 4523 3876 4526
rect 3948 4523 4012 4526
rect 4106 4523 4140 4526
rect 4186 4523 4228 4526
rect 4258 4523 4284 4526
rect 4290 4523 4324 4526
rect 4370 4523 4380 4526
rect 4426 4523 4436 4526
rect 4442 4523 4524 4526
rect 4594 4523 4676 4526
rect 4722 4523 4732 4526
rect 1084 4513 1117 4516
rect 1234 4513 1244 4516
rect 2916 4513 2925 4516
rect 3018 4513 3044 4516
rect 3386 4513 3412 4516
rect 3436 4513 3493 4516
rect 14 4467 4853 4473
rect 972 4423 1005 4426
rect 1084 4423 1093 4426
rect 2852 4423 2877 4426
rect 2932 4423 2965 4426
rect 3402 4423 3420 4426
rect 3444 4423 3477 4426
rect 3906 4423 3932 4426
rect 3946 4423 3956 4426
rect 108 4413 133 4416
rect 178 4413 188 4416
rect 386 4413 404 4416
rect 498 4413 540 4416
rect 594 4413 612 4416
rect 666 4413 700 4416
rect 820 4413 861 4416
rect 900 4413 940 4416
rect 1028 4413 1037 4416
rect 180 4403 189 4406
rect 212 4403 221 4406
rect 226 4403 236 4406
rect 412 4403 453 4406
rect 522 4403 525 4413
rect 666 4406 669 4413
rect 1186 4406 1189 4416
rect 1252 4413 1269 4416
rect 1364 4413 1389 4416
rect 1420 4413 1429 4416
rect 1500 4413 1517 4416
rect 1572 4413 1597 4416
rect 1628 4413 1637 4416
rect 570 4403 620 4406
rect 636 4403 669 4406
rect 812 4403 869 4406
rect 898 4403 932 4406
rect 1010 4403 1020 4406
rect 1090 4403 1100 4406
rect 1124 4403 1133 4406
rect 1146 4403 1172 4406
rect 1186 4403 1236 4406
rect 1426 4405 1429 4413
rect 1466 4403 1476 4406
rect 1508 4403 1533 4406
rect 1634 4405 1637 4413
rect 1714 4413 1748 4416
rect 1754 4413 1804 4416
rect 1836 4413 1861 4416
rect 1650 4403 1684 4406
rect 1714 4405 1717 4413
rect 1722 4403 1740 4406
rect 1828 4403 1884 4406
rect 1916 4403 1996 4406
rect 2018 4403 2021 4414
rect 2026 4413 2036 4416
rect 2066 4413 2092 4416
rect 2284 4413 2293 4416
rect 2404 4413 2421 4416
rect 2458 4413 2484 4416
rect 2548 4413 2565 4416
rect 2692 4413 2701 4416
rect 2826 4413 2836 4416
rect 2900 4413 2909 4416
rect 2930 4413 2973 4416
rect 3220 4413 3253 4416
rect 3364 4413 3389 4416
rect 3396 4413 3405 4416
rect 3682 4413 3724 4416
rect 3786 4413 3812 4416
rect 3834 4413 3852 4416
rect 3962 4413 4004 4416
rect 4010 4413 4044 4416
rect 4050 4413 4060 4416
rect 4090 4413 4116 4416
rect 4170 4413 4180 4416
rect 4212 4413 4221 4416
rect 4300 4413 4341 4416
rect 4378 4413 4404 4416
rect 4442 4413 4468 4416
rect 4498 4413 4508 4416
rect 4522 4413 4565 4416
rect 4748 4413 4773 4416
rect 2260 4403 2269 4406
rect 2802 4403 2828 4406
rect 2892 4403 2901 4406
rect 2932 4403 2965 4406
rect 2970 4405 2973 4413
rect 3002 4403 3012 4406
rect 3036 4403 3061 4406
rect 3100 4403 3117 4406
rect 3250 4405 3253 4413
rect 3386 4405 3389 4413
rect 3748 4403 3765 4406
rect 3820 4403 3853 4406
rect 3876 4403 3925 4406
rect 4012 4403 4029 4406
rect 4050 4405 4053 4413
rect 4162 4403 4188 4406
rect 4204 4403 4237 4406
rect 4260 4403 4285 4406
rect 4306 4403 4340 4406
rect 4428 4403 4453 4406
rect 4516 4403 4533 4406
rect 4538 4403 4548 4406
rect 4570 4403 4596 4406
rect 4770 4405 4773 4413
rect 794 4393 804 4396
rect 978 4393 1012 4396
rect 1026 4393 1036 4396
rect 1138 4393 1164 4396
rect 2858 4393 2884 4396
rect 38 4367 4829 4373
rect 2218 4343 2229 4346
rect 2794 4343 2820 4346
rect 2842 4343 2860 4346
rect 2930 4343 2948 4346
rect 2226 4336 2229 4343
rect 188 4333 205 4336
rect 116 4323 141 4326
rect 186 4323 204 4326
rect 234 4325 237 4336
rect 250 4333 276 4336
rect 556 4333 589 4336
rect 484 4323 509 4326
rect 578 4323 596 4326
rect 626 4325 629 4336
rect 674 4333 764 4336
rect 956 4333 973 4336
rect 996 4333 1052 4336
rect 668 4323 757 4326
rect 772 4323 789 4326
rect 860 4323 885 4326
rect 922 4323 948 4326
rect 1090 4325 1093 4336
rect 1122 4333 1156 4336
rect 1266 4333 1276 4336
rect 1300 4333 1317 4336
rect 1434 4326 1437 4335
rect 1500 4333 1509 4336
rect 1780 4333 1829 4336
rect 1852 4333 1908 4336
rect 1940 4333 1973 4336
rect 2010 4333 2036 4336
rect 2180 4333 2221 4336
rect 2226 4333 2244 4336
rect 2260 4333 2316 4336
rect 2332 4333 2381 4336
rect 2386 4333 2396 4336
rect 2412 4333 2429 4336
rect 2434 4333 2460 4336
rect 2530 4333 2540 4336
rect 2556 4333 2605 4336
rect 2634 4333 2660 4336
rect 2828 4333 2861 4336
rect 2874 4333 2900 4336
rect 2970 4333 3012 4336
rect 3036 4333 3077 4336
rect 3178 4326 3181 4335
rect 3514 4333 3564 4336
rect 3602 4333 3644 4336
rect 3818 4326 3821 4335
rect 3850 4333 3868 4336
rect 3962 4333 3988 4336
rect 4298 4333 4308 4336
rect 4538 4333 4556 4336
rect 4588 4333 4605 4336
rect 4636 4333 4685 4336
rect 1124 4323 1157 4326
rect 1202 4323 1228 4326
rect 1356 4323 1381 4326
rect 1412 4323 1437 4326
rect 1492 4323 1517 4326
rect 1578 4323 1596 4326
rect 1700 4323 1725 4326
rect 1762 4323 1772 4326
rect 1778 4323 1828 4326
rect 1860 4323 1877 4326
rect 1890 4323 1916 4326
rect 1988 4323 1997 4326
rect 2004 4323 2029 4326
rect 2082 4323 2108 4326
rect 2162 4323 2172 4326
rect 2210 4323 2236 4326
rect 2298 4323 2308 4326
rect 2354 4323 2388 4326
rect 2420 4323 2437 4326
rect 2498 4323 2532 4326
rect 2570 4323 2604 4326
rect 2636 4323 2645 4326
rect 2668 4323 2693 4326
rect 2836 4323 2853 4326
rect 2876 4323 2893 4326
rect 3028 4323 3069 4326
rect 3116 4323 3133 4326
rect 3172 4323 3181 4326
rect 3194 4323 3228 4326
rect 3444 4323 3461 4326
rect 3572 4323 3621 4326
rect 3626 4323 3652 4326
rect 3740 4323 3765 4326
rect 3796 4323 3821 4326
rect 3828 4323 3861 4326
rect 3922 4323 3948 4326
rect 4026 4323 4036 4326
rect 4066 4323 4092 4326
rect 4130 4323 4148 4326
rect 4322 4323 4340 4326
rect 4546 4323 4564 4326
rect 4594 4323 4628 4326
rect 1076 4313 1085 4316
rect 1810 4313 1813 4323
rect 2924 4313 2941 4316
rect 14 4267 4853 4273
rect 1076 4223 1101 4226
rect 2868 4223 2893 4226
rect 2924 4223 2949 4226
rect 2986 4223 3052 4226
rect 4250 4223 4260 4226
rect 4284 4223 4293 4226
rect 108 4213 133 4216
rect 170 4213 204 4216
rect 210 4213 228 4216
rect 308 4213 333 4216
rect 402 4213 420 4216
rect 212 4203 229 4206
rect 380 4203 421 4206
rect 450 4203 453 4214
rect 564 4213 589 4216
rect 642 4213 677 4216
rect 570 4203 612 4206
rect 628 4203 669 4206
rect 674 4205 677 4213
rect 730 4213 740 4216
rect 786 4213 796 4216
rect 884 4213 909 4216
rect 946 4213 964 4216
rect 1020 4213 1029 4216
rect 1090 4213 1108 4216
rect 1140 4213 1157 4216
rect 1210 4213 1236 4216
rect 1442 4213 1484 4216
rect 1562 4213 1572 4216
rect 1634 4213 1644 4216
rect 1650 4213 1668 4216
rect 1674 4213 1700 4216
rect 1756 4213 1781 4216
rect 1826 4213 1844 4216
rect 730 4206 733 4213
rect 1874 4206 1877 4214
rect 1882 4213 1916 4216
rect 1922 4213 1940 4216
rect 1946 4213 1972 4216
rect 2108 4213 2157 4216
rect 2172 4213 2213 4216
rect 2330 4213 2340 4216
rect 2418 4213 2485 4216
rect 2634 4213 2644 4216
rect 2708 4213 2741 4216
rect 2836 4213 2845 4216
rect 2882 4213 2908 4216
rect 3140 4213 3189 4216
rect 3258 4213 3284 4216
rect 3388 4213 3396 4216
rect 3482 4213 3524 4216
rect 3586 4213 3604 4216
rect 3634 4213 3676 4216
rect 3682 4213 3700 4216
rect 3730 4213 3756 4216
rect 3860 4213 3885 4216
rect 3954 4213 3964 4216
rect 3994 4213 4020 4216
rect 4108 4213 4125 4216
rect 4164 4213 4181 4216
rect 4188 4213 4197 4216
rect 708 4203 733 4206
rect 946 4203 956 4206
rect 986 4203 1012 4206
rect 1034 4203 1052 4206
rect 1076 4203 1085 4206
rect 1138 4203 1164 4206
rect 1300 4203 1341 4206
rect 1492 4203 1509 4206
rect 1548 4203 1557 4206
rect 1586 4203 1604 4206
rect 1682 4203 1692 4206
rect 1818 4203 1852 4206
rect 1874 4203 1893 4206
rect 1996 4203 2021 4206
rect 2050 4203 2100 4206
rect 2146 4203 2164 4206
rect 2314 4203 2332 4206
rect 2626 4203 2652 4206
rect 2674 4203 2700 4206
rect 2874 4203 2900 4206
rect 2924 4203 2957 4206
rect 2964 4203 2973 4206
rect 2978 4203 3052 4206
rect 3076 4203 3109 4206
rect 3154 4203 3172 4206
rect 3194 4203 3228 4206
rect 3260 4203 3277 4206
rect 3292 4203 3365 4206
rect 3412 4203 3437 4206
rect 3498 4203 3516 4206
rect 3530 4203 3596 4206
rect 3628 4203 3653 4206
rect 3682 4205 3685 4213
rect 3852 4203 3869 4206
rect 3932 4203 3957 4206
rect 4178 4205 4181 4213
rect 4298 4203 4301 4214
rect 4346 4213 4372 4216
rect 4508 4213 4517 4216
rect 4588 4214 4597 4216
rect 4324 4203 4357 4206
rect 4514 4205 4517 4213
rect 4586 4213 4597 4214
rect 4586 4203 4589 4213
rect 4772 4203 4781 4206
rect 970 4193 1004 4196
rect 2930 4193 2956 4196
rect 3634 4183 3637 4203
rect 38 4167 4829 4173
rect 1906 4153 1957 4156
rect 834 4143 868 4146
rect 1026 4143 1052 4146
rect 2722 4143 2756 4146
rect 2770 4143 2868 4146
rect 132 4133 165 4136
rect 188 4133 204 4136
rect 218 4133 237 4136
rect 420 4133 461 4136
rect 564 4133 573 4136
rect 586 4133 604 4136
rect 658 4133 668 4136
rect 866 4133 876 4136
rect 932 4133 988 4136
rect 1012 4133 1021 4136
rect 1050 4133 1060 4136
rect 1066 4133 1085 4136
rect 1090 4133 1108 4136
rect 1146 4133 1172 4136
rect 1282 4133 1316 4136
rect 1346 4133 1380 4136
rect 1402 4133 1420 4136
rect 1452 4133 1485 4136
rect 1586 4133 1620 4136
rect 1652 4133 1693 4136
rect 1812 4133 1861 4136
rect 1884 4133 1964 4136
rect 1996 4133 2044 4136
rect 2066 4133 2117 4136
rect 2306 4133 2396 4136
rect 2490 4133 2525 4136
rect 2548 4133 2597 4136
rect 2764 4133 2869 4136
rect 2876 4133 2901 4136
rect 2906 4133 2940 4136
rect 2964 4133 2989 4136
rect 3020 4133 3037 4136
rect 3084 4133 3109 4136
rect 3154 4133 3164 4136
rect 3196 4133 3229 4136
rect 234 4126 237 4133
rect 114 4123 124 4126
rect 202 4123 229 4126
rect 234 4123 244 4126
rect 348 4123 373 4126
rect 434 4123 460 4126
rect 492 4123 501 4126
rect 506 4123 540 4126
rect 556 4123 565 4126
rect 578 4123 596 4126
rect 628 4123 637 4126
rect 730 4123 740 4126
rect 770 4123 796 4126
rect 884 4123 893 4126
rect 898 4123 908 4126
rect 940 4123 965 4126
rect 970 4123 996 4126
rect 1066 4125 1069 4133
rect 1074 4123 1116 4126
rect 1218 4123 1244 4126
rect 1338 4123 1413 4126
rect 1444 4123 1453 4126
rect 1524 4123 1549 4126
rect 1644 4123 1685 4126
rect 1732 4123 1757 4126
rect 1794 4123 1804 4126
rect 1810 4123 1860 4126
rect 1892 4123 1901 4126
rect 1954 4123 1972 4126
rect 2002 4123 2036 4126
rect 2066 4125 2069 4133
rect 2074 4123 2132 4126
rect 2162 4123 2188 4126
rect 2484 4123 2517 4126
rect 2522 4125 2525 4133
rect 3346 4126 3349 4135
rect 3450 4133 3468 4136
rect 3636 4133 3645 4136
rect 3754 4126 3757 4135
rect 3770 4133 3812 4136
rect 3844 4133 3885 4136
rect 3890 4133 3900 4136
rect 3916 4133 3965 4136
rect 4162 4126 4165 4135
rect 4228 4133 4237 4136
rect 4324 4133 4365 4136
rect 4586 4126 4589 4136
rect 4594 4133 4628 4136
rect 4660 4133 4677 4136
rect 2556 4123 2573 4126
rect 2612 4123 2621 4126
rect 2772 4123 2861 4126
rect 2884 4123 2893 4126
rect 2956 4123 2997 4126
rect 3090 4123 3116 4126
rect 3324 4123 3349 4126
rect 3356 4123 3365 4126
rect 3594 4123 3612 4126
rect 3644 4123 3653 4126
rect 3692 4123 3717 4126
rect 3748 4123 3757 4126
rect 3764 4123 3789 4126
rect 3794 4123 3820 4126
rect 3866 4123 3892 4126
rect 4010 4123 4044 4126
rect 4092 4123 4117 4126
rect 4148 4123 4165 4126
rect 4172 4123 4189 4126
rect 4346 4123 4380 4126
rect 4586 4125 4613 4126
rect 4588 4123 4613 4125
rect 4626 4123 4636 4126
rect 1012 4113 1037 4116
rect 1132 4113 1165 4116
rect 1290 4113 1316 4116
rect 2970 4113 2996 4116
rect 3522 4113 3556 4116
rect 3580 4113 3605 4116
rect 14 4067 4853 4073
rect 898 4043 973 4046
rect 1236 4023 1245 4026
rect 2884 4023 2909 4026
rect 2938 4023 2972 4026
rect 3436 4023 3445 4026
rect 4354 4023 4364 4026
rect 4378 4023 4388 4026
rect 108 4013 117 4016
rect 164 4013 173 4016
rect 242 4013 268 4016
rect 306 4013 324 4016
rect 354 4013 380 4016
rect 468 4013 493 4016
rect 524 4013 541 4016
rect 588 4013 620 4016
rect 652 4013 685 4016
rect 724 4013 749 4016
rect 804 4013 813 4016
rect 860 4013 877 4016
rect 892 4013 973 4016
rect 988 4013 1037 4016
rect 1082 4013 1132 4016
rect 1170 4013 1220 4016
rect 1276 4013 1293 4016
rect 1322 4013 1421 4016
rect 1452 4013 1525 4016
rect 1572 4013 1597 4016
rect 1628 4013 1653 4016
rect 1690 4013 1789 4016
rect 1804 4013 1821 4016
rect 2042 4013 2060 4016
rect 2242 4013 2252 4016
rect 2290 4013 2332 4016
rect 2370 4013 2380 4016
rect 2426 4013 2452 4016
rect 2482 4013 2508 4016
rect 2546 4013 2588 4016
rect 2626 4013 2676 4016
rect 2708 4013 2717 4016
rect 2818 4013 2868 4016
rect 2988 4013 3005 4016
rect 3324 4013 3341 4016
rect 3450 4013 3460 4016
rect 3466 4013 3508 4016
rect 3674 4013 3708 4016
rect 3844 4013 3861 4016
rect 3874 4013 3900 4016
rect 3922 4013 3940 4016
rect 4132 4013 4157 4016
rect 4188 4013 4197 4016
rect 4204 4013 4229 4016
rect 4234 4013 4244 4016
rect 4394 4013 4428 4016
rect 4492 4013 4517 4016
rect 4548 4013 4557 4016
rect 4594 4013 4620 4016
rect 4674 4013 4716 4016
rect 306 4006 309 4013
rect 186 4003 204 4006
rect 250 4003 276 4006
rect 292 4003 309 4006
rect 538 4006 541 4013
rect 538 4003 564 4006
rect 580 4003 589 4006
rect 602 4003 628 4006
rect 658 4003 700 4006
rect 884 4003 917 4006
rect 1034 4003 1037 4013
rect 1322 4006 1325 4013
rect 2426 4006 2429 4013
rect 1042 4003 1052 4006
rect 1068 4003 1093 4006
rect 1106 4003 1140 4006
rect 1156 4003 1212 4006
rect 1250 4003 1260 4006
rect 1316 4003 1325 4006
rect 1330 4003 1348 4006
rect 1402 4003 1428 4006
rect 1634 4003 1660 4006
rect 2042 4003 2052 4006
rect 2178 4003 2196 4006
rect 2250 4003 2260 4006
rect 2276 4003 2309 4006
rect 2348 4003 2373 4006
rect 2378 4003 2388 4006
rect 2404 4003 2429 4006
rect 2554 4003 2596 4006
rect 2612 4003 2669 4006
rect 2674 4003 2684 4006
rect 2706 4003 2756 4006
rect 2842 4003 2860 4006
rect 2884 4003 2893 4006
rect 2898 4003 2972 4006
rect 2996 4003 3029 4006
rect 3130 4003 3164 4006
rect 3338 4005 3341 4013
rect 3396 4003 3405 4006
rect 3466 4005 3469 4013
rect 3602 4003 3636 4006
rect 3668 4003 3693 4006
rect 3724 4003 3741 4006
rect 3858 4005 3861 4013
rect 3956 4003 3973 4006
rect 4194 4005 4197 4013
rect 4210 4003 4236 4006
rect 4282 4003 4308 4006
rect 4324 4003 4357 4006
rect 4436 4003 4453 4006
rect 4588 4003 4605 4006
rect 4610 4003 4628 4006
rect 4644 4003 4653 4006
rect 4724 4003 4781 4006
rect 866 3993 876 3996
rect 38 3967 4829 3973
rect 2882 3943 2908 3946
rect 476 3933 493 3936
rect 516 3933 564 3936
rect 596 3933 637 3936
rect 642 3933 652 3936
rect 674 3933 708 3936
rect 884 3933 909 3936
rect 922 3933 940 3936
rect 1234 3933 1260 3936
rect 1284 3933 1325 3936
rect 1426 3933 1476 3936
rect 1674 3933 1692 3936
rect 1828 3933 1908 3936
rect 1940 3933 2012 3936
rect 2028 3933 2061 3936
rect 2114 3933 2148 3936
rect 2234 3933 2260 3936
rect 2292 3933 2309 3936
rect 2346 3933 2396 3936
rect 2410 3933 2452 3936
rect 2530 3933 2556 3936
rect 2572 3933 2597 3936
rect 2842 3926 2845 3935
rect 2868 3933 2877 3936
rect 2916 3933 2949 3936
rect 3058 3926 3061 3935
rect 3106 3933 3124 3936
rect 3156 3933 3189 3936
rect 3746 3933 3844 3936
rect 3876 3933 3893 3936
rect 4274 3933 4284 3936
rect 4314 3933 4340 3936
rect 4482 3926 4485 3935
rect 4498 3933 4532 3936
rect 4564 3933 4581 3936
rect 4668 3933 4685 3936
rect 108 3923 133 3926
rect 220 3923 245 3926
rect 276 3923 301 3926
rect 388 3923 413 3926
rect 450 3923 468 3926
rect 524 3923 557 3926
rect 588 3923 613 3926
rect 676 3923 685 3926
rect 716 3923 741 3926
rect 786 3923 812 3926
rect 850 3923 876 3926
rect 890 3923 932 3926
rect 1130 3923 1140 3926
rect 1276 3923 1301 3926
rect 1458 3923 1484 3926
rect 1572 3923 1589 3926
rect 1634 3923 1669 3926
rect 1714 3923 1804 3926
rect 1836 3923 1893 3926
rect 1994 3923 2004 3926
rect 2100 3923 2109 3926
rect 2122 3923 2140 3926
rect 2172 3923 2181 3926
rect 2284 3923 2293 3926
rect 2348 3923 2357 3926
rect 2404 3923 2429 3926
rect 2460 3923 2485 3926
rect 2508 3923 2541 3926
rect 2756 3923 2765 3926
rect 2812 3923 2845 3926
rect 2988 3923 3013 3926
rect 3044 3923 3061 3926
rect 3148 3923 3173 3926
rect 3386 3923 3396 3926
rect 3500 3923 3541 3926
rect 3610 3923 3620 3926
rect 3650 3923 3676 3926
rect 3732 3923 3741 3926
rect 3826 3923 3852 3926
rect 3940 3923 3957 3926
rect 4044 3923 4061 3926
rect 4156 3923 4181 3926
rect 4212 3923 4229 3926
rect 4234 3923 4244 3926
rect 4274 3923 4292 3926
rect 4476 3923 4485 3926
rect 4498 3923 4540 3926
rect 4570 3923 4612 3926
rect 4634 3923 4644 3926
rect 1250 3913 1260 3916
rect 2868 3913 2901 3916
rect 1946 3883 1997 3886
rect 14 3867 4853 3873
rect 1108 3823 1157 3826
rect 2772 3823 2789 3826
rect 2860 3823 2869 3826
rect 2882 3823 2892 3826
rect 2938 3823 2956 3826
rect 4346 3823 4356 3826
rect 116 3813 125 3816
rect 172 3813 189 3816
rect 178 3803 204 3806
rect 226 3803 229 3814
rect 242 3813 252 3816
rect 260 3803 293 3806
rect 322 3803 325 3814
rect 364 3813 389 3816
rect 596 3813 613 3816
rect 634 3813 652 3816
rect 684 3813 693 3816
rect 714 3813 732 3816
rect 770 3813 788 3816
rect 826 3813 876 3816
rect 908 3813 949 3816
rect 972 3813 997 3816
rect 1036 3813 1085 3816
rect 1180 3813 1197 3816
rect 1348 3813 1365 3816
rect 1404 3813 1437 3816
rect 1524 3813 1541 3816
rect 1700 3813 1725 3816
rect 1754 3813 1788 3816
rect 1794 3813 1828 3816
rect 1860 3813 1885 3816
rect 1938 3813 1948 3816
rect 1986 3813 2012 3816
rect 2108 3813 2133 3816
rect 2164 3813 2181 3816
rect 2186 3813 2292 3816
rect 2354 3813 2364 3816
rect 2426 3813 2436 3816
rect 2498 3813 2524 3816
rect 2556 3813 2573 3816
rect 2580 3813 2613 3816
rect 2812 3813 2829 3816
rect 714 3806 717 3813
rect 436 3803 485 3806
rect 508 3803 572 3806
rect 604 3803 645 3806
rect 676 3803 717 3806
rect 900 3803 909 3806
rect 964 3803 997 3806
rect 1034 3803 1084 3806
rect 1108 3803 1117 3806
rect 1234 3803 1252 3806
rect 1276 3803 1309 3806
rect 1434 3805 1437 3813
rect 2866 3806 2869 3823
rect 3036 3813 3045 3816
rect 3050 3813 3076 3816
rect 3106 3813 3132 3816
rect 3170 3813 3212 3816
rect 3282 3813 3292 3816
rect 3356 3813 3405 3816
rect 3484 3813 3517 3816
rect 3522 3813 3589 3816
rect 1482 3803 1500 3806
rect 1532 3803 1581 3806
rect 1634 3803 1684 3806
rect 1706 3803 1732 3806
rect 1796 3803 1829 3806
rect 2250 3803 2300 3806
rect 2322 3803 2356 3806
rect 2492 3803 2525 3806
rect 2554 3803 2572 3806
rect 2714 3803 2748 3806
rect 2772 3803 2797 3806
rect 2810 3803 2836 3806
rect 2866 3803 2892 3806
rect 2922 3803 2956 3806
rect 2980 3803 3005 3806
rect 3050 3803 3053 3813
rect 3402 3806 3405 3813
rect 3522 3806 3525 3813
rect 3866 3806 3869 3816
rect 3874 3813 3892 3816
rect 3924 3813 3941 3816
rect 3978 3813 4004 3816
rect 4010 3813 4052 3816
rect 4082 3813 4108 3816
rect 4114 3813 4156 3816
rect 4250 3813 4260 3816
rect 4292 3813 4309 3816
rect 4412 3813 4421 3816
rect 4540 3813 4549 3816
rect 4596 3813 4605 3816
rect 3338 3803 3348 3806
rect 3402 3803 3460 3806
rect 3476 3803 3525 3806
rect 3572 3803 3613 3806
rect 3866 3803 3900 3806
rect 3922 3803 3940 3806
rect 3972 3803 3989 3806
rect 4034 3803 4044 3806
rect 4258 3803 4268 3806
rect 4610 3803 4628 3806
rect 4660 3803 4669 3806
rect 922 3793 956 3796
rect 970 3793 1020 3796
rect 2778 3793 2796 3796
rect 38 3767 4829 3773
rect 922 3743 948 3746
rect 1010 3743 1060 3746
rect 2746 3743 2796 3746
rect 2826 3743 2844 3746
rect 140 3733 173 3736
rect 218 3733 244 3736
rect 412 3733 445 3736
rect 660 3733 669 3736
rect 674 3733 724 3736
rect 970 3733 980 3736
rect 1050 3733 1068 3736
rect 1074 3733 1108 3736
rect 1132 3733 1188 3736
rect 100 3723 109 3726
rect 122 3723 132 3726
rect 162 3723 172 3726
rect 204 3723 221 3726
rect 242 3723 252 3726
rect 332 3723 357 3726
rect 394 3723 404 3726
rect 426 3723 444 3726
rect 476 3723 493 3726
rect 540 3723 557 3726
rect 596 3723 605 3726
rect 668 3723 693 3726
rect 732 3723 741 3726
rect 748 3723 773 3726
rect 820 3723 837 3726
rect 884 3723 893 3726
rect 970 3723 988 3726
rect 1074 3725 1077 3733
rect 1124 3723 1149 3726
rect 1210 3725 1213 3736
rect 1226 3733 1244 3736
rect 1258 3733 1300 3736
rect 1346 3733 1372 3736
rect 1396 3733 1429 3736
rect 1546 3726 1549 3735
rect 1562 3733 1612 3736
rect 1644 3733 1669 3736
rect 1948 3733 1989 3736
rect 1252 3723 1269 3726
rect 1468 3723 1493 3726
rect 1524 3723 1549 3726
rect 1724 3723 1749 3726
rect 1802 3723 1828 3726
rect 1874 3723 1884 3726
rect 1946 3723 1988 3726
rect 2018 3725 2021 3736
rect 2026 3723 2036 3726
rect 2076 3723 2101 3726
rect 2154 3725 2157 3736
rect 2250 3733 2292 3736
rect 2324 3733 2333 3736
rect 2530 3733 2564 3736
rect 2594 3733 2612 3736
rect 2804 3733 2845 3736
rect 2852 3733 2877 3736
rect 2330 3726 2333 3733
rect 2930 3726 2933 3735
rect 2946 3733 2972 3736
rect 3068 3733 3077 3736
rect 3578 3726 3581 3735
rect 3738 3733 3772 3736
rect 3786 3733 3796 3736
rect 3818 3733 3836 3736
rect 4170 3726 4173 3736
rect 4236 3733 4245 3736
rect 4428 3733 4445 3736
rect 4474 3733 4484 3736
rect 4516 3733 4533 3736
rect 4538 3733 4556 3736
rect 4572 3733 4581 3736
rect 2258 3723 2300 3726
rect 2330 3723 2372 3726
rect 2402 3723 2428 3726
rect 2466 3723 2556 3726
rect 2588 3723 2605 3726
rect 2620 3723 2645 3726
rect 2900 3723 2933 3726
rect 2940 3723 2973 3726
rect 3018 3723 3044 3726
rect 3060 3723 3069 3726
rect 3530 3723 3572 3726
rect 3578 3723 3636 3726
rect 3666 3723 3692 3726
rect 3786 3723 3829 3726
rect 3914 3723 3964 3726
rect 3994 3723 4020 3726
rect 4170 3723 4277 3726
rect 4370 3723 4420 3726
rect 4460 3723 4485 3726
rect 218 3703 221 3723
rect 1004 3713 1037 3716
rect 1098 3713 1108 3716
rect 1282 3713 1300 3716
rect 1346 3713 1372 3716
rect 2954 3713 2972 3716
rect 3330 3713 3348 3716
rect 3372 3713 3413 3716
rect 3356 3703 3373 3706
rect 14 3667 4853 3673
rect 1234 3623 1244 3626
rect 1332 3623 1349 3626
rect 2556 3623 2573 3626
rect 2812 3623 2829 3626
rect 2866 3623 2892 3626
rect 2914 3616 2917 3625
rect 3300 3623 3349 3626
rect 4108 3623 4117 3626
rect 164 3613 181 3616
rect 554 3613 564 3616
rect 892 3613 909 3616
rect 948 3613 965 3616
rect 1002 3613 1012 3616
rect 1018 3613 1052 3616
rect 1084 3613 1093 3616
rect 1138 3613 1164 3616
rect 1260 3613 1277 3616
rect 1282 3613 1324 3616
rect 1426 3613 1436 3616
rect 1540 3613 1557 3616
rect 1578 3613 1612 3616
rect 1716 3613 1733 3616
rect 1740 3613 1749 3616
rect 1770 3613 1780 3616
rect 1828 3613 1845 3616
rect 1900 3614 1948 3616
rect 1900 3613 1949 3614
rect 1986 3613 2028 3616
rect 2138 3613 2172 3616
rect 2300 3613 2325 3616
rect 2338 3613 2348 3616
rect 2466 3613 2492 3616
rect 2530 3613 2540 3616
rect 2786 3613 2796 3616
rect 2852 3613 2861 3616
rect 2882 3613 2917 3616
rect 2932 3613 2949 3616
rect 3020 3613 3045 3616
rect 3082 3613 3101 3616
rect 3154 3613 3204 3616
rect 3322 3613 3356 3616
rect 3452 3613 3485 3616
rect 3498 3613 3548 3616
rect 3676 3613 3701 3616
rect 3732 3613 3741 3616
rect 906 3606 909 3613
rect 498 3603 556 3606
rect 906 3603 924 3606
rect 940 3603 973 3606
rect 1020 3603 1037 3606
rect 1082 3603 1101 3606
rect 1140 3603 1165 3606
rect 1188 3603 1197 3606
rect 1234 3603 1244 3606
rect 1306 3603 1316 3606
rect 1482 3603 1516 3606
rect 1548 3603 1605 3606
rect 1730 3605 1733 3613
rect 1796 3603 1821 3606
rect 1836 3603 1869 3606
rect 1946 3603 1949 3613
rect 2322 3606 2325 3613
rect 1986 3603 2036 3606
rect 2052 3603 2100 3606
rect 2132 3603 2165 3606
rect 2180 3603 2189 3606
rect 2322 3603 2356 3606
rect 2778 3603 2788 3606
rect 2844 3603 2893 3606
rect 2940 3603 2981 3606
rect 3082 3603 3116 3606
rect 3148 3603 3197 3606
rect 3212 3603 3253 3606
rect 3380 3603 3421 3606
rect 3514 3603 3540 3606
rect 3754 3603 3757 3614
rect 3788 3613 3877 3616
rect 3882 3613 3949 3616
rect 3980 3613 4044 3616
rect 4236 3613 4245 3616
rect 4250 3613 4276 3616
rect 4322 3613 4356 3616
rect 4490 3613 4508 3616
rect 4538 3613 4572 3616
rect 4634 3613 4660 3616
rect 4690 3613 4748 3616
rect 3780 3603 3789 3606
rect 3794 3603 3797 3613
rect 3994 3603 4036 3606
rect 4132 3603 4141 3606
rect 4274 3603 4284 3606
rect 4300 3603 4341 3606
rect 4482 3603 4500 3606
rect 4620 3603 4645 3606
rect 4684 3603 4741 3606
rect 4756 3603 4773 3606
rect 2826 3593 2836 3596
rect 38 3567 4829 3573
rect 1210 3543 1220 3546
rect 148 3533 189 3536
rect 212 3533 229 3536
rect 340 3533 389 3536
rect 412 3533 492 3536
rect 508 3533 605 3536
rect 636 3533 661 3536
rect 706 3533 764 3536
rect 852 3533 869 3536
rect 916 3533 925 3536
rect 1202 3533 1228 3536
rect 1258 3533 1284 3536
rect 1314 3533 1356 3536
rect 1378 3526 1381 3534
rect 1386 3533 1436 3536
rect 1514 3533 1532 3536
rect 1564 3533 1605 3536
rect 1796 3533 1837 3536
rect 1986 3533 1996 3536
rect 2042 3533 2052 3536
rect 2162 3533 2188 3536
rect 2210 3526 2213 3536
rect 2348 3533 2357 3536
rect 2380 3533 2389 3536
rect 2522 3533 2612 3536
rect 2628 3533 2669 3536
rect 2674 3533 2684 3536
rect 2706 3533 2732 3536
rect 2754 3533 2788 3536
rect 2812 3533 2861 3536
rect 2874 3533 2884 3536
rect 2914 3533 2948 3536
rect 3026 3533 3044 3536
rect 3356 3533 3413 3536
rect 3522 3533 3532 3536
rect 3602 3533 3612 3536
rect 3626 3533 3692 3536
rect 122 3523 140 3526
rect 338 3523 388 3526
rect 420 3523 429 3526
rect 442 3523 484 3526
rect 522 3523 612 3526
rect 642 3523 668 3526
rect 788 3523 797 3526
rect 834 3523 844 3526
rect 882 3523 900 3526
rect 1188 3523 1197 3526
rect 1300 3523 1325 3526
rect 1378 3523 1444 3526
rect 1556 3523 1620 3526
rect 1650 3523 1700 3526
rect 1754 3523 1772 3526
rect 1810 3523 1844 3526
rect 1850 3523 1892 3526
rect 1938 3523 1948 3526
rect 1986 3523 2004 3526
rect 2098 3523 2124 3526
rect 2210 3525 2237 3526
rect 2212 3523 2237 3525
rect 2276 3523 2293 3526
rect 2484 3523 2549 3526
rect 2570 3523 2604 3526
rect 2642 3523 2676 3526
rect 2786 3523 2796 3526
rect 2900 3523 2949 3526
rect 3082 3523 3116 3526
rect 3122 3523 3172 3526
rect 3322 3523 3332 3526
rect 3364 3523 3389 3526
rect 3452 3523 3469 3526
rect 3508 3523 3517 3526
rect 916 3513 965 3516
rect 1314 3513 1356 3516
rect 2812 3513 2869 3516
rect 2914 3513 2948 3516
rect 3202 3513 3244 3516
rect 3268 3513 3325 3516
rect 3522 3506 3525 3533
rect 3754 3523 3764 3526
rect 3794 3525 3797 3536
rect 3986 3526 3989 3534
rect 4274 3526 4277 3534
rect 4290 3533 4316 3536
rect 3980 3523 3989 3526
rect 4212 3523 4229 3526
rect 4268 3523 4277 3526
rect 4290 3523 4324 3526
rect 4530 3523 4533 3534
rect 3514 3503 3525 3506
rect 14 3467 4853 3473
rect 1076 3423 1125 3426
rect 2586 3423 2613 3426
rect 2810 3423 2853 3426
rect 2586 3416 2589 3423
rect 2850 3416 2853 3423
rect 116 3413 125 3416
rect 172 3413 197 3416
rect 316 3413 341 3416
rect 378 3413 404 3416
rect 468 3413 477 3416
rect 482 3413 493 3416
rect 516 3413 533 3416
rect 636 3413 645 3416
rect 724 3413 741 3416
rect 804 3413 813 3416
rect 860 3413 909 3416
rect 988 3413 1029 3416
rect 1164 3413 1173 3416
rect 1220 3413 1237 3416
rect 1274 3413 1300 3416
rect 1372 3413 1389 3416
rect 1428 3413 1453 3416
rect 1484 3413 1493 3416
rect 1562 3413 1572 3416
rect 1740 3413 1749 3416
rect 1794 3413 1812 3416
rect 1842 3413 1868 3416
rect 1948 3413 1973 3416
rect 2010 3413 2028 3416
rect 2092 3413 2117 3416
rect 2154 3413 2180 3416
rect 2306 3413 2340 3416
rect 2378 3413 2388 3416
rect 2476 3413 2509 3416
rect 2548 3413 2565 3416
rect 2580 3413 2589 3416
rect 2594 3413 2660 3416
rect 2706 3413 2716 3416
rect 2804 3413 2845 3416
rect 2850 3413 2868 3416
rect 2964 3413 2997 3416
rect 3100 3413 3109 3416
rect 3268 3413 3285 3416
rect 3436 3413 3461 3416
rect 3492 3413 3501 3416
rect 3676 3413 3709 3416
rect 3740 3413 3781 3416
rect 3826 3413 3844 3416
rect 482 3406 485 3413
rect 178 3403 220 3406
rect 410 3403 444 3406
rect 476 3403 485 3406
rect 490 3403 508 3406
rect 668 3403 685 3406
rect 690 3403 716 3406
rect 1034 3403 1052 3406
rect 1082 3403 1140 3406
rect 1162 3403 1212 3406
rect 1338 3403 1356 3406
rect 1490 3405 1493 3413
rect 3874 3406 3877 3426
rect 4180 3413 4189 3416
rect 4410 3413 4420 3416
rect 4426 3413 4453 3416
rect 4410 3406 4413 3413
rect 2036 3403 2053 3406
rect 2412 3403 2453 3406
rect 2468 3403 2509 3406
rect 2514 3403 2524 3406
rect 2540 3403 2557 3406
rect 2658 3403 2668 3406
rect 2684 3403 2709 3406
rect 2740 3403 2789 3406
rect 2802 3403 2860 3406
rect 2890 3403 2940 3406
rect 3514 3403 3532 3406
rect 3578 3403 3652 3406
rect 3690 3403 3716 3406
rect 3770 3403 3836 3406
rect 3868 3403 3893 3406
rect 3994 3403 4020 3406
rect 4194 3403 4212 3406
rect 4322 3403 4356 3406
rect 4372 3403 4413 3406
rect 4426 3405 4429 3413
rect 4458 3403 4461 3414
rect 4506 3406 4509 3416
rect 4658 3413 4676 3416
rect 4706 3413 4748 3416
rect 4484 3403 4509 3406
rect 4658 3403 4668 3406
rect 4700 3403 4741 3406
rect 4756 3403 4781 3406
rect 410 3393 437 3396
rect 674 3393 708 3396
rect 874 3393 972 3396
rect 2426 3393 2460 3396
rect 2746 3393 2788 3396
rect 38 3367 4829 3373
rect 1178 3343 1212 3346
rect 204 3333 229 3336
rect 266 3333 300 3336
rect 370 3333 388 3336
rect 404 3333 437 3336
rect 500 3333 509 3336
rect 658 3333 700 3336
rect 786 3333 804 3336
rect 996 3333 1029 3336
rect 1076 3333 1148 3336
rect 1210 3333 1220 3336
rect 1226 3333 1276 3336
rect 1306 3333 1356 3336
rect 1380 3333 1453 3336
rect 1492 3333 1509 3336
rect 1514 3333 1548 3336
rect 1578 3333 1628 3336
rect 1660 3333 1717 3336
rect 1748 3333 1781 3336
rect 1820 3333 1837 3336
rect 1876 3333 1925 3336
rect 2146 3333 2164 3336
rect 2180 3333 2236 3336
rect 2258 3333 2284 3336
rect 146 3323 156 3326
rect 370 3323 380 3326
rect 412 3323 476 3326
rect 588 3323 605 3326
rect 900 3323 925 3326
rect 962 3323 988 3326
rect 994 3323 1052 3326
rect 1228 3323 1261 3326
rect 1298 3323 1325 3326
rect 1372 3323 1381 3326
rect 1458 3323 1468 3326
rect 1722 3323 1732 3326
rect 1842 3323 1868 3326
rect 1922 3323 1925 3333
rect 2690 3326 2693 3334
rect 2706 3333 2748 3336
rect 2890 3333 2900 3336
rect 2922 3326 2925 3334
rect 2930 3333 2972 3336
rect 3002 3333 3060 3336
rect 3084 3333 3125 3336
rect 3164 3333 3173 3336
rect 1996 3323 2005 3326
rect 2058 3323 2156 3326
rect 2266 3323 2292 3326
rect 2412 3323 2421 3326
rect 2540 3323 2549 3326
rect 2594 3323 2612 3326
rect 2666 3323 2693 3326
rect 2700 3323 2749 3326
rect 2852 3323 2861 3326
rect 2922 3323 2933 3326
rect 3130 3323 3140 3326
rect 3170 3323 3212 3326
rect 3266 3323 3269 3334
rect 3322 3333 3332 3336
rect 3476 3333 3485 3336
rect 3498 3333 3516 3336
rect 3666 3326 3669 3334
rect 3876 3333 3885 3336
rect 3940 3333 3949 3336
rect 4186 3333 4228 3336
rect 4258 3333 4268 3336
rect 4290 3333 4317 3336
rect 3306 3323 3340 3326
rect 3490 3323 3524 3326
rect 3596 3323 3621 3326
rect 3652 3323 3669 3326
rect 3810 3323 3852 3326
rect 3898 3323 3932 3326
rect 4178 3323 4236 3326
rect 4242 3323 4260 3326
rect 4290 3325 4293 3333
rect 4338 3325 4341 3336
rect 4370 3333 4388 3336
rect 4476 3333 4501 3336
rect 4516 3333 4549 3336
rect 4588 3333 4613 3336
rect 4628 3333 4637 3336
rect 4450 3323 4460 3326
rect 4482 3323 4508 3326
rect 4594 3323 4620 3326
rect 4732 3323 4741 3326
rect 1172 3313 1205 3316
rect 1298 3315 1301 3323
rect 1306 3313 1356 3316
rect 2884 3313 2893 3316
rect 2930 3313 2933 3323
rect 3010 3313 3060 3316
rect 3378 3313 3388 3316
rect 3412 3313 3445 3316
rect 4348 3313 4365 3316
rect 3396 3303 3413 3306
rect 14 3267 4853 3273
rect 3474 3233 3493 3236
rect 964 3223 1005 3226
rect 1306 3223 1332 3226
rect 2418 3223 2437 3226
rect 2556 3223 2581 3226
rect 2970 3223 2980 3226
rect 3354 3223 3388 3226
rect 2418 3216 2421 3223
rect 108 3213 133 3216
rect 178 3213 188 3216
rect 260 3213 269 3216
rect 306 3213 332 3216
rect 412 3213 421 3216
rect 516 3213 549 3216
rect 562 3206 565 3214
rect 618 3213 660 3216
rect 706 3213 772 3216
rect 804 3213 829 3216
rect 850 3213 877 3216
rect 922 3213 948 3216
rect 1028 3213 1069 3216
rect 180 3203 189 3206
rect 212 3203 221 3206
rect 546 3203 565 3206
rect 588 3203 613 3206
rect 618 3183 621 3213
rect 874 3206 877 3213
rect 1074 3206 1077 3214
rect 1162 3213 1172 3216
rect 1204 3213 1213 3216
rect 1268 3213 1277 3216
rect 1348 3213 1381 3216
rect 1452 3213 1461 3216
rect 1572 3213 1605 3216
rect 1708 3213 1717 3216
rect 1722 3213 1732 3216
rect 1770 3213 1796 3216
rect 1842 3213 1868 3216
rect 1898 3213 1908 3216
rect 1978 3213 2084 3216
rect 2348 3213 2357 3216
rect 2362 3213 2380 3216
rect 2412 3213 2421 3216
rect 2426 3213 2460 3216
rect 2490 3213 2540 3216
rect 2684 3213 2693 3216
rect 2924 3213 2933 3216
rect 3034 3213 3093 3216
rect 3138 3213 3148 3216
rect 3306 3213 3332 3216
rect 3474 3215 3477 3233
rect 3490 3226 3493 3233
rect 3490 3223 3532 3226
rect 3546 3223 3556 3226
rect 3562 3223 3596 3226
rect 3620 3223 3709 3226
rect 642 3203 652 3206
rect 770 3203 780 3206
rect 796 3203 869 3206
rect 874 3203 884 3206
rect 890 3203 940 3206
rect 1020 3203 1077 3206
rect 1100 3203 1117 3206
rect 1162 3203 1180 3206
rect 1196 3203 1205 3206
rect 1226 3203 1252 3206
rect 1276 3203 1285 3206
rect 1322 3203 1332 3206
rect 1356 3203 1421 3206
rect 1460 3203 1541 3206
rect 1586 3203 1692 3206
rect 1882 3203 1916 3206
rect 2010 3203 2092 3206
rect 2108 3203 2181 3206
rect 2194 3203 2204 3206
rect 2250 3203 2260 3206
rect 2292 3203 2309 3206
rect 2418 3203 2452 3206
rect 2556 3203 2597 3206
rect 2604 3203 2645 3206
rect 2682 3203 2724 3206
rect 2922 3203 2980 3206
rect 3004 3203 3045 3206
rect 3060 3203 3101 3206
rect 3258 3203 3268 3206
rect 3340 3203 3365 3206
rect 3610 3203 3613 3214
rect 3732 3213 3789 3216
rect 3834 3213 3884 3216
rect 3930 3213 3948 3216
rect 4114 3213 4156 3216
rect 4204 3213 4229 3216
rect 4276 3213 4309 3216
rect 4578 3213 4676 3216
rect 4706 3213 4740 3216
rect 3714 3203 3724 3206
rect 3778 3203 3796 3206
rect 3908 3203 3941 3206
rect 3986 3203 4004 3206
rect 4036 3203 4045 3206
rect 4050 3203 4084 3206
rect 4164 3203 4173 3206
rect 4242 3203 4252 3206
rect 4268 3203 4277 3206
rect 4594 3203 4668 3206
rect 818 3193 876 3196
rect 994 3193 1012 3196
rect 1042 3193 1069 3196
rect 2562 3193 2596 3196
rect 2834 3193 2908 3196
rect 38 3167 4829 3173
rect 2842 3143 2852 3146
rect 2866 3143 2876 3146
rect 180 3133 197 3136
rect 274 3133 284 3136
rect 338 3133 356 3136
rect 378 3133 412 3136
rect 434 3133 468 3136
rect 548 3133 573 3136
rect 578 3133 588 3136
rect 604 3133 613 3136
rect 770 3133 796 3136
rect 812 3133 892 3136
rect 916 3133 965 3136
rect 1012 3133 1100 3136
rect 1124 3133 1197 3136
rect 1210 3133 1268 3136
rect 1292 3133 1317 3136
rect 1322 3133 1348 3136
rect 108 3123 133 3126
rect 172 3123 181 3126
rect 186 3123 196 3126
rect 228 3123 253 3126
rect 266 3123 276 3126
rect 380 3123 405 3126
rect 498 3123 540 3126
rect 546 3123 580 3126
rect 684 3123 709 3126
rect 740 3123 781 3126
rect 820 3123 829 3126
rect 882 3123 900 3126
rect 922 3123 988 3126
rect 1194 3123 1197 3133
rect 1370 3126 1373 3135
rect 1418 3133 1428 3136
rect 1508 3133 1549 3136
rect 2010 3133 2020 3136
rect 2036 3133 2053 3136
rect 2106 3133 2116 3136
rect 2154 3133 2196 3136
rect 2474 3133 2509 3136
rect 2532 3133 2541 3136
rect 2658 3133 2668 3136
rect 2684 3133 2701 3136
rect 1370 3123 1436 3126
rect 1450 3123 1549 3126
rect 1580 3123 1605 3126
rect 1988 3123 2005 3126
rect 2074 3123 2124 3126
rect 2212 3123 2221 3126
rect 2260 3123 2269 3126
rect 2468 3123 2501 3126
rect 2506 3125 2509 3133
rect 2802 3126 2805 3135
rect 2828 3133 2845 3136
rect 2906 3133 2932 3136
rect 2962 3133 3004 3136
rect 3028 3133 3037 3136
rect 3042 3133 3068 3136
rect 3250 3126 3253 3135
rect 3532 3133 3549 3136
rect 3578 3133 3620 3136
rect 3810 3133 3844 3136
rect 2578 3123 2604 3126
rect 2642 3123 2660 3126
rect 2796 3123 2805 3126
rect 2948 3123 3005 3126
rect 3026 3123 3076 3126
rect 3220 3123 3253 3126
rect 3490 3123 3508 3126
rect 3540 3123 3621 3126
rect 3866 3125 3869 3136
rect 3884 3133 3909 3136
rect 4226 3133 4244 3136
rect 4282 3126 4285 3136
rect 4340 3133 4381 3136
rect 4562 3126 4565 3135
rect 4594 3133 4604 3136
rect 916 3113 949 3116
rect 1124 3113 1237 3116
rect 1258 3113 1268 3116
rect 1306 3113 1348 3116
rect 2828 3113 2837 3116
rect 2970 3113 3004 3116
rect 3370 3113 3396 3116
rect 3634 3113 3676 3116
rect 3690 3106 3693 3125
rect 3876 3123 3909 3126
rect 3954 3123 3996 3126
rect 4034 3123 4052 3126
rect 4140 3123 4157 3126
rect 4274 3123 4285 3126
rect 4306 3123 4316 3126
rect 4354 3123 4396 3126
rect 4548 3123 4565 3126
rect 4578 3123 4612 3126
rect 3700 3113 3773 3116
rect 3794 3113 3804 3116
rect 3690 3103 3741 3106
rect 14 3067 4853 3073
rect 900 3023 949 3026
rect 1338 3023 1348 3026
rect 2812 3023 2829 3026
rect 2930 3023 2956 3026
rect 2994 3023 3013 3026
rect 3410 3023 3428 3026
rect 3452 3023 3469 3026
rect 3010 3016 3013 3023
rect 148 3013 173 3016
rect 204 3013 245 3016
rect 340 3013 365 3016
rect 556 3013 589 3016
rect 618 3013 652 3016
rect 706 3013 732 3016
rect 586 3006 589 3013
rect 802 3006 805 3016
rect 820 3013 877 3016
rect 1002 3006 1005 3016
rect 1098 3013 1116 3016
rect 1242 3006 1245 3014
rect 1450 3013 1476 3016
rect 1546 3013 1572 3016
rect 1714 3013 1748 3016
rect 1780 3013 1813 3016
rect 1852 3013 1877 3016
rect 1890 3013 1916 3016
rect 1970 3013 1996 3016
rect 2194 3013 2204 3016
rect 2274 3013 2300 3016
rect 2410 3013 2421 3016
rect 2444 3013 2493 3016
rect 2532 3013 2541 3016
rect 2580 3013 2605 3016
rect 2642 3013 2668 3016
rect 2852 3013 2861 3016
rect 2972 3013 3005 3016
rect 3010 3013 3021 3016
rect 3130 3013 3156 3016
rect 3364 3013 3389 3016
rect 3508 3013 3533 3016
rect 3564 3013 3581 3016
rect 3692 3013 3709 3016
rect 3836 3013 3853 3016
rect 3964 3013 3989 3016
rect 4020 3013 4029 3016
rect 2410 3006 2413 3013
rect 146 3003 180 3006
rect 212 3003 253 3006
rect 412 3003 461 3006
rect 586 3003 644 3006
rect 740 3003 805 3006
rect 818 3003 876 3006
rect 900 3003 909 3006
rect 946 3003 964 3006
rect 1002 3003 1028 3006
rect 1188 3003 1245 3006
rect 1268 3003 1277 3006
rect 1282 3003 1348 3006
rect 1372 3003 1413 3006
rect 1514 3003 1564 3006
rect 1596 3003 1660 3006
rect 1692 3003 1725 3006
rect 1844 3003 1869 3006
rect 2020 3003 2037 3006
rect 2236 3003 2261 3006
rect 2276 3003 2285 3006
rect 2290 3003 2308 3006
rect 2324 3003 2333 3006
rect 2370 3003 2380 3006
rect 2396 3003 2413 3006
rect 2418 3003 2436 3006
rect 2530 3003 2572 3006
rect 2706 3003 2788 3006
rect 2812 3003 2837 3006
rect 2844 3003 2853 3006
rect 2922 3003 2956 3006
rect 2980 3003 3013 3006
rect 3018 3005 3021 3013
rect 3052 3003 3093 3006
rect 3386 3005 3389 3013
rect 3570 3003 3580 3006
rect 3634 3003 3668 3006
rect 3850 3005 3853 3013
rect 4026 3005 4029 3013
rect 4050 3013 4060 3016
rect 4212 3013 4237 3016
rect 4258 3013 4268 3016
rect 4362 3013 4412 3016
rect 4442 3013 4460 3016
rect 4474 3013 4524 3016
rect 4626 3013 4676 3016
rect 4706 3013 4732 3016
rect 4050 3003 4053 3013
rect 4106 3003 4124 3006
rect 4162 3003 4188 3006
rect 4204 3003 4229 3006
rect 4284 3003 4293 3006
rect 4322 3003 4332 3006
rect 4348 3003 4397 3006
rect 4468 3003 4485 3006
rect 4498 3003 4516 3006
rect 4554 3003 4596 3006
rect 4612 3003 4661 3006
rect 4740 3003 4773 3006
rect 770 2993 804 2996
rect 922 2993 956 2996
rect 1162 2993 1180 2996
rect 2826 2993 2836 2996
rect 2850 2993 2853 3003
rect 2858 2993 2900 2996
rect 4770 2993 4773 3003
rect 38 2967 4829 2973
rect 2378 2953 2421 2956
rect 3938 2953 3973 2956
rect 866 2943 932 2946
rect 2770 2943 2828 2946
rect 274 2933 284 2936
rect 212 2923 237 2926
rect 306 2925 309 2936
rect 420 2933 469 2936
rect 530 2933 556 2936
rect 572 2933 636 2936
rect 834 2933 844 2936
rect 940 2933 1021 2936
rect 1044 2933 1061 2936
rect 1082 2933 1164 2936
rect 1180 2933 1268 2936
rect 1292 2933 1309 2936
rect 1314 2933 1348 2936
rect 1372 2933 1381 2936
rect 1402 2933 1428 2936
rect 1452 2933 1493 2936
rect 348 2923 373 2926
rect 538 2923 548 2926
rect 748 2923 773 2926
rect 810 2923 852 2926
rect 948 2923 1005 2926
rect 1018 2925 1021 2933
rect 1618 2926 1621 2935
rect 1682 2933 1716 2936
rect 1858 2933 1908 2936
rect 1052 2923 1069 2926
rect 1090 2923 1156 2926
rect 1226 2923 1276 2926
rect 1532 2923 1557 2926
rect 1588 2923 1621 2926
rect 1732 2923 1749 2926
rect 1796 2923 1813 2926
rect 1852 2923 1869 2926
rect 1874 2923 1900 2926
rect 1930 2925 1933 2936
rect 1980 2933 2013 2936
rect 2114 2933 2164 2936
rect 2554 2933 2588 2936
rect 2610 2933 2644 2936
rect 2842 2933 2868 2936
rect 2892 2933 2917 2936
rect 2922 2933 2932 2936
rect 2962 2933 2988 2936
rect 1954 2923 1972 2926
rect 1978 2923 2012 2926
rect 2044 2923 2061 2926
rect 2066 2923 2084 2926
rect 2116 2923 2125 2926
rect 2138 2923 2156 2926
rect 2188 2923 2197 2926
rect 2442 2923 2460 2926
rect 2490 2923 2516 2926
rect 2562 2923 2580 2926
rect 2612 2923 2621 2926
rect 2652 2923 2669 2926
rect 2866 2923 2876 2926
rect 2914 2923 2940 2926
rect 2962 2916 2965 2933
rect 3010 2926 3013 2935
rect 3426 2926 3429 2935
rect 3442 2933 3484 2936
rect 3516 2933 3597 2936
rect 3916 2933 3957 2936
rect 3962 2933 4004 2936
rect 4186 2933 4204 2936
rect 4282 2933 4300 2936
rect 4618 2926 4621 2935
rect 3010 2923 3092 2926
rect 3356 2923 3381 2926
rect 3412 2923 3429 2926
rect 3436 2923 3485 2926
rect 3666 2923 3676 2926
rect 3706 2923 3732 2926
rect 3882 2923 3892 2926
rect 4354 2923 4380 2926
rect 4588 2923 4621 2926
rect 1292 2913 1325 2916
rect 1338 2913 1348 2916
rect 1386 2913 1428 2916
rect 2956 2913 2965 2916
rect 2970 2913 2988 2916
rect 14 2867 4853 2873
rect 3722 2833 3741 2836
rect 4282 2833 4300 2836
rect 740 2823 813 2826
rect 2844 2823 2861 2826
rect 3626 2816 3629 2826
rect 3698 2823 3708 2826
rect 332 2813 357 2816
rect 394 2813 412 2816
rect 468 2813 493 2816
rect 530 2813 548 2816
rect 578 2813 588 2816
rect 706 2813 724 2816
rect 770 2813 820 2816
rect 852 2813 869 2816
rect 906 2813 916 2816
rect 1028 2813 1045 2816
rect 1140 2813 1149 2816
rect 1252 2813 1261 2816
rect 1476 2813 1549 2816
rect 1596 2813 1621 2816
rect 1652 2813 1661 2816
rect 1780 2813 1805 2816
rect 1842 2813 1876 2816
rect 1940 2813 1957 2816
rect 2036 2813 2061 2816
rect 2098 2813 2108 2816
rect 2138 2813 2156 2816
rect 2282 2813 2364 2816
rect 2498 2813 2548 2816
rect 2580 2813 2613 2816
rect 2620 2813 2645 2816
rect 2788 2813 2813 2816
rect 2884 2813 2925 2816
rect 2954 2813 3029 2816
rect 3060 2813 3069 2816
rect 3140 2813 3165 2816
rect 3196 2813 3205 2816
rect 3316 2813 3341 2816
rect 3372 2813 3389 2816
rect 3396 2813 3405 2816
rect 3426 2813 3564 2816
rect 3618 2813 3652 2816
rect 3722 2815 3725 2833
rect 3738 2826 3741 2833
rect 3738 2823 3788 2826
rect 3812 2823 3909 2826
rect 4274 2823 4284 2826
rect 4308 2823 4317 2826
rect 4004 2813 4013 2816
rect 4100 2813 4133 2816
rect 4180 2813 4205 2816
rect 4428 2813 4437 2816
rect 4442 2813 4452 2816
rect 4490 2813 4516 2816
rect 276 2803 293 2806
rect 394 2803 404 2806
rect 556 2803 565 2806
rect 690 2803 716 2806
rect 802 2803 828 2806
rect 844 2803 853 2806
rect 924 2803 965 2806
rect 1020 2803 1101 2806
rect 1498 2803 1501 2813
rect 1682 2803 1700 2806
rect 1732 2803 1741 2806
rect 1884 2803 1901 2806
rect 2122 2803 2164 2806
rect 2180 2803 2372 2806
rect 2388 2803 2405 2806
rect 2418 2803 2460 2806
rect 2538 2803 2556 2806
rect 2578 2803 2612 2806
rect 2786 2803 2820 2806
rect 2876 2803 2885 2806
rect 2890 2803 2932 2806
rect 2954 2805 2957 2813
rect 2988 2803 3013 2806
rect 3018 2803 3036 2806
rect 3068 2803 3077 2806
rect 3202 2805 3205 2813
rect 3218 2803 3244 2806
rect 3386 2805 3389 2813
rect 3618 2806 3621 2813
rect 4546 2806 4549 2814
rect 4588 2813 4621 2816
rect 4780 2813 4805 2816
rect 3498 2803 3572 2806
rect 3588 2803 3621 2806
rect 3660 2803 3669 2806
rect 4082 2803 4092 2806
rect 4434 2803 4444 2806
rect 4482 2803 4524 2806
rect 4546 2803 4557 2806
rect 4580 2803 4669 2806
rect 3018 2796 3021 2803
rect 2746 2793 2772 2796
rect 2850 2793 2868 2796
rect 3002 2793 3021 2796
rect 4434 2783 4437 2803
rect 38 2767 4829 2773
rect 970 2743 996 2746
rect 3258 2743 3301 2746
rect 3258 2736 3261 2743
rect 252 2733 284 2736
rect 322 2733 332 2736
rect 346 2733 380 2736
rect 396 2733 405 2736
rect 538 2733 636 2736
rect 708 2733 765 2736
rect 788 2733 853 2736
rect 986 2733 1004 2736
rect 1034 2733 1061 2736
rect 1084 2733 1148 2736
rect 538 2726 541 2733
rect 1322 2726 1325 2735
rect 1338 2733 1380 2736
rect 1404 2733 1421 2736
rect 1450 2733 1476 2736
rect 1508 2733 1629 2736
rect 1786 2726 1789 2735
rect 1964 2733 2013 2736
rect 2036 2733 2092 2736
rect 2266 2733 2300 2736
rect 2322 2733 2373 2736
rect 2386 2726 2389 2736
rect 2412 2733 2421 2736
rect 2442 2733 2468 2736
rect 2482 2733 2533 2736
rect 2562 2733 2612 2736
rect 2882 2733 2892 2736
rect 2922 2733 2980 2736
rect 3004 2733 3037 2736
rect 3170 2733 3180 2736
rect 3194 2733 3220 2736
rect 3252 2733 3261 2736
rect 3266 2733 3316 2736
rect 100 2723 109 2726
rect 156 2723 181 2726
rect 196 2723 205 2726
rect 218 2723 228 2726
rect 260 2723 285 2726
rect 322 2723 340 2726
rect 524 2723 541 2726
rect 618 2723 644 2726
rect 674 2723 700 2726
rect 754 2723 764 2726
rect 900 2723 909 2726
rect 956 2723 997 2726
rect 1012 2723 1053 2726
rect 1138 2723 1156 2726
rect 1244 2723 1269 2726
rect 1300 2723 1325 2726
rect 1332 2723 1349 2726
rect 1396 2723 1445 2726
rect 1500 2723 1629 2726
rect 1684 2723 1709 2726
rect 1740 2723 1789 2726
rect 1796 2723 1821 2726
rect 1876 2723 1901 2726
rect 1938 2723 1956 2726
rect 2002 2723 2012 2726
rect 2044 2723 2069 2726
rect 2244 2723 2261 2726
rect 2282 2723 2292 2726
rect 2362 2725 2389 2726
rect 2362 2723 2388 2725
rect 2476 2723 2525 2726
rect 2530 2725 2533 2733
rect 2564 2723 2597 2726
rect 2620 2723 2645 2726
rect 2780 2723 2789 2726
rect 2836 2723 2845 2726
rect 2850 2723 2900 2726
rect 2922 2716 2925 2733
rect 3826 2726 3829 2735
rect 3842 2733 3884 2736
rect 3916 2733 3933 2736
rect 4020 2733 4053 2736
rect 3010 2723 3044 2726
rect 3074 2723 3100 2726
rect 3188 2723 3197 2726
rect 3244 2723 3277 2726
rect 3324 2723 3381 2726
rect 3500 2723 3517 2726
rect 3556 2723 3581 2726
rect 3636 2723 3653 2726
rect 3748 2723 3773 2726
rect 3804 2723 3829 2726
rect 3836 2723 3885 2726
rect 1172 2713 1197 2716
rect 2916 2713 2925 2716
rect 2930 2713 2980 2716
rect 3930 2683 3933 2733
rect 4234 2726 4237 2735
rect 4284 2733 4293 2736
rect 4530 2726 4533 2735
rect 4778 2727 4781 2735
rect 3986 2723 4012 2726
rect 4042 2723 4068 2726
rect 4212 2723 4237 2726
rect 4250 2723 4268 2726
rect 4346 2723 4372 2726
rect 4524 2723 4533 2726
rect 4546 2723 4564 2726
rect 4594 2723 4620 2726
rect 4772 2724 4781 2727
rect 4324 2713 4333 2716
rect 14 2667 4853 2673
rect 4250 2633 4284 2636
rect 1244 2623 1269 2626
rect 1282 2623 1300 2626
rect 1330 2623 1380 2626
rect 2852 2623 2885 2626
rect 2930 2623 2964 2626
rect 3500 2623 3525 2626
rect 4242 2623 4268 2626
rect 4292 2623 4309 2626
rect 4364 2623 4405 2626
rect 92 2613 109 2616
rect 124 2613 164 2616
rect 132 2603 157 2606
rect 162 2603 172 2606
rect 194 2603 197 2614
rect 276 2613 301 2616
rect 338 2613 364 2616
rect 428 2613 469 2616
rect 474 2613 484 2616
rect 516 2613 556 2616
rect 754 2613 804 2616
rect 826 2613 852 2616
rect 890 2613 924 2616
rect 956 2613 997 2616
rect 1052 2613 1077 2616
rect 1114 2613 1124 2616
rect 1316 2613 1349 2616
rect 1402 2613 1436 2616
rect 1442 2613 1484 2616
rect 1514 2613 1540 2616
rect 1634 2613 1652 2616
rect 1740 2613 1765 2616
rect 1876 2613 1893 2616
rect 1930 2613 1956 2616
rect 2252 2613 2277 2616
rect 2316 2613 2325 2616
rect 2442 2613 2500 2616
rect 2530 2613 2556 2616
rect 2594 2613 2620 2616
rect 2626 2613 2668 2616
rect 2772 2613 2821 2616
rect 2826 2613 2836 2616
rect 2890 2613 2901 2616
rect 2908 2613 2965 2616
rect 2980 2613 2989 2616
rect 3034 2613 3076 2616
rect 3114 2613 3132 2616
rect 3236 2613 3261 2616
rect 3316 2613 3341 2616
rect 3346 2613 3356 2616
rect 436 2603 485 2606
rect 508 2603 541 2606
rect 580 2603 613 2606
rect 732 2603 789 2606
rect 850 2603 860 2606
rect 882 2603 932 2606
rect 1164 2603 1173 2606
rect 1178 2603 1220 2606
rect 1244 2603 1261 2606
rect 1282 2603 1300 2606
rect 1330 2603 1380 2606
rect 1402 2605 1405 2613
rect 1442 2605 1445 2613
rect 1578 2603 1604 2606
rect 1660 2603 1677 2606
rect 1682 2603 1724 2606
rect 2330 2603 2412 2606
rect 2594 2603 2612 2606
rect 2666 2603 2676 2606
rect 2692 2603 2749 2606
rect 2770 2603 2828 2606
rect 2852 2603 2893 2606
rect 2898 2605 2901 2613
rect 3410 2606 3413 2614
rect 3562 2613 3660 2616
rect 2922 2603 2964 2606
rect 3036 2603 3061 2606
rect 3322 2603 3348 2606
rect 3362 2603 3381 2606
rect 3410 2603 3453 2606
rect 3564 2603 3573 2606
rect 3578 2603 3652 2606
rect 3770 2605 3773 2616
rect 3778 2613 3852 2616
rect 3884 2613 3956 2616
rect 4010 2613 4060 2616
rect 4090 2613 4124 2616
rect 4130 2613 4148 2616
rect 4178 2613 4204 2616
rect 4324 2613 4333 2616
rect 4410 2613 4420 2616
rect 4548 2613 4573 2616
rect 4604 2613 4613 2616
rect 4658 2613 4676 2616
rect 4706 2613 4732 2616
rect 3834 2603 3860 2606
rect 3876 2603 3885 2606
rect 3980 2603 3997 2606
rect 4026 2603 4052 2606
rect 4130 2605 4133 2613
rect 4306 2603 4316 2606
rect 4370 2603 4412 2606
rect 4444 2603 4453 2606
rect 4484 2603 4493 2606
rect 4650 2603 4668 2606
rect 4740 2603 4789 2606
rect 594 2593 724 2596
rect 1130 2593 1156 2596
rect 2706 2593 2756 2596
rect 3690 2583 3733 2586
rect 38 2567 4829 2573
rect 330 2536 333 2546
rect 946 2543 1004 2546
rect 2866 2543 2900 2546
rect 4434 2536 4437 2546
rect 330 2533 364 2536
rect 380 2533 397 2536
rect 570 2533 596 2536
rect 610 2533 644 2536
rect 740 2533 805 2536
rect 890 2533 916 2536
rect 938 2533 1012 2536
rect 1034 2533 1077 2536
rect 1100 2533 1109 2536
rect 1204 2533 1221 2536
rect 1258 2533 1276 2536
rect 1300 2533 1317 2536
rect 1322 2533 1348 2536
rect 308 2523 333 2526
rect 346 2523 356 2526
rect 388 2523 405 2526
rect 570 2523 604 2526
rect 618 2523 652 2526
rect 714 2523 732 2526
rect 754 2523 804 2526
rect 938 2525 941 2533
rect 1020 2523 1069 2526
rect 1074 2525 1077 2533
rect 1108 2523 1133 2526
rect 1170 2523 1180 2526
rect 1218 2506 1221 2533
rect 1226 2523 1284 2526
rect 1322 2523 1325 2533
rect 1362 2526 1365 2535
rect 1586 2533 1612 2536
rect 1626 2526 1629 2536
rect 1778 2533 1796 2536
rect 1898 2533 1980 2536
rect 1996 2533 2101 2536
rect 2130 2533 2140 2536
rect 2154 2533 2196 2536
rect 2258 2533 2316 2536
rect 2338 2535 2420 2536
rect 2338 2533 2421 2535
rect 2452 2533 2461 2536
rect 2570 2533 2620 2536
rect 2794 2533 2836 2536
rect 2922 2533 2956 2536
rect 2980 2533 2997 2536
rect 3194 2533 3204 2536
rect 3284 2533 3317 2536
rect 1356 2523 1365 2526
rect 1372 2523 1389 2526
rect 1402 2523 1444 2526
rect 1482 2523 1492 2526
rect 1602 2523 1629 2526
rect 1674 2523 1684 2526
rect 1714 2523 1740 2526
rect 1834 2523 1868 2526
rect 1900 2523 1965 2526
rect 2004 2523 2148 2526
rect 2212 2523 2221 2526
rect 2252 2523 2293 2526
rect 2340 2523 2389 2526
rect 2418 2523 2421 2533
rect 2530 2523 2540 2526
rect 2572 2523 2621 2526
rect 2628 2523 2661 2526
rect 2772 2523 2789 2526
rect 2826 2523 2844 2526
rect 2972 2523 2997 2526
rect 3036 2523 3045 2526
rect 3146 2523 3164 2526
rect 3220 2523 3268 2526
rect 3394 2525 3397 2536
rect 3452 2533 3469 2536
rect 3514 2533 3540 2536
rect 3572 2533 3581 2536
rect 3618 2533 3660 2536
rect 1300 2513 1309 2516
rect 1380 2513 1437 2516
rect 2860 2513 2893 2516
rect 3306 2513 3332 2516
rect 3346 2506 3349 2525
rect 3418 2523 3436 2526
rect 3362 2513 3380 2516
rect 3458 2513 3484 2516
rect 3578 2513 3581 2533
rect 3866 2526 3869 2535
rect 3908 2533 3941 2536
rect 4042 2533 4116 2536
rect 4306 2533 4324 2536
rect 4362 2533 4396 2536
rect 4412 2533 4437 2536
rect 4466 2533 4556 2536
rect 4588 2533 4605 2536
rect 4642 2533 4652 2536
rect 3586 2523 3612 2526
rect 3668 2523 3677 2526
rect 3690 2523 3700 2526
rect 3780 2523 3789 2526
rect 3836 2523 3869 2526
rect 3938 2526 3941 2533
rect 4434 2526 4437 2533
rect 3938 2523 3972 2526
rect 4220 2523 4245 2526
rect 4282 2523 4292 2526
rect 4378 2523 4388 2526
rect 4434 2523 4452 2526
rect 4546 2523 4564 2526
rect 4636 2523 4660 2526
rect 3362 2506 3365 2513
rect 1218 2503 1269 2506
rect 3346 2503 3365 2506
rect 14 2467 4853 2473
rect 3322 2433 3341 2436
rect 836 2423 1125 2426
rect 1282 2423 1300 2426
rect 2842 2423 2877 2426
rect 2916 2423 2925 2426
rect 2954 2423 2980 2426
rect 3298 2423 3308 2426
rect 2874 2416 2877 2423
rect 196 2413 228 2416
rect 388 2413 413 2416
rect 450 2413 468 2416
rect 474 2413 500 2416
rect 532 2413 565 2416
rect 618 2413 644 2416
rect 708 2413 717 2416
rect 770 2413 820 2416
rect 1148 2413 1165 2416
rect 1204 2413 1213 2416
rect 1316 2413 1325 2416
rect 1410 2413 1525 2416
rect 1556 2413 1605 2416
rect 1652 2413 1669 2416
rect 1708 2413 1733 2416
rect 1786 2413 1796 2416
rect 1908 2413 2076 2416
rect 2250 2413 2260 2416
rect 2292 2413 2325 2416
rect 2364 2413 2405 2416
rect 2442 2413 2468 2416
rect 2506 2413 2556 2416
rect 2660 2413 2685 2416
rect 2780 2413 2789 2416
rect 2828 2413 2869 2416
rect 2874 2413 2900 2416
rect 132 2403 141 2406
rect 162 2403 172 2406
rect 188 2403 213 2406
rect 252 2403 285 2406
rect 476 2403 485 2406
rect 498 2403 508 2406
rect 524 2403 549 2406
rect 604 2403 613 2406
rect 626 2403 636 2406
rect 770 2403 812 2406
rect 836 2403 845 2406
rect 1274 2403 1300 2406
rect 1324 2403 1381 2406
rect 1410 2405 1413 2413
rect 1476 2403 1485 2406
rect 1564 2403 1589 2406
rect 1730 2405 1733 2413
rect 2922 2406 2925 2423
rect 3042 2413 3060 2416
rect 3106 2413 3132 2416
rect 3242 2413 3252 2416
rect 3322 2415 3325 2433
rect 3338 2426 3341 2433
rect 3338 2423 3372 2426
rect 3396 2423 3429 2426
rect 4322 2423 4332 2426
rect 4356 2423 4365 2426
rect 1812 2403 1821 2406
rect 1916 2403 1933 2406
rect 2058 2403 2068 2406
rect 2242 2403 2268 2406
rect 2284 2403 2325 2406
rect 2330 2403 2356 2406
rect 2546 2403 2564 2406
rect 2580 2403 2629 2406
rect 2642 2403 2652 2406
rect 2826 2403 2892 2406
rect 2922 2403 2980 2406
rect 3004 2403 3013 2406
rect 3084 2403 3125 2406
rect 3212 2403 3229 2406
rect 3442 2403 3445 2414
rect 3476 2413 3501 2416
rect 3548 2413 3557 2416
rect 3618 2413 3636 2416
rect 3716 2413 3725 2416
rect 3772 2413 3813 2416
rect 3850 2413 3860 2416
rect 3978 2413 3988 2416
rect 4034 2413 4044 2416
rect 4122 2413 4140 2416
rect 4170 2413 4196 2416
rect 4274 2413 4292 2416
rect 4404 2413 4429 2416
rect 4500 2413 4525 2416
rect 4556 2413 4573 2416
rect 3468 2403 3509 2406
rect 3618 2403 3621 2413
rect 3660 2403 3677 2406
rect 3810 2405 3813 2413
rect 3876 2403 3925 2406
rect 3972 2403 3981 2406
rect 4122 2405 4125 2413
rect 4274 2403 4284 2406
rect 4570 2405 4573 2413
rect 4586 2406 4589 2416
rect 4642 2413 4668 2416
rect 4642 2406 4645 2413
rect 4586 2403 4604 2406
rect 4620 2403 4645 2406
rect 2322 2396 2325 2403
rect 538 2393 596 2396
rect 2322 2393 2341 2396
rect 2786 2393 2812 2396
rect 38 2367 4829 2373
rect 3226 2353 3349 2356
rect 634 2343 644 2346
rect 2866 2343 2908 2346
rect 2922 2343 2965 2346
rect 2922 2336 2925 2343
rect 180 2333 189 2336
rect 252 2333 316 2336
rect 362 2333 380 2336
rect 402 2333 436 2336
rect 578 2333 612 2336
rect 652 2333 669 2336
rect 578 2326 581 2333
rect 826 2326 829 2335
rect 874 2333 924 2336
rect 946 2333 957 2336
rect 108 2323 125 2326
rect 178 2323 188 2326
rect 220 2323 228 2326
rect 362 2323 372 2326
rect 404 2323 413 2326
rect 564 2323 581 2326
rect 628 2323 637 2326
rect 660 2323 677 2326
rect 772 2323 829 2326
rect 866 2323 916 2326
rect 946 2325 949 2333
rect 986 2316 989 2336
rect 1138 2333 1148 2336
rect 1068 2323 1085 2326
rect 1130 2323 1140 2326
rect 1170 2325 1173 2336
rect 1220 2333 1229 2336
rect 1234 2333 1300 2336
rect 1324 2333 1365 2336
rect 1564 2333 1581 2336
rect 1884 2333 1933 2336
rect 1178 2323 1212 2326
rect 1316 2323 1325 2326
rect 1412 2323 1437 2326
rect 1468 2323 1493 2326
rect 1556 2323 1660 2326
rect 1772 2323 1789 2326
rect 1834 2323 1876 2326
rect 1962 2325 1965 2336
rect 2100 2333 2165 2336
rect 2188 2333 2245 2336
rect 2306 2333 2348 2336
rect 2364 2333 2413 2336
rect 2410 2326 2413 2333
rect 2578 2333 2652 2336
rect 2786 2333 2836 2336
rect 2860 2333 2909 2336
rect 2916 2333 2925 2336
rect 2930 2333 2980 2336
rect 3004 2333 3021 2336
rect 2004 2323 2029 2326
rect 2066 2323 2092 2326
rect 2218 2323 2276 2326
rect 2330 2323 2340 2326
rect 2372 2323 2397 2326
rect 2410 2323 2436 2326
rect 2474 2323 2492 2326
rect 2578 2323 2581 2333
rect 2786 2326 2789 2333
rect 3170 2326 3173 2335
rect 3186 2333 3204 2336
rect 3420 2333 3429 2336
rect 3442 2333 3476 2336
rect 3492 2333 3525 2336
rect 3626 2333 3644 2336
rect 3802 2326 3805 2335
rect 3938 2333 3948 2336
rect 3986 2333 4004 2336
rect 4036 2333 4061 2336
rect 4338 2333 4380 2336
rect 4396 2333 4413 2336
rect 4554 2326 4557 2335
rect 4628 2333 4637 2336
rect 4754 2326 4757 2335
rect 2660 2323 2685 2326
rect 2780 2323 2789 2326
rect 3084 2323 3093 2326
rect 3140 2323 3173 2326
rect 3180 2323 3189 2326
rect 3220 2323 3285 2326
rect 3412 2323 3461 2326
rect 3564 2323 3573 2326
rect 3642 2323 3652 2326
rect 3796 2323 3805 2326
rect 3868 2323 3893 2326
rect 3946 2323 3956 2326
rect 4114 2323 4140 2326
rect 4220 2323 4245 2326
rect 4354 2323 4372 2326
rect 4418 2323 4428 2326
rect 4548 2323 4557 2326
rect 4570 2323 4604 2326
rect 4748 2323 4757 2326
rect 852 2313 909 2316
rect 954 2313 989 2316
rect 1282 2313 1300 2316
rect 2266 2313 2269 2323
rect 2860 2313 2893 2316
rect 2930 2313 2980 2316
rect 4282 2313 4300 2316
rect 4324 2313 4365 2316
rect 4282 2303 4316 2306
rect 14 2267 4853 2273
rect 3330 2233 3421 2236
rect 4242 2233 4261 2236
rect 4300 2233 4309 2236
rect 1282 2223 1300 2226
rect 1362 2223 1420 2226
rect 2820 2223 2869 2226
rect 2914 2223 2924 2226
rect 3306 2223 3316 2226
rect 108 2213 133 2216
rect 188 2213 205 2216
rect 322 2213 364 2216
rect 370 2213 388 2216
rect 426 2213 460 2216
rect 594 2213 620 2216
rect 700 2213 717 2216
rect 858 2213 884 2216
rect 978 2213 988 2216
rect 1026 2213 1180 2216
rect 1212 2213 1285 2216
rect 1316 2213 1325 2216
rect 1516 2213 1541 2216
rect 1596 2213 1605 2216
rect 1738 2213 1748 2216
rect 1778 2213 1804 2216
rect 1842 2213 1876 2216
rect 1930 2213 1940 2216
rect 1972 2213 1989 2216
rect 2028 2213 2053 2216
rect 2090 2213 2100 2216
rect 2106 2213 2172 2216
rect 2284 2213 2309 2216
rect 2322 2213 2332 2216
rect 2364 2213 2381 2216
rect 2436 2213 2477 2216
rect 2490 2213 2564 2216
rect 2732 2213 2797 2216
rect 2876 2213 2925 2216
rect 2940 2213 2949 2216
rect 3034 2213 3060 2216
rect 3186 2213 3228 2216
rect 3258 2213 3268 2216
rect 3330 2215 3333 2233
rect 3340 2223 3421 2226
rect 3346 2213 3389 2216
rect 3394 2213 3428 2216
rect 3474 2213 3484 2216
rect 3522 2213 3556 2216
rect 3788 2213 3797 2216
rect 3900 2213 3932 2216
rect 3970 2213 3988 2216
rect 3994 2213 4005 2216
rect 4042 2213 4068 2216
rect 4074 2213 4084 2216
rect 4114 2213 4140 2216
rect 4242 2215 4245 2233
rect 4258 2226 4261 2233
rect 4258 2223 4292 2226
rect 4316 2223 4325 2226
rect 4364 2213 4381 2216
rect 4386 2213 4405 2216
rect 4556 2213 4565 2216
rect 4620 2213 4637 2216
rect 4698 2213 4756 2216
rect 426 2206 429 2213
rect 372 2203 389 2206
rect 418 2203 429 2206
rect 450 2203 468 2206
rect 490 2203 548 2206
rect 804 2203 813 2206
rect 834 2203 892 2206
rect 938 2203 996 2206
rect 1012 2203 1053 2206
rect 1122 2203 1188 2206
rect 1210 2203 1300 2206
rect 1324 2203 1405 2206
rect 1444 2203 1485 2206
rect 1490 2203 1508 2206
rect 1530 2203 1572 2206
rect 1604 2203 1653 2206
rect 1700 2203 1733 2206
rect 1884 2203 1941 2206
rect 2108 2203 2173 2206
rect 2196 2203 2213 2206
rect 2290 2203 2340 2206
rect 2356 2203 2365 2206
rect 2386 2203 2428 2206
rect 2588 2203 2629 2206
rect 2794 2205 2797 2213
rect 2820 2203 2829 2206
rect 2890 2203 2924 2206
rect 2948 2203 3045 2206
rect 3084 2203 3156 2206
rect 3210 2203 3220 2206
rect 3436 2203 3469 2206
rect 3508 2203 3541 2206
rect 3596 2203 3621 2206
rect 3626 2203 3636 2206
rect 3668 2203 3685 2206
rect 3794 2205 3797 2213
rect 3970 2206 3973 2213
rect 3810 2203 3820 2206
rect 3858 2203 3876 2206
rect 3892 2203 3925 2206
rect 3956 2203 3973 2206
rect 4002 2205 4005 2213
rect 4036 2203 4061 2206
rect 4074 2205 4077 2213
rect 4330 2203 4340 2206
rect 4356 2203 4397 2206
rect 4402 2205 4405 2213
rect 4436 2203 4453 2206
rect 4562 2205 4565 2213
rect 4650 2203 4660 2206
rect 4692 2203 4709 2206
rect 4764 2203 4789 2206
rect 3810 2183 3813 2203
rect 38 2167 4829 2173
rect 2666 2143 2756 2146
rect 2770 2143 2844 2146
rect 116 2133 229 2136
rect 410 2134 420 2136
rect 242 2126 245 2134
rect 410 2133 421 2134
rect 458 2133 524 2136
rect 556 2133 573 2136
rect 604 2133 613 2136
rect 618 2133 644 2136
rect 810 2133 836 2136
rect 866 2133 916 2136
rect 946 2133 980 2136
rect 1004 2133 1013 2136
rect 1034 2133 1076 2136
rect 1100 2133 1125 2136
rect 1282 2133 1388 2136
rect 1412 2133 1437 2136
rect 1516 2133 1533 2136
rect 418 2126 421 2133
rect 1666 2126 1669 2134
rect 2034 2133 2044 2136
rect 2076 2133 2085 2136
rect 2196 2133 2253 2136
rect 2578 2133 2629 2136
rect 2652 2133 2733 2136
rect 2764 2133 2845 2136
rect 2852 2133 2893 2136
rect 3004 2133 3021 2136
rect 3252 2133 3261 2136
rect 3474 2133 3500 2136
rect 3532 2133 3573 2136
rect 3618 2133 3652 2136
rect 3690 2133 3716 2136
rect 194 2123 236 2126
rect 242 2123 269 2126
rect 316 2123 325 2126
rect 372 2123 421 2126
rect 554 2123 580 2126
rect 660 2123 669 2126
rect 674 2123 708 2126
rect 786 2123 828 2126
rect 1178 2123 1252 2126
rect 1284 2123 1301 2126
rect 1306 2123 1396 2126
rect 1580 2123 1589 2126
rect 1636 2123 1669 2126
rect 1682 2123 1700 2126
rect 1788 2123 1813 2126
rect 1844 2123 1901 2126
rect 2068 2123 2172 2126
rect 2386 2123 2420 2126
rect 2458 2123 2492 2126
rect 2572 2123 2621 2126
rect 2626 2125 2629 2133
rect 3906 2126 3909 2134
rect 3922 2133 3956 2136
rect 4004 2133 4029 2136
rect 4242 2126 4245 2134
rect 4258 2133 4356 2136
rect 4394 2133 4444 2136
rect 4474 2133 4492 2136
rect 4522 2133 4532 2136
rect 2772 2123 2829 2126
rect 2924 2123 2957 2126
rect 2996 2123 3005 2126
rect 3010 2123 3028 2126
rect 3058 2123 3084 2126
rect 3156 2123 3173 2126
rect 3218 2123 3236 2126
rect 666 2116 669 2123
rect 1298 2116 1301 2123
rect 666 2113 677 2116
rect 1004 2113 1061 2116
rect 1066 2113 1076 2116
rect 1298 2113 1373 2116
rect 1412 2113 1421 2116
rect 3258 2113 3268 2116
rect 3282 2106 3285 2125
rect 3474 2123 3508 2126
rect 3604 2123 3660 2126
rect 3740 2123 3805 2126
rect 3900 2123 3909 2126
rect 3930 2123 3964 2126
rect 4010 2123 4044 2126
rect 4236 2123 4245 2126
rect 4452 2123 4461 2126
rect 4468 2123 4485 2126
rect 4516 2123 4525 2126
rect 4612 2123 4637 2126
rect 4780 2123 4789 2126
rect 3298 2113 3332 2116
rect 3356 2113 3373 2116
rect 3298 2106 3301 2113
rect 3282 2103 3301 2106
rect 14 2067 4853 2073
rect 1858 2033 1925 2036
rect 202 2003 220 2006
rect 242 2003 260 2006
rect 282 2003 285 2014
rect 306 2013 316 2016
rect 348 2014 365 2016
rect 346 2013 365 2014
rect 484 2013 525 2016
rect 578 2013 596 2016
rect 700 2013 717 2016
rect 972 2013 997 2016
rect 1020 2013 1037 2016
rect 1050 2013 1076 2016
rect 1164 2013 1261 2016
rect 1284 2013 1365 2016
rect 1548 2013 1565 2016
rect 1628 2013 1677 2016
rect 1706 2013 1732 2016
rect 1804 2013 1829 2016
rect 346 2006 349 2013
rect 1858 2006 1861 2033
rect 2836 2023 2901 2026
rect 3258 2023 3276 2026
rect 3450 2023 3492 2026
rect 3516 2023 3661 2026
rect 2898 2016 2901 2023
rect 308 2003 317 2006
rect 346 2003 357 2006
rect 378 2003 468 2006
rect 514 2003 532 2006
rect 564 2003 573 2006
rect 666 2003 676 2006
rect 692 2003 709 2006
rect 1092 2003 1133 2006
rect 1138 2003 1156 2006
rect 1266 2003 1276 2006
rect 1330 2003 1532 2006
rect 1602 2003 1612 2006
rect 1852 2003 1861 2006
rect 1954 2013 2028 2016
rect 2060 2014 2149 2016
rect 2058 2013 2149 2014
rect 2188 2013 2213 2016
rect 2244 2013 2253 2016
rect 2330 2013 2340 2016
rect 2372 2013 2381 2016
rect 2476 2013 2485 2016
rect 2748 2013 2813 2016
rect 2898 2013 2909 2016
rect 2924 2013 2949 2016
rect 2988 2013 3005 2016
rect 3106 2013 3132 2016
rect 3212 2013 3269 2016
rect 3364 2013 3405 2016
rect 3436 2013 3477 2016
rect 3684 2013 3709 2016
rect 1954 2003 1957 2013
rect 2018 2003 2036 2006
rect 2058 2003 2061 2013
rect 2250 2006 2253 2013
rect 2250 2003 2348 2006
rect 2554 2003 2596 2006
rect 2612 2003 2653 2006
rect 2810 2005 2813 2013
rect 2836 2003 2861 2006
rect 2906 2005 2909 2013
rect 3002 2006 3005 2013
rect 3810 2006 3813 2026
rect 3844 2013 3877 2016
rect 2932 2003 2941 2006
rect 2954 2003 2964 2006
rect 3002 2003 3012 2006
rect 3044 2003 3069 2006
rect 3170 2003 3196 2006
rect 3330 2003 3340 2006
rect 3370 2003 3412 2006
rect 3538 2003 3660 2006
rect 3810 2003 3820 2006
rect 3898 2003 3901 2014
rect 4050 2013 4060 2016
rect 4090 2013 4108 2016
rect 4114 2013 4132 2016
rect 4162 2013 4188 2016
rect 4260 2013 4285 2016
rect 4316 2013 4325 2016
rect 4476 2013 4493 2016
rect 4532 2013 4573 2016
rect 4594 2013 4604 2016
rect 4618 2013 4644 2016
rect 3924 2003 3949 2006
rect 4114 2005 4117 2013
rect 4322 2005 4325 2013
rect 4370 2003 4452 2006
rect 4570 2003 4573 2013
rect 4612 2003 4629 2006
rect 354 1993 357 2003
rect 858 1993 956 1996
rect 978 1993 1004 1996
rect 1098 1993 1148 1996
rect 38 1967 4829 1973
rect 594 1943 652 1946
rect 2930 1943 2980 1946
rect 4338 1936 4341 1946
rect 66 1933 84 1936
rect 106 1933 116 1936
rect 106 1926 109 1933
rect 100 1923 109 1926
rect 132 1923 141 1926
rect 180 1923 197 1926
rect 250 1923 253 1934
rect 466 1933 484 1936
rect 522 1933 540 1936
rect 588 1933 621 1936
rect 660 1933 669 1936
rect 740 1933 789 1936
rect 804 1933 829 1936
rect 1044 1933 1053 1936
rect 1122 1933 1164 1936
rect 1180 1933 1213 1936
rect 1490 1933 1548 1936
rect 1578 1933 1604 1936
rect 1644 1933 1677 1936
rect 1748 1933 1765 1936
rect 1810 1933 1828 1936
rect 1914 1933 1964 1936
rect 1980 1933 2013 1936
rect 2332 1933 2357 1936
rect 2410 1933 2452 1936
rect 2738 1933 2788 1936
rect 2812 1933 2821 1936
rect 1762 1926 1765 1933
rect 2898 1926 2901 1934
rect 2924 1933 2973 1936
rect 2988 1933 3013 1936
rect 3036 1933 3045 1936
rect 3068 1933 3077 1936
rect 3260 1933 3269 1936
rect 3324 1933 3365 1936
rect 3370 1933 3380 1936
rect 3362 1926 3365 1933
rect 3418 1926 3421 1936
rect 3516 1933 3533 1936
rect 3748 1933 3781 1936
rect 3804 1933 3829 1936
rect 4316 1933 4341 1936
rect 3530 1926 3533 1933
rect 292 1923 301 1926
rect 508 1923 533 1926
rect 668 1923 693 1926
rect 716 1923 725 1926
rect 732 1923 741 1926
rect 852 1923 861 1926
rect 962 1923 1020 1926
rect 1052 1923 1085 1926
rect 1138 1923 1156 1926
rect 1188 1923 1245 1926
rect 1356 1923 1365 1926
rect 1412 1923 1421 1926
rect 1434 1923 1460 1926
rect 1506 1923 1556 1926
rect 1620 1923 1628 1926
rect 1700 1923 1725 1926
rect 1762 1923 1788 1926
rect 1908 1923 1949 1926
rect 2050 1923 2076 1926
rect 2266 1923 2324 1926
rect 2404 1923 2445 1926
rect 2482 1923 2548 1926
rect 2580 1923 2621 1926
rect 2634 1923 2708 1926
rect 2890 1923 2901 1926
rect 3002 1923 3020 1926
rect 3050 1923 3060 1926
rect 3274 1923 3300 1926
rect 3362 1923 3421 1926
rect 3482 1923 3492 1926
rect 3530 1923 3588 1926
rect 3610 1923 3620 1926
rect 3650 1923 3676 1926
rect 3714 1923 3740 1926
rect 3746 1923 3780 1926
rect 3938 1923 3948 1926
rect 3978 1923 4004 1926
rect 4100 1923 4125 1926
rect 4228 1923 4237 1926
rect 4412 1923 4437 1926
rect 4666 1923 4692 1926
rect 2890 1916 2893 1923
rect 2812 1913 2893 1916
rect 3074 1913 3124 1916
rect 3154 1913 3188 1916
rect 3154 1906 3157 1913
rect 3138 1903 3157 1906
rect 14 1867 4853 1873
rect 2738 1823 2804 1826
rect 2874 1823 2909 1826
rect 2924 1823 2933 1826
rect 3002 1823 3012 1826
rect 3074 1823 3124 1826
rect 2874 1816 2877 1823
rect 3002 1816 3005 1823
rect 180 1813 205 1816
rect 276 1814 316 1816
rect 274 1813 316 1814
rect 242 1803 251 1806
rect 274 1803 277 1813
rect 346 1806 349 1814
rect 476 1813 493 1816
rect 532 1813 597 1816
rect 602 1813 628 1816
rect 666 1813 708 1816
rect 738 1813 748 1816
rect 842 1813 892 1816
rect 954 1813 972 1816
rect 1004 1813 1013 1816
rect 1076 1813 1133 1816
rect 1140 1813 1149 1816
rect 1252 1813 1261 1816
rect 1332 1813 1341 1816
rect 1346 1813 1404 1816
rect 1660 1813 1701 1816
rect 1738 1813 1788 1816
rect 1898 1813 1908 1816
rect 1956 1813 1965 1816
rect 1978 1813 2036 1816
rect 2066 1813 2108 1816
rect 2146 1813 2172 1816
rect 2202 1813 2277 1816
rect 602 1806 605 1813
rect 738 1806 741 1813
rect 1698 1806 1701 1813
rect 298 1803 324 1806
rect 346 1803 373 1806
rect 378 1803 396 1806
rect 412 1803 437 1806
rect 570 1803 605 1806
rect 666 1803 700 1806
rect 732 1803 741 1806
rect 908 1803 957 1806
rect 962 1803 980 1806
rect 996 1803 1013 1806
rect 1026 1803 1068 1806
rect 1090 1803 1132 1806
rect 1258 1803 1308 1806
rect 1340 1803 1397 1806
rect 1428 1803 1445 1806
rect 1698 1803 1708 1806
rect 1740 1803 1781 1806
rect 2060 1803 2069 1806
rect 2282 1803 2285 1814
rect 2372 1813 2381 1816
rect 2412 1813 2429 1816
rect 2484 1813 2525 1816
rect 2540 1813 2573 1816
rect 2610 1813 2636 1816
rect 2732 1813 2805 1816
rect 2812 1813 2861 1816
rect 2868 1813 2877 1816
rect 2882 1813 2980 1816
rect 2994 1813 3005 1816
rect 3028 1813 3052 1816
rect 3178 1813 3196 1816
rect 3218 1813 3244 1816
rect 3300 1813 3333 1816
rect 3524 1813 3533 1816
rect 3586 1813 3604 1816
rect 3652 1813 3717 1816
rect 3724 1813 3764 1816
rect 3826 1813 3852 1816
rect 3932 1813 3972 1816
rect 4130 1813 4164 1816
rect 4258 1813 4276 1816
rect 4404 1813 4413 1816
rect 4452 1813 4477 1816
rect 4516 1813 4525 1816
rect 4562 1813 4588 1816
rect 4708 1813 4717 1816
rect 2378 1803 2388 1806
rect 2418 1803 2460 1806
rect 2820 1803 2860 1806
rect 2874 1803 2908 1806
rect 2922 1803 2972 1806
rect 2994 1805 2997 1813
rect 3002 1803 3012 1806
rect 3076 1803 3109 1806
rect 3260 1803 3269 1806
rect 3274 1803 3292 1806
rect 3626 1803 3644 1806
rect 3732 1803 3749 1806
rect 3900 1803 3925 1806
rect 3946 1803 3964 1806
rect 4138 1803 4156 1806
rect 4194 1803 4220 1806
rect 4252 1803 4269 1806
rect 4466 1803 4492 1806
rect 4626 1803 4636 1806
rect 4780 1803 4789 1806
rect 1018 1793 1060 1796
rect 38 1767 4829 1773
rect 890 1743 940 1746
rect 2202 1743 2244 1746
rect 178 1733 220 1736
rect 236 1733 245 1736
rect 372 1733 389 1736
rect 412 1733 452 1736
rect 540 1733 557 1736
rect 588 1733 597 1736
rect 610 1733 636 1736
rect 668 1733 693 1736
rect 804 1733 853 1736
rect 948 1733 965 1736
rect 1100 1733 1197 1736
rect 1316 1733 1325 1736
rect 1402 1733 1460 1736
rect 1556 1733 1589 1736
rect 1660 1733 1717 1736
rect 1740 1733 1757 1736
rect 1834 1733 1884 1736
rect 1754 1726 1757 1733
rect 116 1723 133 1726
rect 172 1723 205 1726
rect 300 1723 325 1726
rect 370 1723 388 1726
rect 426 1723 460 1726
rect 490 1723 532 1726
rect 538 1723 564 1726
rect 596 1723 621 1726
rect 626 1723 644 1726
rect 732 1723 741 1726
rect 796 1723 805 1726
rect 842 1723 852 1726
rect 884 1723 893 1726
rect 956 1723 1069 1726
rect 1186 1723 1204 1726
rect 1242 1723 1292 1726
rect 1322 1723 1372 1726
rect 1402 1723 1452 1726
rect 1484 1723 1532 1726
rect 1602 1723 1652 1726
rect 1698 1723 1716 1726
rect 1754 1723 1796 1726
rect 1906 1725 1909 1736
rect 2196 1733 2245 1736
rect 2258 1733 2276 1736
rect 2324 1733 2365 1736
rect 2436 1733 2445 1736
rect 2450 1726 2453 1733
rect 2466 1726 2469 1744
rect 2938 1743 2948 1746
rect 2610 1733 2628 1736
rect 2804 1733 2813 1736
rect 2916 1733 2933 1736
rect 3004 1733 3021 1736
rect 3042 1726 3045 1744
rect 3052 1733 3069 1736
rect 3410 1733 3420 1736
rect 3434 1733 3460 1736
rect 3492 1733 3501 1736
rect 3572 1733 3589 1736
rect 3772 1733 3789 1736
rect 3988 1733 4005 1736
rect 3706 1726 3709 1733
rect 3938 1726 3941 1733
rect 4002 1726 4005 1733
rect 4034 1733 4044 1736
rect 4100 1733 4125 1736
rect 4364 1733 4397 1736
rect 4426 1733 4444 1736
rect 4588 1733 4597 1736
rect 4602 1733 4644 1736
rect 4682 1733 4700 1736
rect 4034 1726 4037 1733
rect 1962 1723 1972 1726
rect 2010 1723 2044 1726
rect 2074 1723 2116 1726
rect 2154 1723 2172 1726
rect 2290 1723 2357 1726
rect 2402 1723 2412 1726
rect 2442 1723 2453 1726
rect 2460 1723 2469 1726
rect 2554 1723 2572 1726
rect 2618 1723 2636 1726
rect 2796 1723 2805 1726
rect 2842 1723 2884 1726
rect 2970 1723 3045 1726
rect 3434 1723 3468 1726
rect 3498 1723 3508 1726
rect 3514 1723 3556 1726
rect 3628 1723 3653 1726
rect 3684 1723 3709 1726
rect 3716 1723 3748 1726
rect 3778 1723 3804 1726
rect 3844 1723 3869 1726
rect 3900 1723 3941 1726
rect 3948 1723 3964 1726
rect 4002 1723 4037 1726
rect 4068 1723 4092 1726
rect 4330 1723 4340 1726
rect 4370 1723 4404 1726
rect 4442 1723 4452 1726
rect 4482 1723 4524 1726
rect 4586 1723 4652 1726
rect 4730 1723 4756 1726
rect 842 1703 845 1723
rect 2442 1716 2445 1723
rect 2554 1716 2557 1723
rect 2618 1716 2621 1723
rect 2434 1713 2445 1716
rect 2490 1713 2524 1716
rect 2548 1713 2557 1716
rect 2604 1713 2621 1716
rect 2674 1713 2716 1716
rect 3098 1713 3116 1716
rect 3146 1713 3172 1716
rect 3196 1713 3205 1716
rect 3210 1713 3236 1716
rect 3260 1713 3285 1716
rect 3722 1713 3725 1723
rect 1818 1703 1853 1706
rect 2650 1703 2660 1706
rect 2674 1703 2732 1706
rect 3090 1703 3132 1706
rect 3146 1703 3149 1713
rect 3170 1703 3188 1706
rect 3210 1703 3252 1706
rect 14 1667 4853 1673
rect 1218 1643 1245 1646
rect 2796 1633 2845 1636
rect 2954 1633 2964 1636
rect 3122 1633 3172 1636
rect 3218 1633 3260 1636
rect 4562 1633 4581 1636
rect 2812 1623 2829 1626
rect 2922 1623 2948 1626
rect 2972 1623 2997 1626
rect 3050 1623 3068 1626
rect 3130 1623 3156 1626
rect 3226 1623 3244 1626
rect 3396 1623 3421 1626
rect 2826 1616 2829 1623
rect 2994 1616 2997 1623
rect 3418 1616 3421 1623
rect 108 1613 133 1616
rect 178 1613 196 1616
rect 180 1603 189 1606
rect 202 1605 205 1616
rect 244 1613 269 1616
rect 306 1613 324 1616
rect 330 1613 348 1616
rect 420 1613 429 1616
rect 468 1613 493 1616
rect 538 1613 572 1616
rect 604 1613 621 1616
rect 732 1613 741 1616
rect 786 1613 812 1616
rect 850 1613 876 1616
rect 964 1613 989 1616
rect 1026 1613 1060 1616
rect 1106 1613 1132 1616
rect 1276 1613 1325 1616
rect 1340 1613 1349 1616
rect 1388 1613 1421 1616
rect 1474 1613 1492 1616
rect 1588 1613 1637 1616
rect 1674 1613 1684 1616
rect 1722 1613 1756 1616
rect 1786 1613 1812 1616
rect 1874 1613 1916 1616
rect 1962 1613 1980 1616
rect 2076 1613 2132 1616
rect 2236 1613 2253 1616
rect 2292 1613 2324 1616
rect 2420 1613 2445 1616
rect 2476 1613 2485 1616
rect 2554 1613 2580 1616
rect 2714 1613 2724 1616
rect 2738 1613 2780 1616
rect 2826 1613 2852 1616
rect 2916 1613 2941 1616
rect 2994 1613 3005 1616
rect 3194 1613 3212 1616
rect 3234 1613 3252 1616
rect 3290 1613 3316 1616
rect 3340 1613 3381 1616
rect 3418 1613 3428 1616
rect 3468 1613 3501 1616
rect 3532 1613 3549 1616
rect 3674 1613 3692 1616
rect 3898 1613 3948 1616
rect 3978 1613 4020 1616
rect 4058 1613 4076 1616
rect 4114 1613 4148 1616
rect 4186 1613 4220 1616
rect 4250 1613 4300 1616
rect 4338 1613 4380 1616
rect 4532 1613 4604 1616
rect 1722 1606 1725 1613
rect 1962 1606 1965 1613
rect 332 1603 349 1606
rect 386 1603 396 1606
rect 540 1603 573 1606
rect 596 1603 613 1606
rect 740 1603 765 1606
rect 780 1603 813 1606
rect 1068 1603 1133 1606
rect 1156 1603 1221 1606
rect 1242 1603 1252 1606
rect 1284 1603 1333 1606
rect 1348 1603 1357 1606
rect 1668 1603 1685 1606
rect 1708 1603 1725 1606
rect 1914 1603 1924 1606
rect 1940 1603 1965 1606
rect 2004 1603 2013 1606
rect 2018 1603 2060 1606
rect 2298 1603 2332 1606
rect 2714 1603 2732 1606
rect 2738 1596 2741 1613
rect 3002 1607 3005 1613
rect 3378 1607 3381 1613
rect 2754 1603 2772 1606
rect 2860 1603 2869 1606
rect 2882 1603 2908 1606
rect 3028 1603 3061 1606
rect 3108 1603 3125 1606
rect 3274 1603 3324 1606
rect 3498 1603 3501 1613
rect 3722 1603 3764 1606
rect 3900 1603 3940 1606
rect 4050 1603 4068 1606
rect 4178 1603 4212 1606
rect 4324 1603 4333 1606
rect 4338 1603 4372 1606
rect 4482 1603 4508 1606
rect 2340 1593 2365 1596
rect 2716 1593 2725 1596
rect 2738 1595 2749 1596
rect 2740 1593 2749 1595
rect 3482 1593 3508 1596
rect 38 1567 4829 1573
rect 890 1543 916 1546
rect 930 1543 996 1546
rect 3514 1543 3556 1546
rect 170 1533 188 1536
rect 324 1533 357 1536
rect 386 1533 420 1536
rect 570 1533 596 1536
rect 612 1533 660 1536
rect 692 1533 709 1536
rect 818 1533 852 1536
rect 914 1533 924 1536
rect 1004 1533 1013 1536
rect 1194 1533 1236 1536
rect 1258 1533 1308 1536
rect 1340 1533 1404 1536
rect 1434 1533 1452 1536
rect 1722 1533 1740 1536
rect 1930 1533 1948 1536
rect 1970 1533 1988 1536
rect 2866 1533 2892 1536
rect 3058 1533 3084 1536
rect 3098 1533 3108 1536
rect 3132 1533 3149 1536
rect 3186 1533 3196 1536
rect 3324 1533 3333 1536
rect 3338 1533 3348 1536
rect 3458 1533 3476 1536
rect 3508 1533 3557 1536
rect 3586 1533 3604 1536
rect 3684 1533 3693 1536
rect 3706 1533 3716 1536
rect 3794 1533 3804 1536
rect 3852 1533 3877 1536
rect 3900 1533 3925 1536
rect 4034 1533 4044 1536
rect 4068 1533 4077 1536
rect 170 1526 173 1533
rect 706 1526 709 1533
rect 1194 1526 1197 1533
rect 1722 1526 1725 1533
rect 108 1523 133 1526
rect 164 1523 173 1526
rect 252 1523 277 1526
rect 322 1523 356 1526
rect 500 1523 517 1526
rect 556 1523 581 1526
rect 706 1523 724 1526
rect 770 1523 780 1526
rect 932 1523 989 1526
rect 1012 1523 1069 1526
rect 1116 1523 1125 1526
rect 1172 1523 1197 1526
rect 1202 1523 1228 1526
rect 1260 1523 1293 1526
rect 1332 1523 1341 1526
rect 1428 1523 1445 1526
rect 1460 1523 1485 1526
rect 1522 1523 1548 1526
rect 1644 1523 1653 1526
rect 1700 1523 1725 1526
rect 1778 1523 1820 1526
rect 1914 1523 1956 1526
rect 2004 1523 2021 1526
rect 2026 1523 2044 1526
rect 2082 1523 2100 1526
rect 2338 1523 2348 1526
rect 2378 1523 2404 1526
rect 2442 1523 2492 1526
rect 2586 1523 2700 1526
rect 2866 1523 2900 1526
rect 2922 1523 2932 1526
rect 3092 1523 3116 1526
rect 3138 1523 3156 1526
rect 3210 1523 3220 1526
rect 3356 1523 3373 1526
rect 3378 1523 3404 1526
rect 3428 1523 3445 1526
rect 3466 1523 3484 1526
rect 3554 1525 3557 1533
rect 3642 1526 3645 1533
rect 3826 1526 3829 1533
rect 4130 1526 4133 1536
rect 4148 1533 4197 1536
rect 4242 1533 4300 1536
rect 4330 1533 4372 1536
rect 4474 1533 4484 1536
rect 4466 1526 4469 1533
rect 4522 1526 4525 1536
rect 4580 1533 4589 1536
rect 4628 1533 4637 1536
rect 3628 1523 3645 1526
rect 3652 1523 3669 1526
rect 3676 1523 3693 1526
rect 3826 1523 3837 1526
rect 3874 1523 3884 1526
rect 3906 1523 3940 1526
rect 4130 1523 4140 1526
rect 4146 1523 4236 1526
rect 4466 1523 4477 1526
rect 4500 1523 4525 1526
rect 4634 1526 4637 1533
rect 4634 1523 4652 1526
rect 4780 1523 4797 1526
rect 3138 1516 3141 1523
rect 3378 1516 3381 1523
rect 2220 1513 2237 1516
rect 2794 1513 2836 1516
rect 2860 1513 2885 1516
rect 3132 1513 3141 1516
rect 3364 1513 3381 1516
rect 3690 1516 3693 1523
rect 3690 1513 3716 1516
rect 3834 1515 3837 1523
rect 3948 1513 3965 1516
rect 4068 1513 4100 1516
rect 4244 1513 4261 1516
rect 4266 1513 4300 1516
rect 4402 1513 4444 1516
rect 2170 1503 2212 1506
rect 2810 1503 2852 1506
rect 14 1467 4853 1473
rect 2188 1423 2197 1426
rect 3068 1423 3093 1426
rect 3138 1423 3148 1426
rect 3666 1423 3685 1426
rect 3706 1423 3716 1426
rect 3804 1423 3821 1426
rect 108 1413 133 1416
rect 178 1413 196 1416
rect 228 1413 268 1416
rect 300 1413 373 1416
rect 444 1413 469 1416
rect 514 1413 524 1416
rect 530 1413 548 1416
rect 554 1413 580 1416
rect 738 1413 764 1416
rect 770 1413 812 1416
rect 892 1413 933 1416
rect 948 1413 997 1416
rect 1020 1413 1093 1416
rect 1100 1413 1125 1416
rect 1130 1413 1188 1416
rect 1220 1413 1277 1416
rect 1420 1413 1445 1416
rect 1476 1413 1509 1416
rect 1546 1413 1572 1416
rect 1674 1413 1700 1416
rect 1732 1413 1757 1416
rect 1770 1413 1780 1416
rect 1874 1413 1908 1416
rect 1922 1413 1972 1416
rect 2004 1413 2036 1416
rect 180 1403 197 1406
rect 242 1403 276 1406
rect 388 1403 405 1406
rect 532 1403 541 1406
rect 556 1403 573 1406
rect 578 1403 588 1406
rect 604 1403 613 1406
rect 642 1403 668 1406
rect 772 1403 813 1406
rect 884 1403 909 1406
rect 940 1403 965 1406
rect 1012 1403 1053 1406
rect 1108 1403 1165 1406
rect 1170 1403 1196 1406
rect 1212 1403 1284 1406
rect 1316 1403 1396 1406
rect 1412 1403 1437 1406
rect 1458 1403 1468 1406
rect 1660 1403 1701 1406
rect 1916 1403 1973 1406
rect 1996 1403 2021 1406
rect 2178 1403 2181 1414
rect 2250 1413 2276 1416
rect 2364 1413 2389 1416
rect 2548 1413 2580 1416
rect 2674 1413 2684 1416
rect 2786 1413 2804 1416
rect 3108 1413 3133 1416
rect 3164 1413 3181 1416
rect 3236 1413 3277 1416
rect 3308 1413 3341 1416
rect 3372 1413 3412 1416
rect 3666 1413 3724 1416
rect 3778 1413 3788 1416
rect 3178 1406 3181 1413
rect 3826 1406 3829 1425
rect 4020 1423 4069 1426
rect 4074 1423 4084 1426
rect 4482 1423 4524 1426
rect 4554 1423 4573 1426
rect 4586 1423 4596 1426
rect 3842 1413 3876 1416
rect 3970 1413 4012 1416
rect 4018 1413 4092 1416
rect 4226 1413 4236 1416
rect 4274 1413 4300 1416
rect 4306 1413 4324 1416
rect 4354 1413 4380 1416
rect 4460 1413 4517 1416
rect 4540 1413 4597 1416
rect 4612 1413 4637 1416
rect 4756 1413 4773 1416
rect 4306 1407 4309 1413
rect 2786 1403 2796 1406
rect 3082 1403 3100 1406
rect 3114 1403 3148 1406
rect 3178 1403 3212 1406
rect 3234 1403 3292 1406
rect 3378 1403 3404 1406
rect 3732 1403 3749 1406
rect 3754 1403 3780 1406
rect 3804 1403 3829 1406
rect 3844 1403 3869 1406
rect 3906 1403 3932 1406
rect 3956 1403 3965 1406
rect 4100 1403 4117 1406
rect 4252 1403 4261 1406
rect 4418 1403 4444 1406
rect 4482 1403 4524 1406
rect 4554 1403 4596 1406
rect 4634 1403 4644 1406
rect 1170 1396 1173 1403
rect 850 1393 876 1396
rect 890 1393 932 1396
rect 946 1393 1004 1396
rect 1162 1393 1173 1396
rect 3308 1393 3325 1396
rect 3330 1393 3348 1396
rect 2938 1383 2973 1386
rect 38 1367 4829 1373
rect 282 1336 285 1346
rect 778 1343 948 1346
rect 1050 1343 1188 1346
rect 3036 1343 3045 1346
rect 4218 1336 4221 1346
rect 260 1333 285 1336
rect 554 1333 564 1336
rect 580 1333 628 1336
rect 660 1333 669 1336
rect 882 1333 956 1336
rect 1036 1333 1181 1336
rect 1196 1333 1229 1336
rect 1234 1333 1252 1336
rect 1268 1333 1293 1336
rect 1418 1333 1436 1336
rect 1468 1333 1477 1336
rect 1594 1333 1612 1336
rect 1684 1333 1725 1336
rect 1748 1333 1781 1336
rect 1956 1333 1997 1336
rect 1418 1326 1421 1333
rect 1474 1326 1477 1333
rect 1778 1326 1781 1333
rect 116 1323 141 1326
rect 178 1323 252 1326
rect 332 1323 341 1326
rect 484 1323 509 1326
rect 540 1323 549 1326
rect 588 1323 613 1326
rect 618 1323 636 1326
rect 674 1323 684 1326
rect 964 1323 1021 1326
rect 1204 1323 1237 1326
rect 1396 1323 1421 1326
rect 1460 1323 1469 1326
rect 1474 1323 1500 1326
rect 1530 1323 1556 1326
rect 1634 1323 1660 1326
rect 1690 1323 1724 1326
rect 1778 1323 1788 1326
rect 1818 1323 1844 1326
rect 1938 1323 1948 1326
rect 1962 1323 1996 1326
rect 2034 1323 2052 1326
rect 2082 1323 2108 1326
rect 2194 1323 2197 1335
rect 2306 1333 2316 1336
rect 2340 1333 2357 1336
rect 2380 1333 2397 1336
rect 2516 1333 2540 1336
rect 2602 1333 2628 1336
rect 2746 1333 2788 1336
rect 2924 1333 2965 1336
rect 2994 1333 3013 1336
rect 3034 1333 3052 1336
rect 3098 1333 3108 1336
rect 3122 1333 3140 1336
rect 3164 1333 3173 1336
rect 3202 1333 3236 1336
rect 3650 1333 3676 1336
rect 3796 1333 3821 1336
rect 4026 1333 4044 1336
rect 4082 1333 4108 1336
rect 4180 1333 4221 1336
rect 4236 1333 4261 1336
rect 4300 1333 4333 1336
rect 4434 1333 4452 1336
rect 4634 1333 4652 1336
rect 4690 1333 4740 1336
rect 4772 1333 4789 1336
rect 2250 1323 2268 1326
rect 2332 1323 2341 1326
rect 2508 1323 2525 1326
rect 2690 1323 2716 1326
rect 2930 1323 2972 1326
rect 2994 1325 2997 1333
rect 3634 1326 3637 1333
rect 4610 1326 4613 1333
rect 3002 1323 3012 1326
rect 3036 1323 3053 1326
rect 3116 1323 3125 1326
rect 3156 1323 3165 1326
rect 3204 1323 3229 1326
rect 3252 1323 3285 1326
rect 3548 1323 3573 1326
rect 3604 1323 3637 1326
rect 3644 1323 3684 1326
rect 3858 1323 3884 1326
rect 3956 1323 3981 1326
rect 4012 1323 4045 1326
rect 4146 1323 4172 1326
rect 4178 1323 4253 1326
rect 4468 1323 4485 1326
rect 4524 1323 4533 1326
rect 4580 1323 4613 1326
rect 1474 1313 1477 1323
rect 3282 1316 3285 1323
rect 2146 1313 2164 1316
rect 2346 1313 2364 1316
rect 3282 1313 3308 1316
rect 4068 1313 4077 1316
rect 4434 1313 4452 1316
rect 14 1267 4853 1273
rect 2996 1223 3013 1226
rect 3026 1223 3044 1226
rect 3068 1223 3189 1226
rect 132 1213 149 1216
rect 188 1213 197 1216
rect 234 1203 237 1214
rect 282 1213 292 1216
rect 370 1213 388 1216
rect 420 1214 477 1216
rect 418 1213 477 1214
rect 516 1213 541 1216
rect 586 1213 612 1216
rect 698 1213 724 1216
rect 778 1213 796 1216
rect 828 1213 837 1216
rect 930 1213 948 1216
rect 1084 1213 1133 1216
rect 1148 1213 1229 1216
rect 1324 1213 1341 1216
rect 1380 1213 1421 1216
rect 1436 1213 1445 1216
rect 1484 1213 1493 1216
rect 1516 1213 1533 1216
rect 1572 1213 1597 1216
rect 1602 1213 1620 1216
rect 1772 1213 1781 1216
rect 1834 1213 1844 1216
rect 2026 1213 2052 1216
rect 2244 1213 2269 1216
rect 2300 1213 2309 1216
rect 2338 1213 2356 1216
rect 2402 1213 2412 1216
rect 2490 1213 2508 1216
rect 2522 1213 2532 1216
rect 2596 1213 2637 1216
rect 2738 1213 2748 1216
rect 2842 1213 2868 1216
rect 2988 1213 3037 1216
rect 3122 1213 3173 1216
rect 3266 1213 3332 1216
rect 3356 1213 3485 1216
rect 3532 1213 3557 1216
rect 3588 1213 3597 1216
rect 3658 1213 3700 1216
rect 3770 1213 3836 1216
rect 3916 1213 3941 1216
rect 4004 1213 4060 1216
rect 4372 1213 4420 1216
rect 4466 1213 4509 1216
rect 4580 1213 4597 1216
rect 4650 1213 4765 1216
rect 260 1203 284 1206
rect 418 1203 421 1213
rect 2306 1207 2309 1213
rect 3770 1206 3773 1213
rect 4650 1207 4653 1213
rect 588 1203 613 1206
rect 650 1203 676 1206
rect 698 1203 716 1206
rect 748 1203 781 1206
rect 826 1203 876 1206
rect 1178 1203 1244 1206
rect 1282 1203 1316 1206
rect 1330 1203 1356 1206
rect 1378 1203 1428 1206
rect 1482 1203 1508 1206
rect 1580 1203 1605 1206
rect 1644 1203 1661 1206
rect 2372 1203 2389 1206
rect 2434 1203 2468 1206
rect 2540 1203 2549 1206
rect 2588 1203 2621 1206
rect 2842 1203 2860 1206
rect 3348 1203 3357 1206
rect 3602 1203 3612 1206
rect 3644 1203 3677 1206
rect 3682 1203 3692 1206
rect 3724 1203 3773 1206
rect 4330 1203 4348 1206
rect 4468 1203 4501 1206
rect 4562 1203 4572 1206
rect 4586 1203 4620 1206
rect 4724 1203 4789 1206
rect 1090 1193 1132 1196
rect 2436 1193 2453 1196
rect 2484 1193 2501 1196
rect 3322 1193 3332 1196
rect 38 1167 4829 1173
rect 874 1143 908 1146
rect 922 1143 940 1146
rect 4218 1136 4221 1146
rect 156 1133 205 1136
rect 186 1123 204 1126
rect 234 1125 237 1136
rect 250 1133 260 1136
rect 394 1133 444 1136
rect 812 1133 837 1136
rect 860 1133 877 1136
rect 916 1133 933 1136
rect 1068 1133 1093 1136
rect 1108 1133 1149 1136
rect 1706 1133 1724 1136
rect 1740 1133 1757 1136
rect 1788 1133 1829 1136
rect 1844 1133 1909 1136
rect 1932 1133 1941 1136
rect 1962 1133 1972 1136
rect 2364 1133 2388 1136
rect 2500 1133 2509 1136
rect 2514 1133 2532 1136
rect 2570 1133 2604 1136
rect 2620 1133 2637 1136
rect 2738 1133 2748 1136
rect 2866 1133 2884 1136
rect 3018 1133 3028 1136
rect 3042 1133 3068 1136
rect 3114 1133 3132 1136
rect 3218 1133 3236 1136
rect 3250 1133 3268 1136
rect 3284 1133 3301 1136
rect 3306 1133 3340 1136
rect 3594 1133 3604 1136
rect 3682 1133 3772 1136
rect 3804 1133 3813 1136
rect 3906 1133 3940 1136
rect 4034 1133 4068 1136
rect 4172 1133 4221 1136
rect 4226 1133 4244 1136
rect 4276 1133 4301 1136
rect 4330 1133 4348 1136
rect 4564 1133 4581 1136
rect 4612 1133 4621 1136
rect 562 1126 565 1133
rect 874 1126 877 1133
rect 3114 1126 3117 1133
rect 3250 1126 3253 1133
rect 3562 1126 3565 1133
rect 4634 1126 4637 1136
rect 306 1123 332 1126
rect 514 1123 556 1126
rect 562 1123 621 1126
rect 724 1123 749 1126
rect 786 1123 804 1126
rect 826 1123 836 1126
rect 874 1123 909 1126
rect 924 1123 941 1126
rect 996 1123 1021 1126
rect 1066 1123 1100 1126
rect 1122 1123 1156 1126
rect 1316 1123 1325 1126
rect 1372 1123 1381 1126
rect 1386 1123 1396 1126
rect 1442 1123 1452 1126
rect 1532 1123 1557 1126
rect 1594 1123 1620 1126
rect 1652 1123 1669 1126
rect 1754 1123 1780 1126
rect 2026 1123 2036 1126
rect 2098 1123 2124 1126
rect 2188 1113 2197 1116
rect 2218 1113 2236 1116
rect 2242 1106 2245 1125
rect 2330 1123 2356 1126
rect 2562 1123 2596 1126
rect 2698 1123 2756 1126
rect 2882 1123 2892 1126
rect 3012 1123 3029 1126
rect 3036 1123 3069 1126
rect 3076 1123 3085 1126
rect 3100 1123 3117 1126
rect 3148 1123 3181 1126
rect 3244 1123 3253 1126
rect 3292 1123 3325 1126
rect 3364 1123 3373 1126
rect 3484 1123 3508 1126
rect 3554 1123 3565 1126
rect 3580 1123 3605 1126
rect 3612 1123 3621 1126
rect 3746 1123 3780 1126
rect 3818 1123 3836 1126
rect 3866 1123 3892 1126
rect 3964 1123 4012 1126
rect 4092 1123 4164 1126
rect 4226 1123 4252 1126
rect 4282 1123 4333 1126
rect 4556 1123 4581 1126
rect 4604 1123 4637 1126
rect 4732 1123 4757 1126
rect 3554 1116 3557 1123
rect 2260 1113 2285 1116
rect 2322 1113 2348 1116
rect 3044 1113 3061 1116
rect 3162 1113 3188 1116
rect 3212 1113 3229 1116
rect 3516 1113 3557 1116
rect 2172 1103 2189 1106
rect 2194 1103 2245 1106
rect 14 1067 4853 1073
rect 2138 1023 2164 1026
rect 2178 1023 2188 1026
rect 3050 1023 3068 1026
rect 4466 1023 4500 1026
rect 164 1013 181 1016
rect 268 1013 285 1016
rect 324 1013 349 1016
rect 500 1013 517 1016
rect 556 1013 597 1016
rect 650 1013 668 1016
rect 714 1013 732 1016
rect 826 1013 844 1016
rect 850 1013 884 1016
rect 988 1013 1013 1016
rect 1044 1013 1085 1016
rect 1124 1013 1149 1016
rect 1188 1013 1221 1016
rect 1252 1013 1261 1016
rect 1378 1013 1404 1016
rect 1436 1013 1445 1016
rect 1458 1013 1476 1016
rect 1522 1013 1532 1016
rect 1570 1013 1580 1016
rect 178 1006 181 1013
rect 714 1006 717 1013
rect 1458 1006 1461 1013
rect 1634 1006 1637 1016
rect 1666 1013 1684 1016
rect 1812 1013 1829 1016
rect 1970 1013 1988 1016
rect 2034 1013 2044 1016
rect 2194 1013 2212 1016
rect 2354 1013 2365 1016
rect 2434 1013 2452 1016
rect 2482 1013 2492 1016
rect 1666 1006 1669 1013
rect 178 1003 204 1006
rect 226 1003 244 1006
rect 578 1003 612 1006
rect 628 1003 660 1006
rect 692 1003 717 1006
rect 852 1003 877 1006
rect 882 1003 892 1006
rect 908 1003 933 1006
rect 1116 1003 1125 1006
rect 1138 1003 1180 1006
rect 1186 1003 1228 1006
rect 1260 1003 1381 1006
rect 1386 1003 1412 1006
rect 1428 1003 1461 1006
rect 1588 1003 1637 1006
rect 1660 1003 1669 1006
rect 1708 1003 1756 1006
rect 1778 1003 1804 1006
rect 1930 1003 1996 1006
rect 2194 1003 2204 1006
rect 2314 1003 2332 1006
rect 2362 1005 2365 1013
rect 2554 1007 2557 1016
rect 2596 1013 2605 1016
rect 2730 1013 2748 1016
rect 3012 1013 3029 1016
rect 3036 1013 3061 1016
rect 3084 1013 3093 1016
rect 3130 1013 3172 1016
rect 3178 1013 3212 1016
rect 3244 1013 3261 1016
rect 3274 1013 3292 1016
rect 3324 1013 3349 1016
rect 3354 1013 3364 1016
rect 3130 1006 3133 1013
rect 3474 1006 3477 1016
rect 3482 1013 3500 1016
rect 3516 1013 3549 1016
rect 3618 1013 3661 1016
rect 3842 1013 3868 1016
rect 3906 1013 3940 1016
rect 3658 1007 3661 1013
rect 4114 1007 4117 1016
rect 4194 1013 4236 1016
rect 4346 1013 4380 1016
rect 4410 1013 4469 1016
rect 4482 1013 4501 1016
rect 4516 1013 4549 1016
rect 4580 1013 4597 1016
rect 4498 1007 4501 1013
rect 2468 1003 2477 1006
rect 2722 1003 2740 1006
rect 2986 1003 3004 1006
rect 3018 1003 3028 1006
rect 3092 1003 3101 1006
rect 3116 1003 3133 1006
rect 3180 1003 3189 1006
rect 3236 1003 3245 1006
rect 3322 1003 3356 1006
rect 3468 1003 3477 1006
rect 3482 1003 3492 1006
rect 3546 1003 3556 1006
rect 3692 1003 3733 1006
rect 3964 1003 4012 1006
rect 4116 1003 4149 1006
rect 4260 1003 4300 1006
rect 4404 1003 4437 1006
rect 4460 1003 4493 1006
rect 4524 1003 4533 1006
rect 4588 1003 4645 1006
rect 4690 1003 4732 1006
rect 4764 1003 4773 1006
rect 1130 993 1172 996
rect 38 967 4829 973
rect 1010 943 1052 946
rect 188 933 197 936
rect 116 923 141 926
rect 186 923 204 926
rect 234 925 237 936
rect 250 933 260 936
rect 596 933 644 936
rect 676 933 717 936
rect 858 933 908 936
rect 924 933 933 936
rect 978 933 988 936
rect 1034 933 1060 936
rect 1098 933 1124 936
rect 1140 933 1165 936
rect 1170 926 1173 944
rect 3026 943 3077 946
rect 3106 936 3109 944
rect 1180 933 1189 936
rect 1194 933 1220 936
rect 1252 933 1285 936
rect 1412 933 1429 936
rect 1450 933 1508 936
rect 1530 933 1588 936
rect 1668 933 1701 936
rect 2234 933 2252 936
rect 2276 933 2285 936
rect 2306 933 2316 936
rect 2340 933 2349 936
rect 2500 933 2509 936
rect 2522 933 2532 936
rect 2578 933 2604 936
rect 2730 933 2748 936
rect 2866 933 2996 936
rect 3066 933 3092 936
rect 3106 933 3132 936
rect 3218 933 3236 936
rect 3258 933 3332 936
rect 3370 933 3380 936
rect 3498 933 3532 936
rect 3578 933 3588 936
rect 3652 933 3661 936
rect 3666 933 3692 936
rect 3716 933 3725 936
rect 3804 933 3853 936
rect 242 923 268 926
rect 316 923 341 926
rect 378 923 396 926
rect 524 923 557 926
rect 604 923 637 926
rect 756 923 781 926
rect 818 923 844 926
rect 866 923 900 926
rect 970 923 996 926
rect 1068 923 1109 926
rect 1162 923 1173 926
rect 1188 923 1213 926
rect 1244 923 1261 926
rect 1162 913 1165 923
rect 1426 883 1429 933
rect 1516 923 1525 926
rect 1604 923 1629 926
rect 1666 923 1716 926
rect 1746 923 1804 926
rect 1834 923 1860 926
rect 1898 923 1916 926
rect 1962 923 1972 926
rect 2106 913 2156 916
rect 2170 906 2173 925
rect 2194 913 2204 916
rect 2210 906 2213 925
rect 2234 916 2237 933
rect 3626 926 3629 933
rect 3754 926 3757 933
rect 3898 926 3901 933
rect 3946 926 3949 936
rect 4028 933 4045 936
rect 4108 933 4149 936
rect 4180 933 4189 936
rect 4194 933 4228 936
rect 4258 933 4284 936
rect 2300 923 2317 926
rect 2460 923 2485 926
rect 2562 923 2596 926
rect 2746 923 2756 926
rect 3004 923 3077 926
rect 3210 923 3228 926
rect 3260 923 3293 926
rect 3356 923 3373 926
rect 3556 923 3573 926
rect 3626 923 3637 926
rect 3754 923 3765 926
rect 3778 923 3796 926
rect 3802 923 3868 926
rect 3890 923 3901 926
rect 3916 923 3949 926
rect 3994 926 3997 933
rect 4074 926 4077 933
rect 4154 926 4157 933
rect 4314 926 4317 936
rect 4322 933 4340 936
rect 4386 926 4389 936
rect 4394 933 4404 936
rect 4508 933 4541 936
rect 4588 933 4605 936
rect 4610 933 4636 936
rect 3994 923 4005 926
rect 4010 923 4020 926
rect 4074 923 4085 926
rect 4090 923 4100 926
rect 4130 923 4157 926
rect 4300 923 4317 926
rect 4356 923 4389 926
rect 4420 923 4429 926
rect 4500 923 4549 926
rect 4652 923 4669 926
rect 4716 923 4741 926
rect 4780 923 4797 926
rect 2228 913 2237 916
rect 2314 915 2317 923
rect 3114 913 3132 916
rect 3188 913 3221 916
rect 3634 915 3637 923
rect 3762 916 3765 923
rect 3890 916 3893 923
rect 3762 913 3788 916
rect 3876 913 3893 916
rect 4002 916 4005 923
rect 4082 916 4085 923
rect 4002 913 4012 916
rect 4082 913 4092 916
rect 4194 913 4228 916
rect 4314 913 4340 916
rect 4370 913 4404 916
rect 4594 913 4636 916
rect 2170 903 2213 906
rect 2234 903 2237 913
rect 14 867 4853 873
rect 3028 823 3045 826
rect 3090 823 3100 826
rect 3124 823 3189 826
rect 3524 823 3533 826
rect 4172 823 4189 826
rect 108 813 133 816
rect 170 813 180 816
rect 266 813 388 816
rect 420 813 437 816
rect 476 813 501 816
rect 564 813 581 816
rect 668 813 685 816
rect 714 813 732 816
rect 762 813 796 816
rect 826 813 836 816
rect 868 813 885 816
rect 1044 813 1061 816
rect 1180 813 1197 816
rect 1284 813 1317 816
rect 1354 813 1396 816
rect 1442 813 1452 816
rect 1524 813 1549 816
rect 1626 813 1636 816
rect 1674 813 1716 816
rect 1748 813 1757 816
rect 1826 813 1852 816
rect 1940 813 1957 816
rect 1978 813 1996 816
rect 2042 813 2068 816
rect 2186 813 2212 816
rect 2252 813 2277 816
rect 2308 813 2317 816
rect 2548 813 2581 816
rect 682 806 685 813
rect 188 803 205 806
rect 226 803 236 806
rect 252 803 277 806
rect 370 803 396 806
rect 586 803 596 806
rect 612 803 637 806
rect 682 803 692 806
rect 756 803 781 806
rect 820 803 837 806
rect 866 803 900 806
rect 1036 803 1053 806
rect 1066 803 1076 806
rect 1186 803 1220 806
rect 1236 803 1261 806
rect 1282 803 1324 806
rect 1354 805 1357 813
rect 2618 806 2621 814
rect 2626 813 2644 816
rect 2738 813 2756 816
rect 2850 813 2868 816
rect 3020 813 3061 816
rect 3228 813 3260 816
rect 3292 813 3333 816
rect 3436 813 3477 816
rect 3498 813 3516 816
rect 3556 813 3589 816
rect 3612 813 3653 816
rect 3714 813 3732 816
rect 3746 813 3796 816
rect 3834 813 3876 816
rect 3906 813 3948 816
rect 4044 813 4085 816
rect 4122 813 4164 816
rect 4170 813 4244 816
rect 4282 813 4316 816
rect 4410 813 4452 816
rect 4506 813 4516 816
rect 1596 803 1637 806
rect 1660 803 1724 806
rect 1746 803 1780 806
rect 1898 803 1916 806
rect 1938 803 1956 806
rect 1970 803 2004 806
rect 2034 803 2060 806
rect 2194 803 2204 806
rect 2570 803 2596 806
rect 2618 803 2637 806
rect 2850 803 2860 806
rect 2978 803 3012 806
rect 3050 803 3060 806
rect 3220 803 3229 806
rect 3290 803 3332 806
rect 3386 803 3412 806
rect 3570 803 3604 806
rect 3626 803 3676 806
rect 3740 803 3781 806
rect 3820 803 3861 806
rect 3900 803 3909 806
rect 3972 803 4020 806
rect 4052 803 4077 806
rect 4082 803 4092 806
rect 4354 803 4372 806
rect 4482 803 4508 806
rect 4602 803 4628 806
rect 4660 803 4677 806
rect 1010 793 1028 796
rect 38 767 4829 773
rect 1010 743 1020 746
rect 1034 743 1060 746
rect 2484 743 2525 746
rect 3130 743 3156 746
rect 188 733 221 736
rect 226 733 236 736
rect 404 733 429 736
rect 116 723 141 726
rect 210 723 244 726
rect 324 723 349 726
rect 386 723 396 726
rect 458 725 461 736
rect 466 733 492 736
rect 564 733 573 736
rect 586 733 604 736
rect 748 733 765 736
rect 804 733 829 736
rect 1180 733 1213 736
rect 1242 733 1284 736
rect 1644 733 1676 736
rect 1708 733 1733 736
rect 1898 733 1932 736
rect 2290 733 2308 736
rect 2332 733 2405 736
rect 2450 733 2461 736
rect 754 726 757 733
rect 500 723 517 726
rect 522 723 540 726
rect 572 723 621 726
rect 716 723 725 726
rect 754 723 780 726
rect 810 723 836 726
rect 868 723 876 726
rect 882 723 900 726
rect 938 723 964 726
rect 1036 723 1053 726
rect 1076 723 1117 726
rect 1122 723 1172 726
rect 1178 723 1212 726
rect 1244 723 1261 726
rect 1330 723 1356 726
rect 1394 723 1428 726
rect 1474 723 1484 726
rect 1706 723 1757 726
rect 1892 723 1909 726
rect 1914 723 1924 726
rect 2074 723 2092 726
rect 2138 723 2148 726
rect 2324 723 2373 726
rect 2378 723 2412 726
rect 2458 725 2461 733
rect 2522 726 2525 743
rect 2540 733 2549 736
rect 2586 733 2612 736
rect 2812 733 2860 736
rect 2890 733 2940 736
rect 3074 733 3108 736
rect 3138 733 3164 736
rect 3514 733 3532 736
rect 3586 733 3596 736
rect 3660 733 3709 736
rect 3772 733 3781 736
rect 3786 733 3812 736
rect 4098 733 4164 736
rect 4298 733 4332 736
rect 4452 733 4469 736
rect 4610 733 4644 736
rect 4690 733 4716 736
rect 4772 733 4789 736
rect 3074 726 3077 733
rect 2522 723 2532 726
rect 2586 723 2604 726
rect 2642 723 2652 726
rect 2762 723 2788 726
rect 2948 723 2981 726
rect 2988 723 2997 726
rect 3012 723 3045 726
rect 3060 723 3077 726
rect 3124 723 3149 726
rect 3210 723 3236 726
rect 3404 723 3413 726
rect 3540 723 3581 726
rect 3594 723 3636 726
rect 3674 723 3748 726
rect 3786 723 3820 726
rect 3978 723 4172 726
rect 4210 723 4268 726
rect 4298 723 4340 726
rect 4522 723 4580 726
rect 4634 723 4652 726
rect 4706 723 4724 726
rect 4754 723 4764 726
rect 2378 716 2381 723
rect 2058 713 2077 716
rect 2354 713 2381 716
rect 2956 713 2973 716
rect 3018 713 3044 716
rect 3204 713 3221 716
rect 14 667 4853 673
rect 2980 633 3013 636
rect 2338 623 2356 626
rect 330 613 356 616
rect 362 613 388 616
rect 578 613 604 616
rect 668 613 677 616
rect 786 613 836 616
rect 890 613 924 616
rect 954 613 980 616
rect 1100 613 1125 616
rect 1170 613 1180 616
rect 1212 613 1244 616
rect 1250 613 1269 616
rect 1402 613 1420 616
rect 1452 613 1461 616
rect 1468 613 1477 616
rect 1618 613 1644 616
rect 1722 613 1740 616
rect 1772 613 1780 616
rect 1906 613 1916 616
rect 2244 613 2269 616
rect 2300 613 2317 616
rect 2394 613 2412 616
rect 2458 613 2468 616
rect 2642 613 2684 616
rect 2898 613 2908 616
rect 3002 613 3020 616
rect 3508 613 3533 616
rect 3540 613 3581 616
rect 3634 613 3644 616
rect 3778 613 3804 616
rect 4146 613 4196 616
rect 4338 613 4388 616
rect 4474 613 4524 616
rect 4554 613 4564 616
rect 4666 613 4716 616
rect 890 606 893 613
rect 180 603 189 606
rect 202 603 212 606
rect 228 603 245 606
rect 266 603 300 606
rect 316 603 341 606
rect 364 603 389 606
rect 602 603 612 606
rect 634 603 660 606
rect 818 603 844 606
rect 860 603 893 606
rect 1172 603 1181 606
rect 1250 605 1253 613
rect 1258 603 1284 606
rect 1316 603 1349 606
rect 1394 603 1428 606
rect 1450 603 1460 606
rect 1474 603 1516 606
rect 1716 603 1733 606
rect 1770 603 1788 606
rect 2306 603 2356 606
rect 2380 603 2413 606
rect 2458 596 2461 613
rect 2476 603 2517 606
rect 2556 603 2596 606
rect 2644 603 2661 606
rect 2802 603 2828 606
rect 3028 603 3045 606
rect 3092 603 3117 606
rect 3162 603 3172 606
rect 3178 603 3268 606
rect 3282 603 3292 606
rect 3530 605 3533 613
rect 3634 606 3637 613
rect 3620 603 3637 606
rect 3658 603 3676 606
rect 3812 603 3837 606
rect 3922 603 3956 606
rect 4068 603 4109 606
rect 4220 603 4229 606
rect 4500 603 4509 606
rect 4594 603 4628 606
rect 4724 603 4789 606
rect 1018 593 1044 596
rect 2436 593 2461 596
rect 3180 593 3237 596
rect 3274 593 3284 596
rect 38 567 4829 573
rect 978 543 1012 546
rect 1026 543 1036 546
rect 1178 543 1196 546
rect 1210 543 1244 546
rect 2970 543 2988 546
rect 162 533 180 536
rect 202 533 220 536
rect 364 533 389 536
rect 442 533 452 536
rect 210 523 228 526
rect 292 523 317 526
rect 362 523 388 526
rect 420 523 437 526
rect 564 523 589 526
rect 626 525 629 536
rect 658 525 661 536
rect 730 533 756 536
rect 788 533 813 536
rect 842 533 852 536
rect 866 533 916 536
rect 938 533 964 536
rect 1044 533 1061 536
rect 1204 533 1237 536
rect 1258 533 1276 536
rect 1308 533 1325 536
rect 1386 533 1396 536
rect 1418 533 1444 536
rect 1586 533 1596 536
rect 1636 533 1669 536
rect 1708 533 1773 536
rect 1970 533 2012 536
rect 1666 526 1669 533
rect 666 523 676 526
rect 730 523 764 526
rect 794 523 812 526
rect 850 523 860 526
rect 866 523 908 526
rect 940 523 957 526
rect 962 523 972 526
rect 1028 523 1037 526
rect 1052 523 1069 526
rect 1108 523 1133 526
rect 1164 523 1189 526
rect 1212 523 1245 526
rect 1260 523 1269 526
rect 1300 523 1309 526
rect 1410 523 1436 526
rect 1522 523 1532 526
rect 1612 523 1620 526
rect 1666 523 1684 526
rect 1796 523 1845 526
rect 1946 523 1964 526
rect 1970 523 2004 526
rect 2034 525 2037 536
rect 2042 533 2060 536
rect 2314 533 2348 536
rect 2362 533 2388 536
rect 2436 533 2445 536
rect 2898 533 2916 536
rect 2964 533 2973 536
rect 2978 533 2996 536
rect 3394 533 3436 536
rect 3490 533 3524 536
rect 3724 533 3756 536
rect 3788 533 3844 536
rect 3858 533 3884 536
rect 3970 533 4004 536
rect 4058 533 4076 536
rect 3858 526 3861 533
rect 4226 526 4229 534
rect 4276 533 4293 536
rect 4628 533 4645 536
rect 2068 523 2093 526
rect 2130 523 2156 526
rect 2338 523 2356 526
rect 2386 523 2412 526
rect 2484 523 2501 526
rect 2924 523 2956 526
rect 3004 523 3021 526
rect 3060 523 3109 526
rect 3260 523 3293 526
rect 3388 523 3429 526
rect 3444 523 3453 526
rect 3532 523 3549 526
rect 3556 523 3565 526
rect 3604 523 3629 526
rect 3786 523 3861 526
rect 3908 523 3956 526
rect 4050 523 4084 526
rect 4140 523 4165 526
rect 4196 523 4229 526
rect 4236 523 4252 526
rect 4410 523 4436 526
rect 4538 523 4564 526
rect 4620 523 4637 526
rect 4780 523 4789 526
rect 794 513 797 523
rect 2364 513 2381 516
rect 3066 513 3116 516
rect 3540 513 3548 516
rect 14 467 4853 473
rect 3036 433 3053 436
rect 2938 423 2972 426
rect 3018 423 3028 426
rect 3404 423 3413 426
rect 108 413 133 416
rect 220 413 285 416
rect 324 413 349 416
rect 380 413 397 416
rect 426 406 429 414
rect 602 413 612 416
rect 676 413 685 416
rect 730 413 740 416
rect 778 413 796 416
rect 890 413 908 416
rect 1036 413 1045 416
rect 1084 413 1109 416
rect 1140 413 1157 416
rect 1196 413 1221 416
rect 1450 413 1460 416
rect 1570 413 1596 416
rect 1762 413 1772 416
rect 1842 413 1868 416
rect 1972 413 1981 416
rect 2068 413 2093 416
rect 2130 413 2156 416
rect 2332 413 2357 416
rect 2474 413 2492 416
rect 2538 413 2556 416
rect 2820 413 2837 416
rect 2980 413 2996 416
rect 3044 413 3060 416
rect 3066 413 3092 416
rect 3196 413 3213 416
rect 3252 413 3261 416
rect 3308 413 3341 416
rect 3356 413 3381 416
rect 3402 413 3460 416
rect 3474 413 3485 416
rect 3506 413 3525 416
rect 3588 413 3613 416
rect 3644 413 3685 416
rect 4004 413 4021 416
rect 4106 413 4132 416
rect 4252 413 4277 416
rect 4314 413 4348 416
rect 4378 413 4413 416
rect 4444 413 4461 416
rect 4604 413 4629 416
rect 4634 413 4668 416
rect 778 406 781 413
rect 180 403 189 406
rect 386 403 429 406
rect 458 403 484 406
rect 594 403 620 406
rect 642 403 668 406
rect 722 403 732 406
rect 764 403 781 406
rect 1162 403 1172 406
rect 1202 403 1244 406
rect 1266 403 1276 406
rect 1314 403 1332 406
rect 1442 403 1468 406
rect 1490 403 1524 406
rect 1652 403 1685 406
rect 1730 403 1780 406
rect 1796 403 1805 406
rect 1906 403 1948 406
rect 1964 403 2004 406
rect 2020 403 2029 406
rect 2034 403 2060 406
rect 2338 403 2381 406
rect 2994 403 3004 406
rect 3068 403 3085 406
rect 3314 403 3348 406
rect 3362 403 3388 406
rect 3418 403 3452 406
rect 3474 405 3477 413
rect 3506 405 3509 413
rect 4410 406 4413 413
rect 3514 403 3524 406
rect 3650 403 3692 406
rect 4330 403 4340 406
rect 4410 403 4420 406
rect 4628 403 4653 406
rect 1002 393 1020 396
rect 38 367 4829 373
rect 794 343 828 346
rect 970 343 1020 346
rect 2674 343 2692 346
rect 354 333 380 336
rect 580 333 605 336
rect 746 333 756 336
rect 788 333 821 336
rect 842 333 876 336
rect 906 333 932 336
rect 946 333 964 336
rect 1010 333 1028 336
rect 1100 333 1125 336
rect 1140 333 1181 336
rect 1186 333 1204 336
rect 1236 333 1245 336
rect 1300 333 1325 336
rect 1346 333 1356 336
rect 1764 333 1773 336
rect 1812 333 1845 336
rect 1970 333 2020 336
rect 2042 333 2092 336
rect 2516 333 2541 336
rect 2594 333 2612 336
rect 2660 333 2669 336
rect 2700 333 2733 336
rect 2844 333 2861 336
rect 2884 333 2925 336
rect 3068 333 3085 336
rect 3114 333 3132 336
rect 3290 333 3340 336
rect 3362 333 3372 336
rect 3426 333 3452 336
rect 3466 333 3492 336
rect 3522 333 3532 336
rect 3556 333 3573 336
rect 3610 333 3636 336
rect 3924 333 3948 336
rect 3980 333 4004 336
rect 4108 333 4148 336
rect 108 323 133 326
rect 164 323 181 326
rect 276 323 301 326
rect 338 323 348 326
rect 492 323 517 326
rect 554 323 572 326
rect 578 323 604 326
rect 844 323 861 326
rect 900 323 917 326
rect 940 323 949 326
rect 972 323 1021 326
rect 1036 323 1085 326
rect 1106 323 1132 326
rect 1394 323 1420 326
rect 1514 323 1524 326
rect 1636 323 1645 326
rect 1826 323 1852 326
rect 1946 323 1964 326
rect 1970 323 2012 326
rect 2044 323 2061 326
rect 2164 323 2173 326
rect 2276 323 2301 326
rect 2474 323 2500 326
rect 2620 323 2645 326
rect 2652 323 2661 326
rect 2772 323 2797 326
rect 2858 325 2861 333
rect 3020 323 3029 326
rect 3036 323 3045 326
rect 3074 323 3092 326
rect 3140 323 3157 326
rect 3252 323 3261 326
rect 3268 323 3277 326
rect 3290 325 3293 333
rect 4402 326 4405 335
rect 4426 333 4444 336
rect 4666 333 4692 336
rect 4740 333 4789 336
rect 3348 323 3357 326
rect 3380 323 3389 326
rect 3460 323 3500 326
rect 3522 323 3540 326
rect 3588 323 3644 326
rect 3698 323 3716 326
rect 3796 323 3821 326
rect 3858 323 3900 326
rect 3972 323 4005 326
rect 4100 323 4117 326
rect 4130 323 4156 326
rect 4340 323 4365 326
rect 4396 323 4405 326
rect 4412 323 4452 326
rect 4732 323 4741 326
rect 2516 313 2556 316
rect 2580 313 2589 316
rect 2564 303 2597 306
rect 14 267 4853 273
rect 3348 223 3365 226
rect 3396 223 3405 226
rect 3436 223 3453 226
rect 108 213 133 216
rect 260 213 268 216
rect 426 213 436 216
rect 474 213 492 216
rect 530 213 540 216
rect 572 213 644 216
rect 676 213 693 216
rect 700 213 709 216
rect 714 213 724 216
rect 828 213 853 216
rect 868 213 885 216
rect 890 213 900 216
rect 946 213 956 216
rect 1002 213 1012 216
rect 1148 213 1157 216
rect 1242 213 1292 216
rect 1338 213 1348 216
rect 1452 213 1461 216
rect 1466 213 1492 216
rect 1636 213 1669 216
rect 1684 213 1701 216
rect 1706 213 1716 216
rect 1748 213 1772 216
rect 1820 213 1845 216
rect 1892 213 1909 216
rect 1940 213 1957 216
rect 1962 213 1972 216
rect 2010 213 2044 216
rect 2146 213 2164 216
rect 2210 213 2220 216
rect 2300 213 2325 216
rect 2356 213 2373 216
rect 2490 213 2508 216
rect 2522 213 2540 216
rect 2682 213 2708 216
rect 2818 213 2844 216
rect 2850 213 2900 216
rect 2938 213 2972 216
rect 2978 213 2988 216
rect 3082 213 3092 216
rect 3316 213 3333 216
rect 3340 213 3349 216
rect 3394 213 3420 216
rect 3460 213 3477 216
rect 3516 213 3541 216
rect 3572 213 3581 216
rect 3586 213 3620 216
rect 3730 213 3772 216
rect 3802 213 3820 216
rect 3916 213 3941 216
rect 4100 213 4125 216
rect 4282 213 4292 216
rect 4340 213 4356 216
rect 4452 213 4468 216
rect 4564 213 4580 216
rect 4586 213 4645 216
rect 2682 206 2685 213
rect 180 203 189 206
rect 212 203 221 206
rect 226 203 236 206
rect 298 203 316 206
rect 338 203 356 206
rect 372 203 381 206
rect 466 203 484 206
rect 564 203 645 206
rect 674 203 692 206
rect 788 203 813 206
rect 826 203 860 206
rect 1004 203 1013 206
rect 1162 203 1172 206
rect 1194 203 1204 206
rect 1236 203 1285 206
rect 1386 203 1412 206
rect 1434 203 1444 206
rect 1466 203 1500 206
rect 1522 203 1564 206
rect 1596 203 1605 206
rect 1690 203 1724 206
rect 1740 203 1757 206
rect 1802 203 1812 206
rect 1826 203 1868 206
rect 1884 203 1917 206
rect 1946 203 1980 206
rect 2474 203 2500 206
rect 2514 203 2532 206
rect 2562 203 2596 206
rect 2626 203 2644 206
rect 2660 203 2685 206
rect 2722 203 2748 206
rect 2812 203 2837 206
rect 2850 205 2853 213
rect 2866 203 2908 206
rect 2978 205 2981 213
rect 3330 205 3333 213
rect 4642 206 4645 213
rect 3346 203 3380 206
rect 3442 203 3452 206
rect 3578 203 3612 206
rect 3644 203 3700 206
rect 3732 203 3764 206
rect 3778 203 3812 206
rect 3844 203 3892 206
rect 4276 203 4285 206
rect 4306 203 4316 206
rect 4364 203 4397 206
rect 4402 203 4428 206
rect 4476 203 4509 206
rect 4514 203 4540 206
rect 4588 203 4613 206
rect 4642 203 4660 206
rect 794 193 812 196
rect 826 193 852 196
rect 38 167 4829 173
rect 826 133 844 136
rect 1156 133 1165 136
rect 1218 133 1244 136
rect 1266 133 1284 136
rect 2458 135 2468 136
rect 2458 133 2469 135
rect 2466 126 2469 133
rect 2746 126 2749 135
rect 2930 126 2933 135
rect 3330 126 3333 135
rect 3570 126 3573 135
rect 3746 126 3749 135
rect 4036 133 4061 136
rect 4074 126 4077 135
rect 172 123 197 126
rect 292 123 301 126
rect 474 123 484 126
rect 548 123 557 126
rect 770 123 796 126
rect 828 123 845 126
rect 890 123 916 126
rect 988 123 997 126
rect 1084 123 1109 126
rect 1196 123 1205 126
rect 1330 123 1356 126
rect 1458 123 1468 126
rect 1618 123 1628 126
rect 1778 123 1796 126
rect 1842 123 1852 126
rect 1898 123 1908 126
rect 1954 123 1964 126
rect 2050 123 2076 126
rect 2388 123 2413 126
rect 2444 123 2469 126
rect 2476 123 2485 126
rect 2684 123 2709 126
rect 2740 123 2749 126
rect 2756 123 2765 126
rect 2780 123 2852 126
rect 2898 123 2924 126
rect 2930 123 2956 126
rect 2986 123 3012 126
rect 3050 123 3108 126
rect 3316 123 3333 126
rect 3340 123 3365 126
rect 3380 123 3389 126
rect 3404 123 3428 126
rect 3492 123 3517 126
rect 3548 123 3573 126
rect 3580 123 3589 126
rect 3652 123 3677 126
rect 3708 123 3749 126
rect 3804 123 3829 126
rect 4028 123 4037 126
rect 4050 123 4068 126
rect 4074 123 4084 126
rect 4114 123 4140 126
rect 4228 123 4253 126
rect 4284 123 4301 126
rect 4668 123 4677 126
rect 2594 113 2628 116
rect 3388 113 3397 116
rect 3444 113 3453 116
rect 14 67 4853 73
rect 38 37 4829 57
rect 14 13 4853 33
<< metal2 >>
rect 2 273 5 3216
rect 14 13 34 4727
rect 38 37 58 4703
rect 1170 4626 1173 4706
rect 1650 4656 1653 4736
rect 1866 4656 1869 4676
rect 1650 4653 1661 4656
rect 90 4593 93 4606
rect 122 4523 125 4616
rect 170 4533 173 4546
rect 170 4513 173 4526
rect 178 4523 181 4606
rect 186 4523 189 4546
rect 82 4366 85 4406
rect 82 4363 93 4366
rect 90 4256 93 4363
rect 82 4253 93 4256
rect 82 4103 85 4253
rect 122 4136 125 4416
rect 130 4413 133 4426
rect 162 4413 165 4436
rect 170 4413 173 4426
rect 178 4386 181 4416
rect 186 4396 189 4406
rect 194 4403 197 4436
rect 218 4416 221 4526
rect 202 4396 205 4416
rect 210 4413 221 4416
rect 186 4393 205 4396
rect 178 4383 189 4386
rect 138 4313 141 4326
rect 170 4303 173 4326
rect 178 4313 181 4326
rect 186 4323 189 4383
rect 218 4366 221 4406
rect 226 4403 229 4526
rect 234 4506 237 4526
rect 266 4523 269 4616
rect 274 4533 277 4556
rect 282 4543 301 4546
rect 282 4523 285 4543
rect 290 4523 293 4536
rect 298 4533 301 4543
rect 298 4513 301 4526
rect 234 4503 245 4506
rect 242 4446 245 4503
rect 234 4443 245 4446
rect 218 4363 229 4366
rect 202 4343 221 4346
rect 202 4333 205 4343
rect 130 4213 133 4226
rect 162 4193 165 4216
rect 170 4213 173 4226
rect 202 4223 205 4326
rect 210 4303 213 4336
rect 218 4323 221 4343
rect 226 4316 229 4363
rect 234 4333 237 4443
rect 242 4386 245 4416
rect 258 4413 261 4426
rect 250 4403 261 4406
rect 266 4403 269 4436
rect 242 4383 269 4386
rect 226 4313 237 4316
rect 162 4143 181 4146
rect 122 4133 133 4136
rect 162 4133 165 4143
rect 82 3886 85 4036
rect 114 4013 117 4126
rect 130 4066 133 4133
rect 162 4113 165 4126
rect 122 4063 133 4066
rect 122 4006 125 4063
rect 114 4003 125 4006
rect 82 3883 93 3886
rect 90 3746 93 3883
rect 82 3743 93 3746
rect 82 3603 85 3743
rect 90 3713 93 3736
rect 106 3613 109 3726
rect 114 3706 117 4003
rect 130 3913 133 3926
rect 146 3923 149 3976
rect 154 3856 157 4026
rect 170 4013 173 4136
rect 178 4123 181 4143
rect 210 4136 213 4216
rect 178 3966 181 4106
rect 186 3973 189 4136
rect 194 4133 213 4136
rect 218 4133 221 4226
rect 226 4196 229 4206
rect 234 4203 237 4313
rect 250 4303 253 4336
rect 242 4196 245 4216
rect 258 4213 261 4226
rect 226 4193 245 4196
rect 250 4193 253 4206
rect 258 4186 261 4206
rect 250 4183 261 4186
rect 194 4123 197 4133
rect 202 4113 205 4126
rect 226 4106 229 4136
rect 218 4103 229 4106
rect 218 4036 221 4103
rect 218 4033 229 4036
rect 194 4013 197 4026
rect 178 3963 197 3966
rect 162 3923 165 3936
rect 178 3933 181 3946
rect 194 3933 197 3963
rect 210 3943 213 4016
rect 218 3933 221 4006
rect 170 3913 173 3926
rect 154 3853 165 3856
rect 122 3723 125 3816
rect 162 3776 165 3853
rect 178 3803 181 3926
rect 226 3916 229 4033
rect 222 3913 229 3916
rect 222 3826 225 3913
rect 222 3823 229 3826
rect 186 3793 189 3816
rect 194 3813 205 3816
rect 154 3773 165 3776
rect 114 3703 125 3706
rect 122 3606 125 3703
rect 114 3603 125 3606
rect 114 3536 117 3603
rect 106 3533 117 3536
rect 106 3466 109 3533
rect 106 3463 117 3466
rect 90 3403 93 3426
rect 114 3366 117 3463
rect 122 3413 125 3526
rect 154 3456 157 3773
rect 162 3723 165 3736
rect 170 3733 173 3746
rect 178 3556 181 3736
rect 186 3713 189 3726
rect 194 3723 197 3806
rect 210 3743 213 3816
rect 218 3733 221 3806
rect 226 3733 229 3823
rect 234 3726 237 4096
rect 242 4073 245 4126
rect 250 4106 253 4183
rect 258 4123 261 4136
rect 250 4103 257 4106
rect 242 4013 245 4056
rect 254 4026 257 4103
rect 250 4023 257 4026
rect 250 4003 253 4023
rect 266 4016 269 4383
rect 282 4223 285 4426
rect 290 4333 293 4356
rect 298 4323 301 4336
rect 306 4333 309 4526
rect 314 4523 317 4616
rect 322 4566 325 4596
rect 346 4593 349 4606
rect 322 4563 333 4566
rect 330 4436 333 4563
rect 370 4513 373 4536
rect 378 4523 381 4606
rect 402 4593 405 4606
rect 426 4603 429 4616
rect 394 4533 397 4546
rect 410 4533 413 4556
rect 386 4503 389 4526
rect 402 4513 405 4526
rect 426 4496 429 4556
rect 322 4433 333 4436
rect 418 4493 429 4496
rect 322 4416 325 4433
rect 318 4413 325 4416
rect 318 4316 321 4413
rect 330 4323 333 4416
rect 386 4323 389 4416
rect 418 4376 421 4493
rect 442 4476 445 4506
rect 434 4473 445 4476
rect 450 4473 453 4526
rect 434 4396 437 4473
rect 450 4413 453 4426
rect 450 4396 453 4406
rect 458 4403 461 4536
rect 466 4483 469 4526
rect 474 4493 477 4536
rect 490 4533 493 4616
rect 546 4613 549 4626
rect 538 4576 541 4606
rect 538 4573 549 4576
rect 490 4496 493 4526
rect 506 4503 509 4526
rect 530 4523 533 4536
rect 538 4496 541 4566
rect 546 4523 549 4573
rect 554 4563 557 4616
rect 586 4613 589 4626
rect 690 4613 693 4626
rect 730 4613 733 4626
rect 634 4593 637 4606
rect 650 4586 653 4606
rect 706 4593 709 4606
rect 634 4583 653 4586
rect 554 4533 557 4556
rect 490 4493 501 4496
rect 466 4396 469 4416
rect 482 4413 485 4476
rect 498 4413 501 4493
rect 530 4493 541 4496
rect 434 4393 445 4396
rect 450 4393 469 4396
rect 474 4393 477 4406
rect 418 4373 429 4376
rect 426 4356 429 4373
rect 426 4353 433 4356
rect 318 4313 325 4316
rect 282 4203 285 4216
rect 282 4176 285 4196
rect 282 4173 293 4176
rect 274 4133 277 4156
rect 282 4093 285 4166
rect 290 4133 293 4173
rect 306 4163 309 4226
rect 298 4086 301 4136
rect 282 4083 301 4086
rect 266 4013 277 4016
rect 282 4013 285 4083
rect 242 3813 245 3926
rect 274 3856 277 4013
rect 298 3946 301 4076
rect 306 4023 309 4126
rect 322 4033 325 4313
rect 330 4213 333 4226
rect 362 4193 365 4216
rect 370 4213 373 4226
rect 386 4156 389 4176
rect 386 4153 393 4156
rect 370 4113 373 4126
rect 390 4086 393 4153
rect 402 4143 405 4216
rect 410 4136 413 4336
rect 430 4306 433 4353
rect 426 4303 433 4306
rect 418 4213 421 4226
rect 418 4196 421 4206
rect 426 4203 429 4303
rect 442 4296 445 4393
rect 522 4366 525 4406
rect 530 4403 533 4493
rect 554 4413 557 4486
rect 546 4393 549 4406
rect 522 4363 529 4366
rect 458 4323 461 4336
rect 442 4293 453 4296
rect 434 4196 437 4216
rect 418 4193 437 4196
rect 442 4193 445 4206
rect 410 4133 421 4136
rect 402 4103 405 4126
rect 410 4113 413 4126
rect 386 4083 393 4086
rect 386 4046 389 4083
rect 418 4076 421 4133
rect 370 4043 389 4046
rect 402 4073 421 4076
rect 322 4013 333 4016
rect 354 4013 357 4026
rect 290 3943 301 3946
rect 274 3853 285 3856
rect 210 3723 237 3726
rect 210 3696 213 3723
rect 202 3693 213 3696
rect 202 3566 205 3693
rect 218 3636 221 3706
rect 218 3633 237 3636
rect 202 3563 213 3566
rect 170 3553 181 3556
rect 170 3506 173 3553
rect 186 3543 205 3546
rect 186 3533 189 3543
rect 186 3513 189 3526
rect 170 3503 181 3506
rect 154 3453 165 3456
rect 162 3376 165 3453
rect 178 3403 181 3503
rect 194 3393 197 3536
rect 202 3523 205 3543
rect 110 3363 117 3366
rect 154 3373 165 3376
rect 98 3323 101 3346
rect 110 3286 113 3363
rect 146 3313 149 3326
rect 110 3283 117 3286
rect 82 2756 85 3206
rect 114 3173 117 3283
rect 130 3203 133 3216
rect 146 3183 149 3236
rect 130 3123 133 3136
rect 98 3003 101 3026
rect 106 2923 109 3016
rect 114 2986 117 3036
rect 130 3013 133 3026
rect 122 2993 125 3006
rect 114 2983 125 2986
rect 74 2753 85 2756
rect 74 2596 77 2753
rect 90 2713 93 2736
rect 106 2723 109 2816
rect 82 2603 85 2626
rect 74 2593 85 2596
rect 82 2506 85 2593
rect 106 2523 109 2616
rect 122 2613 125 2983
rect 138 2966 141 3016
rect 146 3013 149 3176
rect 154 3106 157 3373
rect 210 3366 213 3563
rect 218 3523 221 3633
rect 242 3563 245 3726
rect 250 3723 253 3826
rect 258 3733 261 3776
rect 226 3533 229 3546
rect 206 3363 213 3366
rect 178 3293 181 3336
rect 194 3313 197 3326
rect 206 3306 209 3363
rect 226 3356 229 3526
rect 242 3423 245 3556
rect 266 3546 269 3836
rect 274 3733 277 3816
rect 282 3786 285 3853
rect 290 3813 293 3943
rect 298 3933 309 3936
rect 290 3796 293 3806
rect 298 3803 301 3926
rect 306 3823 309 3926
rect 306 3796 309 3816
rect 314 3813 317 3936
rect 330 3933 333 4013
rect 370 3996 373 4043
rect 402 4003 405 4073
rect 426 4046 429 4146
rect 434 4123 437 4136
rect 450 4133 453 4293
rect 466 4186 469 4216
rect 482 4203 485 4326
rect 506 4313 509 4326
rect 526 4306 529 4363
rect 538 4323 541 4336
rect 562 4333 565 4406
rect 546 4313 549 4326
rect 526 4303 533 4306
rect 530 4256 533 4303
rect 522 4253 533 4256
rect 466 4183 485 4186
rect 458 4143 477 4146
rect 458 4133 461 4143
rect 466 4103 469 4136
rect 474 4123 477 4143
rect 482 4123 485 4183
rect 498 4113 501 4126
rect 506 4123 509 4216
rect 522 4176 525 4253
rect 570 4203 573 4406
rect 578 4303 581 4426
rect 586 4383 589 4526
rect 586 4313 589 4336
rect 586 4203 589 4216
rect 522 4173 541 4176
rect 538 4146 541 4173
rect 530 4143 541 4146
rect 422 4043 429 4046
rect 370 3993 381 3996
rect 322 3833 325 3926
rect 290 3793 309 3796
rect 282 3783 289 3786
rect 286 3706 289 3783
rect 314 3766 317 3806
rect 322 3793 325 3806
rect 314 3763 333 3766
rect 286 3703 293 3706
rect 290 3566 293 3703
rect 306 3613 309 3756
rect 286 3563 293 3566
rect 266 3543 277 3546
rect 266 3523 269 3536
rect 274 3416 277 3543
rect 286 3486 289 3563
rect 330 3543 333 3763
rect 338 3676 341 3956
rect 362 3933 365 3956
rect 378 3946 381 3993
rect 422 3986 425 4043
rect 490 4013 493 4026
rect 422 3983 429 3986
rect 426 3966 429 3983
rect 426 3963 433 3966
rect 378 3943 397 3946
rect 394 3896 397 3943
rect 410 3913 413 3926
rect 386 3893 397 3896
rect 386 3836 389 3893
rect 430 3886 433 3963
rect 442 3953 445 4006
rect 530 3966 533 4143
rect 546 4133 557 4136
rect 530 3963 541 3966
rect 442 3923 445 3946
rect 490 3943 509 3946
rect 490 3933 493 3943
rect 450 3913 453 3926
rect 490 3893 493 3926
rect 378 3833 389 3836
rect 426 3883 433 3886
rect 426 3836 429 3883
rect 498 3856 501 3936
rect 506 3923 509 3943
rect 514 3933 517 3946
rect 522 3906 525 3926
rect 490 3853 501 3856
rect 514 3903 525 3906
rect 426 3833 437 3836
rect 354 3713 357 3726
rect 338 3673 357 3676
rect 354 3576 357 3673
rect 338 3573 357 3576
rect 338 3553 341 3573
rect 378 3556 381 3833
rect 386 3813 389 3826
rect 418 3793 421 3816
rect 426 3813 429 3826
rect 386 3723 389 3746
rect 394 3713 397 3726
rect 426 3706 429 3726
rect 418 3703 429 3706
rect 434 3706 437 3833
rect 442 3763 445 3826
rect 482 3813 485 3836
rect 482 3796 485 3806
rect 490 3803 493 3853
rect 498 3796 501 3816
rect 482 3793 501 3796
rect 506 3793 509 3806
rect 514 3766 517 3903
rect 498 3763 517 3766
rect 442 3743 461 3746
rect 442 3733 445 3743
rect 450 3723 453 3736
rect 458 3723 461 3743
rect 434 3703 445 3706
rect 418 3626 421 3703
rect 418 3623 429 3626
rect 370 3553 381 3556
rect 314 3523 325 3526
rect 330 3523 333 3536
rect 338 3513 341 3526
rect 370 3496 373 3553
rect 386 3543 405 3546
rect 386 3533 389 3543
rect 386 3503 389 3526
rect 394 3523 397 3536
rect 402 3523 405 3543
rect 410 3533 413 3546
rect 370 3493 381 3496
rect 286 3483 293 3486
rect 290 3463 293 3483
rect 242 3413 277 3416
rect 234 3383 237 3406
rect 250 3393 253 3406
rect 218 3353 229 3356
rect 218 3313 221 3353
rect 274 3346 277 3413
rect 290 3393 293 3406
rect 226 3343 245 3346
rect 226 3333 229 3343
rect 206 3303 213 3306
rect 210 3243 213 3303
rect 226 3256 229 3326
rect 218 3253 229 3256
rect 162 3213 165 3226
rect 162 3123 165 3146
rect 170 3133 173 3216
rect 178 3213 181 3236
rect 178 3123 181 3206
rect 186 3193 189 3206
rect 194 3203 197 3226
rect 218 3216 221 3253
rect 154 3103 165 3106
rect 162 3036 165 3103
rect 154 3033 165 3036
rect 186 3033 189 3186
rect 202 3166 205 3216
rect 210 3213 221 3216
rect 194 3163 205 3166
rect 194 3133 197 3163
rect 202 3133 205 3146
rect 210 3123 213 3196
rect 210 3086 213 3106
rect 202 3083 213 3086
rect 146 2993 149 3006
rect 138 2963 149 2966
rect 130 2733 133 2746
rect 138 2713 141 2726
rect 146 2603 149 2963
rect 154 2906 157 3033
rect 202 3026 205 3083
rect 202 3023 213 3026
rect 162 2923 165 3006
rect 170 2963 173 3016
rect 186 3003 189 3016
rect 194 2973 197 3006
rect 186 2933 189 2956
rect 210 2946 213 3023
rect 218 3013 221 3206
rect 226 3003 229 3246
rect 234 2983 237 3336
rect 242 3323 245 3343
rect 250 3333 253 3346
rect 274 3343 285 3346
rect 242 3296 245 3316
rect 242 3293 249 3296
rect 246 3226 249 3293
rect 242 3223 249 3226
rect 242 3103 245 3223
rect 258 3206 261 3326
rect 266 3233 269 3336
rect 266 3213 269 3226
rect 250 3193 253 3206
rect 258 3203 269 3206
rect 250 3113 253 3126
rect 258 3096 261 3146
rect 254 3093 261 3096
rect 254 3026 257 3093
rect 266 3053 269 3203
rect 274 3133 277 3216
rect 282 3153 285 3343
rect 306 3243 309 3326
rect 314 3323 317 3336
rect 306 3213 309 3226
rect 282 3066 285 3136
rect 290 3123 293 3196
rect 322 3176 325 3466
rect 378 3436 381 3493
rect 362 3433 381 3436
rect 338 3413 341 3426
rect 330 3333 333 3346
rect 298 3133 301 3176
rect 318 3173 325 3176
rect 306 3093 309 3126
rect 318 3106 321 3173
rect 330 3116 333 3156
rect 338 3123 341 3146
rect 346 3123 349 3156
rect 330 3113 341 3116
rect 318 3103 325 3106
rect 282 3063 293 3066
rect 242 3013 245 3026
rect 254 3023 261 3026
rect 250 2996 253 3006
rect 258 3003 261 3023
rect 266 3003 269 3016
rect 282 3013 285 3026
rect 250 2993 269 2996
rect 274 2993 277 3006
rect 290 3003 293 3063
rect 322 3056 325 3103
rect 298 2996 301 3056
rect 314 3053 325 3056
rect 338 3056 341 3113
rect 338 3053 349 3056
rect 314 3023 317 3053
rect 282 2993 301 2996
rect 210 2943 221 2946
rect 154 2903 165 2906
rect 162 2846 165 2903
rect 218 2896 221 2943
rect 250 2936 253 2956
rect 266 2936 269 2993
rect 250 2933 257 2936
rect 234 2903 237 2926
rect 154 2843 165 2846
rect 210 2893 221 2896
rect 154 2723 157 2843
rect 162 2743 165 2816
rect 178 2793 181 2806
rect 178 2723 181 2736
rect 186 2713 189 2736
rect 202 2723 205 2816
rect 210 2783 213 2893
rect 254 2886 257 2933
rect 266 2933 277 2936
rect 266 2923 269 2933
rect 282 2926 285 2993
rect 274 2923 285 2926
rect 250 2883 257 2886
rect 250 2826 253 2883
rect 246 2823 253 2826
rect 218 2683 221 2736
rect 234 2733 237 2756
rect 246 2746 249 2823
rect 246 2743 253 2746
rect 242 2713 245 2726
rect 162 2613 173 2616
rect 178 2613 181 2626
rect 154 2593 157 2606
rect 114 2566 117 2586
rect 114 2563 125 2566
rect 122 2516 125 2563
rect 162 2523 165 2606
rect 170 2596 173 2613
rect 170 2593 177 2596
rect 174 2526 177 2593
rect 170 2523 177 2526
rect 66 2503 85 2506
rect 114 2513 125 2516
rect 66 2476 69 2503
rect 66 2473 77 2476
rect 74 2396 77 2473
rect 114 2426 117 2513
rect 170 2506 173 2523
rect 162 2503 173 2506
rect 162 2436 165 2503
rect 162 2433 173 2436
rect 66 2393 77 2396
rect 106 2423 117 2426
rect 66 1933 69 2393
rect 106 2376 109 2423
rect 82 1993 85 2376
rect 106 2373 113 2376
rect 110 2316 113 2373
rect 122 2323 125 2416
rect 138 2403 141 2426
rect 170 2416 173 2433
rect 162 2413 173 2416
rect 178 2413 181 2426
rect 170 2406 173 2413
rect 162 2323 165 2406
rect 170 2403 181 2406
rect 186 2403 189 2606
rect 194 2583 197 2606
rect 250 2586 253 2743
rect 258 2733 261 2816
rect 266 2813 269 2906
rect 274 2836 277 2923
rect 274 2833 285 2836
rect 282 2796 285 2833
rect 290 2803 293 2926
rect 298 2883 301 2986
rect 314 2976 317 3016
rect 314 2973 325 2976
rect 306 2903 309 2966
rect 322 2856 325 2973
rect 338 2963 341 3006
rect 306 2853 325 2856
rect 306 2803 309 2853
rect 330 2796 333 2886
rect 274 2793 285 2796
rect 322 2793 333 2796
rect 274 2746 277 2793
rect 274 2743 285 2746
rect 282 2713 285 2743
rect 290 2693 293 2786
rect 298 2633 301 2736
rect 306 2656 309 2786
rect 314 2733 317 2746
rect 322 2733 325 2793
rect 346 2783 349 3053
rect 354 2953 357 3366
rect 362 3253 365 3433
rect 370 3333 373 3416
rect 378 3413 381 3426
rect 370 3306 373 3326
rect 370 3303 377 3306
rect 374 3246 377 3303
rect 370 3243 377 3246
rect 370 3173 373 3243
rect 362 3143 381 3146
rect 362 3123 365 3143
rect 370 3123 373 3136
rect 378 3133 381 3143
rect 362 3013 365 3026
rect 386 3013 389 3396
rect 394 3323 397 3406
rect 402 3243 405 3416
rect 410 3403 413 3526
rect 426 3523 429 3623
rect 442 3586 445 3703
rect 434 3583 445 3586
rect 434 3506 437 3583
rect 426 3503 437 3506
rect 426 3426 429 3503
rect 426 3423 437 3426
rect 410 3376 413 3396
rect 410 3373 417 3376
rect 414 3236 417 3373
rect 410 3233 417 3236
rect 402 3113 405 3176
rect 410 3116 413 3233
rect 418 3123 421 3216
rect 410 3113 417 3116
rect 394 3013 397 3056
rect 402 3013 405 3026
rect 414 2956 417 3113
rect 414 2953 421 2956
rect 370 2923 373 2936
rect 402 2923 405 2946
rect 410 2923 413 2936
rect 418 2906 421 2953
rect 410 2903 421 2906
rect 354 2813 357 2826
rect 386 2773 389 2816
rect 394 2813 397 2826
rect 394 2766 397 2806
rect 410 2796 413 2903
rect 410 2793 421 2796
rect 386 2763 397 2766
rect 322 2713 325 2726
rect 346 2723 349 2736
rect 306 2653 317 2656
rect 298 2613 301 2626
rect 226 2583 253 2586
rect 202 2493 205 2536
rect 210 2513 213 2526
rect 226 2483 229 2583
rect 314 2576 317 2653
rect 306 2573 317 2576
rect 250 2513 253 2526
rect 226 2413 229 2436
rect 242 2413 245 2496
rect 110 2313 117 2316
rect 114 2136 117 2313
rect 162 2296 165 2316
rect 154 2293 165 2296
rect 154 2236 157 2293
rect 154 2233 165 2236
rect 130 2213 133 2226
rect 162 2213 165 2233
rect 170 2223 173 2326
rect 178 2323 181 2403
rect 186 2343 205 2346
rect 186 2333 189 2343
rect 178 2203 181 2236
rect 186 2183 189 2326
rect 194 2313 197 2336
rect 202 2323 205 2343
rect 210 2303 213 2406
rect 234 2333 237 2406
rect 226 2253 229 2326
rect 242 2233 245 2326
rect 258 2323 261 2416
rect 282 2403 285 2416
rect 290 2386 293 2486
rect 298 2393 301 2406
rect 282 2383 293 2386
rect 306 2383 309 2573
rect 322 2556 325 2696
rect 318 2553 325 2556
rect 318 2436 321 2553
rect 330 2543 333 2616
rect 338 2613 341 2626
rect 318 2433 325 2436
rect 314 2393 317 2406
rect 258 2286 261 2306
rect 258 2283 265 2286
rect 202 2213 205 2226
rect 242 2213 245 2226
rect 218 2193 221 2206
rect 114 2133 125 2136
rect 106 2013 109 2126
rect 122 2006 125 2133
rect 194 2106 197 2126
rect 186 2103 197 2106
rect 186 2056 189 2103
rect 186 2053 197 2056
rect 162 2013 165 2026
rect 114 2003 125 2006
rect 82 1826 85 1936
rect 82 1823 93 1826
rect 82 1756 85 1806
rect 74 1753 85 1756
rect 74 1646 77 1753
rect 90 1656 93 1823
rect 98 1813 101 1986
rect 114 1956 117 2003
rect 110 1953 117 1956
rect 110 1896 113 1953
rect 122 1906 125 1946
rect 138 1923 141 1936
rect 154 1933 157 1996
rect 170 1983 173 2016
rect 178 1976 181 2036
rect 186 1993 189 2006
rect 178 1973 185 1976
rect 122 1903 133 1906
rect 110 1893 117 1896
rect 114 1816 117 1893
rect 110 1813 117 1816
rect 110 1756 113 1813
rect 130 1806 133 1903
rect 182 1896 185 1973
rect 194 1923 197 2053
rect 202 2003 205 2026
rect 210 2003 213 2186
rect 218 2013 221 2056
rect 226 2013 229 2136
rect 250 2123 253 2256
rect 262 2146 265 2283
rect 282 2266 285 2383
rect 298 2306 301 2336
rect 322 2323 325 2433
rect 330 2403 333 2526
rect 346 2386 349 2716
rect 362 2696 365 2756
rect 370 2713 373 2726
rect 386 2723 389 2763
rect 402 2733 405 2776
rect 402 2703 405 2726
rect 418 2713 421 2793
rect 362 2693 373 2696
rect 370 2646 373 2693
rect 426 2686 429 3406
rect 434 3393 437 3423
rect 434 3116 437 3336
rect 442 3323 445 3526
rect 458 3523 461 3566
rect 466 3513 469 3746
rect 490 3713 493 3736
rect 498 3706 501 3763
rect 514 3733 517 3756
rect 538 3746 541 3963
rect 554 3923 557 4096
rect 562 4023 565 4126
rect 570 4013 573 4136
rect 578 4113 581 4186
rect 586 4096 589 4136
rect 582 4093 589 4096
rect 582 4026 585 4093
rect 582 4023 589 4026
rect 562 3993 565 4006
rect 570 3816 573 3926
rect 578 3823 581 3936
rect 586 3923 589 4023
rect 594 3986 597 4416
rect 610 4413 613 4526
rect 634 4523 637 4583
rect 786 4556 789 4616
rect 810 4566 813 4606
rect 858 4603 861 4616
rect 778 4553 789 4556
rect 794 4563 813 4566
rect 650 4523 653 4536
rect 682 4533 685 4546
rect 626 4413 637 4416
rect 642 4413 645 4426
rect 602 4333 613 4336
rect 618 4333 621 4406
rect 650 4396 653 4486
rect 642 4393 653 4396
rect 610 4313 613 4326
rect 602 4213 605 4226
rect 618 4213 621 4326
rect 602 4133 605 4206
rect 602 4106 605 4126
rect 610 4123 613 4136
rect 618 4133 621 4206
rect 602 4103 609 4106
rect 606 4026 609 4103
rect 602 4023 609 4026
rect 602 4003 605 4023
rect 618 4013 621 4026
rect 594 3983 601 3986
rect 598 3916 601 3983
rect 594 3913 601 3916
rect 594 3816 597 3913
rect 570 3813 581 3816
rect 594 3813 601 3816
rect 538 3743 545 3746
rect 498 3703 517 3706
rect 482 3526 485 3656
rect 490 3533 493 3546
rect 474 3523 485 3526
rect 498 3523 501 3606
rect 450 3403 453 3446
rect 474 3413 477 3523
rect 490 3486 493 3516
rect 514 3503 517 3703
rect 542 3696 545 3743
rect 538 3693 545 3696
rect 522 3523 525 3546
rect 490 3483 501 3486
rect 498 3436 501 3483
rect 490 3433 501 3436
rect 490 3413 493 3433
rect 458 3403 469 3406
rect 482 3303 485 3336
rect 490 3323 493 3406
rect 506 3333 509 3346
rect 506 3313 509 3326
rect 466 3143 469 3216
rect 506 3203 509 3226
rect 434 3113 445 3116
rect 442 3006 445 3113
rect 458 3103 461 3126
rect 474 3036 477 3126
rect 482 3053 485 3136
rect 490 3113 493 3126
rect 434 3003 445 3006
rect 458 3033 477 3036
rect 458 3003 461 3033
rect 498 3013 501 3126
rect 506 3096 509 3116
rect 506 3093 513 3096
rect 510 3026 513 3093
rect 506 3023 513 3026
rect 506 3006 509 3023
rect 522 3006 525 3426
rect 530 3413 533 3436
rect 538 3273 541 3693
rect 554 3613 557 3726
rect 578 3676 581 3813
rect 586 3763 589 3806
rect 570 3673 581 3676
rect 570 3596 573 3673
rect 562 3593 573 3596
rect 562 3466 565 3593
rect 586 3576 589 3756
rect 598 3746 601 3813
rect 578 3573 589 3576
rect 594 3743 601 3746
rect 578 3486 581 3573
rect 594 3496 597 3743
rect 610 3736 613 3926
rect 618 3913 621 4006
rect 626 3846 629 4386
rect 642 4326 645 4393
rect 658 4333 661 4416
rect 690 4413 693 4536
rect 706 4533 717 4536
rect 722 4533 725 4546
rect 778 4543 781 4553
rect 698 4483 701 4526
rect 714 4513 717 4526
rect 754 4443 757 4536
rect 778 4513 781 4526
rect 794 4523 797 4563
rect 818 4513 821 4526
rect 642 4323 653 4326
rect 674 4323 677 4336
rect 754 4323 757 4416
rect 778 4336 781 4406
rect 794 4393 797 4406
rect 770 4333 781 4336
rect 650 4306 653 4323
rect 634 4093 637 4306
rect 650 4303 661 4306
rect 658 4226 661 4303
rect 770 4266 773 4333
rect 770 4263 781 4266
rect 650 4223 661 4226
rect 642 4193 645 4216
rect 650 4146 653 4223
rect 714 4216 717 4246
rect 666 4193 669 4206
rect 682 4146 685 4216
rect 698 4213 717 4216
rect 778 4213 781 4263
rect 786 4213 789 4326
rect 834 4323 837 4526
rect 874 4456 877 4526
rect 882 4523 885 4606
rect 906 4543 925 4546
rect 906 4533 909 4543
rect 890 4473 893 4526
rect 874 4453 893 4456
rect 858 4383 861 4416
rect 866 4413 869 4436
rect 882 4413 885 4446
rect 866 4336 869 4406
rect 874 4396 877 4406
rect 890 4403 893 4453
rect 898 4396 901 4406
rect 914 4403 917 4536
rect 922 4523 925 4543
rect 938 4533 941 4616
rect 1026 4613 1029 4626
rect 1018 4576 1021 4606
rect 1018 4573 1029 4576
rect 946 4533 949 4546
rect 938 4413 941 4526
rect 946 4403 949 4416
rect 874 4393 901 4396
rect 866 4333 873 4336
rect 690 4203 701 4206
rect 706 4193 709 4206
rect 714 4186 717 4213
rect 706 4183 717 4186
rect 646 4143 653 4146
rect 674 4143 685 4146
rect 646 4096 649 4143
rect 658 4103 661 4136
rect 674 4113 677 4143
rect 682 4133 693 4136
rect 698 4133 701 4146
rect 690 4116 693 4126
rect 706 4116 709 4183
rect 818 4163 821 4216
rect 834 4143 837 4156
rect 690 4113 709 4116
rect 646 4093 653 4096
rect 634 4003 637 4016
rect 642 4003 645 4016
rect 634 3923 637 3936
rect 642 3933 645 3986
rect 642 3903 645 3926
rect 622 3843 629 3846
rect 622 3796 625 3843
rect 634 3803 637 3836
rect 622 3793 629 3796
rect 642 3793 645 3806
rect 610 3733 617 3736
rect 602 3636 605 3726
rect 614 3676 617 3733
rect 610 3673 617 3676
rect 610 3653 613 3673
rect 626 3656 629 3793
rect 650 3753 653 4093
rect 658 3993 661 4006
rect 658 3943 677 3946
rect 658 3923 661 3943
rect 666 3923 669 3936
rect 674 3933 677 3943
rect 682 3926 685 4016
rect 682 3923 693 3926
rect 658 3896 661 3916
rect 658 3893 669 3896
rect 666 3836 669 3893
rect 658 3833 669 3836
rect 658 3736 661 3833
rect 666 3753 669 3816
rect 674 3793 677 3806
rect 642 3733 661 3736
rect 666 3743 685 3746
rect 666 3733 669 3743
rect 622 3653 629 3656
rect 602 3633 613 3636
rect 610 3566 613 3633
rect 602 3563 613 3566
rect 602 3533 605 3563
rect 622 3536 625 3653
rect 634 3563 637 3726
rect 642 3696 645 3733
rect 650 3723 661 3726
rect 666 3713 669 3726
rect 674 3723 677 3736
rect 682 3713 685 3743
rect 690 3723 693 3923
rect 642 3693 661 3696
rect 658 3556 661 3693
rect 706 3636 709 4113
rect 714 3983 717 4006
rect 730 4003 733 4126
rect 738 3913 741 3926
rect 746 3896 749 4116
rect 770 4086 773 4126
rect 762 4083 773 4086
rect 762 4013 765 4083
rect 754 4003 765 4006
rect 778 3966 781 4096
rect 818 4066 821 4136
rect 858 4093 861 4326
rect 870 4256 873 4333
rect 882 4313 885 4326
rect 898 4323 901 4393
rect 954 4386 957 4426
rect 946 4383 957 4386
rect 914 4323 917 4346
rect 922 4313 925 4326
rect 870 4253 893 4256
rect 890 4196 893 4253
rect 946 4246 949 4383
rect 962 4366 965 4536
rect 986 4523 989 4536
rect 1002 4523 1005 4546
rect 994 4496 997 4516
rect 986 4493 997 4496
rect 986 4426 989 4493
rect 1010 4453 1013 4536
rect 1026 4523 1029 4573
rect 1034 4533 1037 4616
rect 1066 4613 1069 4626
rect 1170 4623 1181 4626
rect 1114 4593 1117 4606
rect 1058 4533 1061 4556
rect 1082 4533 1085 4546
rect 1042 4513 1045 4526
rect 1058 4506 1061 4526
rect 1054 4503 1061 4506
rect 986 4423 997 4426
rect 970 4383 973 4406
rect 958 4363 965 4366
rect 958 4266 961 4363
rect 978 4353 981 4396
rect 994 4366 997 4423
rect 1002 4373 1005 4426
rect 1010 4386 1013 4406
rect 1026 4393 1029 4496
rect 1054 4436 1057 4503
rect 1054 4433 1061 4436
rect 1034 4413 1045 4416
rect 1010 4383 1017 4386
rect 994 4363 1005 4366
rect 970 4343 989 4346
rect 970 4333 973 4343
rect 958 4263 965 4266
rect 946 4243 957 4246
rect 906 4213 909 4226
rect 930 4213 941 4216
rect 946 4213 949 4226
rect 882 4193 893 4196
rect 882 4176 885 4193
rect 878 4173 885 4176
rect 866 4076 869 4136
rect 878 4116 881 4173
rect 890 4123 893 4146
rect 898 4123 901 4176
rect 878 4113 885 4116
rect 858 4073 869 4076
rect 818 4063 829 4066
rect 770 3963 781 3966
rect 754 3923 765 3926
rect 730 3893 749 3896
rect 730 3776 733 3893
rect 770 3886 773 3963
rect 810 3933 813 4016
rect 826 3976 829 4063
rect 826 3973 837 3976
rect 786 3913 789 3926
rect 770 3883 781 3886
rect 778 3826 781 3883
rect 778 3823 785 3826
rect 730 3773 749 3776
rect 738 3733 741 3756
rect 746 3736 749 3773
rect 746 3733 757 3736
rect 698 3633 709 3636
rect 618 3533 625 3536
rect 594 3493 601 3496
rect 578 3483 589 3486
rect 562 3463 581 3466
rect 578 3443 581 3463
rect 578 3413 581 3436
rect 554 3366 557 3406
rect 586 3373 589 3483
rect 598 3366 601 3493
rect 618 3456 621 3533
rect 634 3526 637 3556
rect 626 3523 637 3526
rect 642 3553 661 3556
rect 642 3523 645 3553
rect 682 3536 685 3576
rect 658 3533 693 3536
rect 634 3506 637 3523
rect 634 3503 645 3506
rect 618 3453 625 3456
rect 622 3366 625 3453
rect 642 3436 645 3503
rect 682 3453 685 3526
rect 634 3433 645 3436
rect 554 3363 565 3366
rect 562 3333 565 3363
rect 594 3363 601 3366
rect 546 3213 549 3236
rect 546 3123 549 3206
rect 554 3106 557 3246
rect 562 3213 565 3316
rect 570 3203 573 3216
rect 578 3213 581 3226
rect 586 3203 589 3306
rect 594 3153 597 3363
rect 602 3233 605 3326
rect 610 3216 613 3366
rect 622 3363 629 3366
rect 626 3276 629 3363
rect 602 3213 613 3216
rect 622 3273 629 3276
rect 602 3146 605 3213
rect 622 3206 625 3273
rect 434 2923 437 3003
rect 474 2953 477 3006
rect 498 3003 509 3006
rect 514 3003 525 3006
rect 546 3103 557 3106
rect 562 3143 581 3146
rect 546 3006 549 3103
rect 562 3013 565 3143
rect 570 3113 573 3136
rect 578 3133 581 3143
rect 586 3143 605 3146
rect 546 3003 557 3006
rect 466 2943 485 2946
rect 466 2933 469 2943
rect 466 2913 469 2926
rect 474 2923 477 2936
rect 482 2923 485 2943
rect 490 2933 493 2946
rect 498 2923 501 3003
rect 490 2813 493 2826
rect 514 2806 517 3003
rect 530 2883 533 2936
rect 538 2913 541 2926
rect 554 2896 557 3003
rect 546 2893 557 2896
rect 522 2813 525 2836
rect 530 2813 533 2826
rect 362 2643 373 2646
rect 418 2683 429 2686
rect 362 2623 365 2643
rect 362 2413 365 2536
rect 370 2523 373 2606
rect 330 2333 333 2346
rect 338 2323 341 2386
rect 346 2383 357 2386
rect 346 2313 349 2336
rect 354 2333 357 2383
rect 362 2373 365 2406
rect 362 2333 365 2366
rect 394 2363 397 2626
rect 418 2566 421 2683
rect 442 2573 445 2806
rect 514 2803 525 2806
rect 466 2613 469 2726
rect 474 2613 477 2716
rect 482 2596 485 2606
rect 490 2603 493 2626
rect 498 2596 501 2616
rect 506 2613 517 2616
rect 482 2593 501 2596
rect 418 2563 429 2566
rect 402 2483 405 2526
rect 426 2456 429 2563
rect 426 2453 433 2456
rect 410 2413 413 2426
rect 430 2376 433 2453
rect 482 2436 485 2576
rect 506 2513 509 2526
rect 482 2433 493 2436
rect 442 2383 445 2416
rect 450 2413 453 2426
rect 474 2403 477 2416
rect 482 2403 485 2426
rect 426 2373 433 2376
rect 386 2343 405 2346
rect 298 2303 309 2306
rect 282 2263 293 2266
rect 258 2143 265 2146
rect 234 2003 237 2016
rect 242 2013 245 2036
rect 242 1966 245 2006
rect 250 2003 253 2016
rect 258 2013 261 2143
rect 290 2133 293 2263
rect 306 2236 309 2303
rect 298 2233 309 2236
rect 298 2213 301 2233
rect 362 2226 365 2326
rect 378 2316 381 2336
rect 386 2323 389 2343
rect 394 2323 397 2336
rect 402 2333 405 2343
rect 378 2313 389 2316
rect 386 2236 389 2313
rect 410 2236 413 2336
rect 426 2246 429 2373
rect 442 2313 445 2326
rect 426 2243 437 2246
rect 386 2233 397 2236
rect 410 2233 421 2236
rect 354 2223 365 2226
rect 266 2096 269 2126
rect 266 2093 277 2096
rect 274 2036 277 2093
rect 266 2033 277 2036
rect 266 2013 269 2033
rect 274 1983 277 2016
rect 282 1973 285 2006
rect 234 1963 245 1966
rect 234 1923 237 1963
rect 266 1933 269 1946
rect 242 1906 245 1926
rect 178 1893 185 1896
rect 234 1903 245 1906
rect 178 1846 181 1893
rect 234 1846 237 1903
rect 250 1866 253 1926
rect 250 1863 261 1866
rect 178 1843 189 1846
rect 234 1843 245 1846
rect 122 1803 133 1806
rect 110 1753 117 1756
rect 90 1653 109 1656
rect 74 1643 85 1646
rect 82 1356 85 1643
rect 106 1436 109 1653
rect 114 1443 117 1753
rect 106 1433 117 1436
rect 66 1353 85 1356
rect 66 1296 69 1353
rect 66 1293 77 1296
rect 74 1076 77 1293
rect 90 1236 93 1376
rect 114 1346 117 1433
rect 122 1373 125 1803
rect 154 1793 157 1806
rect 130 1723 133 1786
rect 186 1776 189 1843
rect 202 1813 205 1826
rect 242 1823 245 1843
rect 234 1803 237 1816
rect 242 1813 253 1816
rect 258 1813 261 1863
rect 266 1806 269 1896
rect 290 1813 293 2126
rect 322 2123 325 2216
rect 354 2176 357 2223
rect 370 2176 373 2216
rect 386 2196 389 2206
rect 394 2203 397 2233
rect 402 2196 405 2216
rect 418 2213 421 2233
rect 386 2193 405 2196
rect 354 2173 365 2176
rect 370 2173 389 2176
rect 298 1923 301 2016
rect 306 2003 309 2016
rect 314 1996 317 2006
rect 322 2003 325 2016
rect 330 1996 333 2016
rect 354 2006 357 2016
rect 362 2013 365 2173
rect 386 2056 389 2173
rect 410 2133 413 2206
rect 370 2053 389 2056
rect 370 2033 373 2053
rect 314 1993 333 1996
rect 338 1983 341 2006
rect 346 2003 357 2006
rect 314 1956 317 1976
rect 310 1953 317 1956
rect 310 1886 313 1953
rect 310 1883 317 1886
rect 314 1826 317 1883
rect 338 1836 341 1966
rect 346 1923 349 2003
rect 354 1963 357 1996
rect 354 1903 357 1936
rect 362 1913 365 1926
rect 338 1833 349 1836
rect 314 1823 321 1826
rect 154 1773 189 1776
rect 154 1756 157 1773
rect 154 1753 165 1756
rect 162 1686 165 1753
rect 154 1683 165 1686
rect 154 1666 157 1683
rect 150 1663 157 1666
rect 130 1613 133 1626
rect 150 1606 153 1663
rect 178 1636 181 1736
rect 202 1723 205 1736
rect 210 1666 213 1746
rect 218 1733 237 1736
rect 242 1733 245 1806
rect 258 1803 269 1806
rect 249 1783 261 1786
rect 218 1673 221 1733
rect 162 1633 181 1636
rect 194 1663 213 1666
rect 162 1613 165 1633
rect 150 1603 157 1606
rect 130 1523 133 1536
rect 154 1483 157 1603
rect 170 1533 173 1616
rect 178 1613 181 1626
rect 130 1413 133 1426
rect 146 1403 149 1446
rect 162 1413 165 1436
rect 170 1413 173 1426
rect 178 1413 181 1596
rect 186 1576 189 1606
rect 194 1593 197 1663
rect 202 1613 205 1656
rect 186 1573 197 1576
rect 186 1533 189 1556
rect 194 1523 197 1573
rect 202 1506 205 1606
rect 218 1576 221 1666
rect 226 1653 229 1726
rect 234 1723 245 1726
rect 249 1723 252 1783
rect 258 1733 261 1776
rect 274 1743 277 1806
rect 258 1683 261 1726
rect 242 1603 245 1676
rect 274 1663 277 1736
rect 298 1733 301 1806
rect 306 1723 309 1816
rect 318 1746 321 1823
rect 330 1773 333 1816
rect 346 1813 349 1833
rect 378 1813 381 2006
rect 418 1973 421 2206
rect 434 2146 437 2243
rect 458 2233 461 2336
rect 482 2313 485 2326
rect 490 2236 493 2433
rect 514 2413 517 2426
rect 498 2383 501 2406
rect 466 2233 493 2236
rect 434 2143 445 2146
rect 450 2143 453 2216
rect 466 2176 469 2233
rect 474 2196 477 2216
rect 482 2203 485 2216
rect 490 2213 493 2226
rect 490 2196 493 2206
rect 474 2193 493 2196
rect 466 2173 485 2176
rect 426 2113 429 2126
rect 434 2103 437 2136
rect 442 2093 445 2143
rect 450 2023 453 2136
rect 458 2116 461 2136
rect 458 2113 469 2116
rect 466 2046 469 2113
rect 458 2043 469 2046
rect 458 1993 461 2043
rect 482 2026 485 2173
rect 506 2153 509 2376
rect 522 2276 525 2803
rect 546 2796 549 2893
rect 562 2803 565 2926
rect 570 2833 573 2936
rect 578 2923 581 3126
rect 586 3086 589 3143
rect 610 3133 613 3206
rect 622 3203 629 3206
rect 594 3113 597 3126
rect 610 3103 613 3126
rect 586 3083 597 3086
rect 594 2926 597 3083
rect 618 3013 621 3186
rect 626 3113 629 3203
rect 634 3096 637 3433
rect 642 3343 645 3416
rect 650 3413 661 3416
rect 658 3363 661 3413
rect 682 3403 685 3426
rect 674 3386 677 3396
rect 690 3386 693 3406
rect 666 3383 677 3386
rect 686 3383 693 3386
rect 658 3333 661 3346
rect 642 3306 645 3326
rect 642 3303 649 3306
rect 646 3236 649 3303
rect 642 3233 649 3236
rect 642 3203 645 3233
rect 658 3213 661 3276
rect 666 3173 669 3206
rect 630 3093 637 3096
rect 642 3096 645 3156
rect 674 3153 677 3376
rect 686 3226 689 3383
rect 686 3223 693 3226
rect 682 3143 685 3206
rect 658 3103 661 3136
rect 690 3126 693 3223
rect 686 3123 693 3126
rect 642 3093 649 3096
rect 630 2976 633 3093
rect 646 3046 649 3093
rect 646 3043 669 3046
rect 630 2973 637 2976
rect 626 2936 629 2956
rect 586 2923 597 2926
rect 618 2933 629 2936
rect 578 2813 581 2826
rect 546 2793 557 2796
rect 554 2736 557 2793
rect 554 2733 565 2736
rect 538 2603 541 2726
rect 562 2656 565 2733
rect 554 2653 565 2656
rect 554 2636 557 2653
rect 586 2636 589 2923
rect 602 2856 605 2906
rect 618 2876 621 2933
rect 618 2873 629 2876
rect 598 2853 605 2856
rect 626 2853 629 2873
rect 598 2776 601 2853
rect 634 2826 637 2973
rect 642 2923 645 3016
rect 658 2983 661 3006
rect 666 2976 669 3043
rect 674 3003 677 3056
rect 658 2973 669 2976
rect 650 2933 653 2956
rect 658 2923 661 2973
rect 686 2946 689 3123
rect 698 2956 701 3633
rect 706 3533 709 3546
rect 706 3323 709 3446
rect 714 3423 717 3616
rect 738 3613 741 3726
rect 714 3333 717 3366
rect 722 3303 725 3436
rect 730 3383 733 3456
rect 738 3413 741 3526
rect 730 3333 733 3356
rect 706 3213 709 3256
rect 754 3216 757 3733
rect 770 3723 773 3816
rect 782 3766 785 3823
rect 810 3783 813 3836
rect 834 3833 837 3973
rect 850 3923 853 3936
rect 826 3793 829 3816
rect 778 3763 785 3766
rect 778 3723 781 3763
rect 794 3723 797 3736
rect 778 3533 789 3536
rect 794 3533 797 3716
rect 818 3696 821 3726
rect 834 3703 837 3726
rect 810 3693 821 3696
rect 810 3603 813 3693
rect 842 3626 845 3796
rect 858 3766 861 4073
rect 874 4003 877 4016
rect 866 3983 869 3996
rect 882 3843 885 4113
rect 914 4106 917 4136
rect 922 4123 925 4196
rect 930 4133 933 4213
rect 946 4193 949 4206
rect 954 4146 957 4243
rect 962 4153 965 4263
rect 970 4233 973 4326
rect 978 4323 981 4336
rect 986 4323 989 4343
rect 994 4333 997 4346
rect 1002 4323 1005 4363
rect 1014 4326 1017 4383
rect 1010 4323 1017 4326
rect 1010 4306 1013 4323
rect 1002 4303 1013 4306
rect 1002 4226 1005 4303
rect 1002 4223 1013 4226
rect 970 4193 973 4206
rect 954 4143 973 4146
rect 962 4106 965 4126
rect 914 4103 925 4106
rect 890 3903 893 3926
rect 882 3803 885 3836
rect 858 3763 865 3766
rect 862 3686 865 3763
rect 874 3723 877 3756
rect 890 3733 893 3816
rect 858 3683 865 3686
rect 842 3623 849 3626
rect 770 3433 773 3526
rect 794 3443 797 3526
rect 834 3523 837 3616
rect 846 3516 849 3623
rect 842 3513 849 3516
rect 842 3456 845 3513
rect 858 3506 861 3683
rect 882 3626 885 3716
rect 890 3703 893 3726
rect 878 3623 885 3626
rect 878 3546 881 3623
rect 866 3533 869 3546
rect 878 3543 885 3546
rect 882 3523 885 3543
rect 890 3533 893 3616
rect 898 3586 901 4046
rect 906 3913 909 3936
rect 914 3896 917 4006
rect 922 3916 925 4103
rect 954 4103 965 4106
rect 954 4026 957 4103
rect 970 4043 973 4143
rect 986 4036 989 4206
rect 954 4023 965 4026
rect 922 3913 933 3916
rect 946 3913 949 3926
rect 910 3893 917 3896
rect 910 3826 913 3893
rect 930 3866 933 3913
rect 922 3863 933 3866
rect 922 3833 925 3863
rect 938 3826 941 3846
rect 910 3823 917 3826
rect 906 3753 909 3806
rect 914 3626 917 3823
rect 934 3823 941 3826
rect 922 3793 925 3816
rect 922 3743 925 3776
rect 934 3726 937 3823
rect 930 3723 937 3726
rect 930 3646 933 3723
rect 930 3643 941 3646
rect 906 3623 917 3626
rect 906 3606 909 3623
rect 922 3616 925 3626
rect 914 3613 925 3616
rect 906 3603 917 3606
rect 898 3583 905 3586
rect 902 3526 905 3583
rect 898 3523 905 3526
rect 898 3506 901 3523
rect 858 3503 869 3506
rect 842 3453 849 3456
rect 746 3213 757 3216
rect 706 3013 709 3126
rect 722 3086 725 3166
rect 746 3126 749 3213
rect 770 3133 773 3206
rect 778 3163 781 3406
rect 786 3306 789 3336
rect 810 3323 813 3416
rect 846 3376 849 3453
rect 866 3426 869 3503
rect 842 3373 849 3376
rect 858 3423 869 3426
rect 890 3503 901 3506
rect 786 3303 797 3306
rect 794 3236 797 3303
rect 786 3233 797 3236
rect 786 3213 789 3233
rect 818 3193 821 3326
rect 842 3226 845 3373
rect 858 3356 861 3423
rect 874 3393 877 3406
rect 890 3376 893 3503
rect 914 3426 917 3603
rect 930 3543 933 3616
rect 922 3523 925 3536
rect 938 3506 941 3643
rect 946 3623 949 3836
rect 954 3813 957 4006
rect 962 3833 965 4023
rect 970 4013 973 4036
rect 986 4033 997 4036
rect 978 4003 981 4026
rect 994 3966 997 4033
rect 986 3963 997 3966
rect 978 3936 981 3956
rect 974 3933 981 3936
rect 974 3846 977 3933
rect 974 3843 981 3846
rect 970 3793 973 3826
rect 930 3503 941 3506
rect 930 3446 933 3503
rect 930 3443 937 3446
rect 914 3423 925 3426
rect 890 3373 901 3376
rect 854 3353 861 3356
rect 854 3306 857 3353
rect 854 3303 861 3306
rect 838 3223 845 3226
rect 746 3123 757 3126
rect 778 3123 781 3146
rect 810 3133 813 3146
rect 722 3083 733 3086
rect 730 3006 733 3083
rect 722 3003 733 3006
rect 698 2953 705 2956
rect 666 2933 669 2946
rect 686 2943 693 2946
rect 682 2906 685 2926
rect 674 2903 685 2906
rect 674 2846 677 2903
rect 674 2843 685 2846
rect 630 2823 637 2826
rect 598 2773 605 2776
rect 550 2633 557 2636
rect 578 2633 589 2636
rect 550 2516 553 2633
rect 562 2523 565 2606
rect 570 2533 573 2616
rect 578 2613 581 2633
rect 550 2513 557 2516
rect 570 2513 573 2526
rect 538 2413 541 2486
rect 530 2393 541 2396
rect 546 2373 549 2406
rect 554 2366 557 2513
rect 546 2363 557 2366
rect 518 2273 525 2276
rect 530 2323 541 2326
rect 518 2186 521 2273
rect 518 2183 525 2186
rect 514 2136 517 2166
rect 466 2023 485 2026
rect 506 2133 517 2136
rect 466 2003 469 2023
rect 402 1913 405 1926
rect 338 1793 341 1806
rect 314 1743 321 1746
rect 314 1683 317 1743
rect 322 1713 325 1726
rect 354 1723 357 1746
rect 362 1713 365 1726
rect 370 1693 373 1806
rect 378 1726 381 1806
rect 386 1803 389 1816
rect 394 1803 397 1876
rect 402 1813 405 1906
rect 386 1743 405 1746
rect 386 1733 389 1743
rect 394 1726 397 1736
rect 378 1723 397 1726
rect 402 1723 405 1743
rect 410 1733 413 1746
rect 266 1613 269 1626
rect 298 1593 301 1616
rect 306 1613 309 1626
rect 330 1613 333 1686
rect 338 1613 357 1616
rect 218 1573 229 1576
rect 210 1513 213 1526
rect 202 1503 217 1506
rect 214 1436 217 1503
rect 114 1343 125 1346
rect 122 1296 125 1343
rect 138 1313 141 1326
rect 162 1316 165 1406
rect 186 1346 189 1416
rect 194 1396 197 1406
rect 202 1403 205 1436
rect 214 1433 221 1436
rect 210 1396 213 1416
rect 194 1393 213 1396
rect 186 1343 197 1346
rect 170 1323 173 1336
rect 162 1313 173 1316
rect 178 1313 181 1326
rect 86 1233 93 1236
rect 106 1293 125 1296
rect 86 1186 89 1233
rect 106 1203 109 1293
rect 170 1256 173 1313
rect 170 1253 177 1256
rect 86 1183 93 1186
rect 66 1073 77 1076
rect 66 973 69 1073
rect 90 1056 93 1183
rect 98 1113 101 1136
rect 106 1106 109 1126
rect 146 1123 149 1216
rect 174 1176 177 1253
rect 194 1246 197 1343
rect 170 1173 177 1176
rect 186 1243 197 1246
rect 170 1106 173 1173
rect 186 1106 189 1243
rect 218 1216 221 1433
rect 226 1363 229 1573
rect 274 1513 277 1526
rect 306 1523 309 1546
rect 314 1513 317 1526
rect 322 1523 325 1536
rect 234 1336 237 1486
rect 242 1386 245 1406
rect 242 1383 249 1386
rect 230 1333 237 1336
rect 230 1236 233 1333
rect 246 1326 249 1383
rect 242 1323 249 1326
rect 230 1233 237 1236
rect 194 1123 197 1216
rect 218 1213 229 1216
rect 202 1143 221 1146
rect 202 1133 205 1143
rect 210 1123 213 1136
rect 218 1123 221 1143
rect 106 1103 117 1106
rect 82 1053 93 1056
rect 82 956 85 1053
rect 114 1036 117 1103
rect 162 1103 173 1106
rect 162 1046 165 1103
rect 162 1043 173 1046
rect 106 1033 117 1036
rect 106 1013 109 1033
rect 74 953 85 956
rect 74 836 77 953
rect 90 856 93 976
rect 170 966 173 1043
rect 178 973 181 1106
rect 186 1103 197 1106
rect 194 1036 197 1103
rect 186 1033 197 1036
rect 170 963 181 966
rect 186 963 189 1033
rect 194 1003 197 1016
rect 210 1013 213 1116
rect 226 1103 229 1213
rect 234 1133 237 1233
rect 242 1116 245 1323
rect 250 1133 253 1216
rect 258 1143 261 1366
rect 266 1303 269 1416
rect 274 1403 277 1506
rect 338 1503 341 1613
rect 346 1596 349 1606
rect 354 1603 357 1613
rect 362 1596 365 1616
rect 346 1593 365 1596
rect 370 1593 373 1606
rect 378 1596 381 1626
rect 386 1603 389 1636
rect 394 1613 397 1723
rect 418 1706 421 1816
rect 434 1803 437 1856
rect 458 1853 461 1926
rect 466 1893 469 1936
rect 498 1933 501 1956
rect 490 1856 493 1926
rect 506 1906 509 2133
rect 522 2113 525 2183
rect 530 2133 533 2323
rect 546 2236 549 2363
rect 562 2303 565 2416
rect 542 2233 549 2236
rect 542 2186 545 2233
rect 554 2213 557 2226
rect 562 2213 573 2216
rect 542 2183 549 2186
rect 546 2163 549 2183
rect 514 2003 517 2016
rect 522 2013 525 2036
rect 530 2016 533 2126
rect 538 2023 541 2136
rect 546 2096 549 2126
rect 554 2123 557 2156
rect 570 2133 573 2213
rect 578 2136 581 2596
rect 586 2523 589 2616
rect 594 2593 597 2636
rect 602 2436 605 2773
rect 610 2603 613 2626
rect 610 2533 613 2546
rect 594 2433 605 2436
rect 594 2266 597 2433
rect 610 2413 613 2426
rect 618 2413 621 2786
rect 630 2736 633 2823
rect 642 2743 645 2816
rect 666 2803 669 2816
rect 630 2733 637 2736
rect 650 2733 653 2766
rect 666 2733 669 2756
rect 634 2606 637 2733
rect 658 2673 661 2726
rect 674 2723 677 2746
rect 682 2656 685 2843
rect 690 2833 693 2943
rect 702 2896 705 2953
rect 722 2923 725 3003
rect 702 2893 709 2896
rect 706 2836 709 2893
rect 698 2833 709 2836
rect 690 2723 693 2826
rect 698 2716 701 2833
rect 706 2746 709 2816
rect 722 2756 725 2836
rect 722 2753 729 2756
rect 706 2743 717 2746
rect 630 2603 637 2606
rect 674 2653 685 2656
rect 690 2713 701 2716
rect 714 2713 717 2743
rect 690 2656 693 2713
rect 726 2706 729 2753
rect 722 2703 729 2706
rect 690 2653 701 2656
rect 630 2436 633 2603
rect 630 2433 637 2436
rect 610 2373 613 2406
rect 626 2403 629 2416
rect 594 2263 605 2266
rect 594 2213 597 2226
rect 578 2133 585 2136
rect 546 2093 557 2096
rect 554 2016 557 2093
rect 530 2013 541 2016
rect 554 2013 565 2016
rect 546 1993 549 2006
rect 514 1913 517 1936
rect 506 1903 517 1906
rect 490 1853 501 1856
rect 450 1736 453 1826
rect 442 1733 453 1736
rect 466 1733 469 1776
rect 474 1733 485 1736
rect 410 1703 421 1706
rect 410 1646 413 1703
rect 410 1643 421 1646
rect 418 1623 421 1643
rect 378 1593 397 1596
rect 354 1543 373 1546
rect 354 1533 357 1543
rect 354 1513 357 1526
rect 362 1523 365 1536
rect 370 1523 373 1543
rect 378 1533 381 1546
rect 386 1533 389 1556
rect 394 1526 397 1593
rect 402 1583 405 1616
rect 426 1613 429 1726
rect 410 1563 413 1606
rect 426 1593 429 1606
rect 386 1523 397 1526
rect 314 1436 317 1456
rect 282 1343 285 1416
rect 290 1333 293 1406
rect 298 1316 301 1416
rect 306 1333 309 1436
rect 314 1433 325 1436
rect 322 1376 325 1433
rect 386 1426 389 1523
rect 370 1423 389 1426
rect 370 1413 373 1423
rect 314 1373 325 1376
rect 290 1313 301 1316
rect 290 1256 293 1313
rect 314 1256 317 1373
rect 322 1333 325 1356
rect 330 1333 341 1336
rect 338 1313 341 1326
rect 290 1253 301 1256
rect 266 1136 269 1236
rect 298 1233 301 1253
rect 306 1253 317 1256
rect 258 1133 269 1136
rect 234 1113 245 1116
rect 226 1013 229 1026
rect 202 993 205 1006
rect 218 983 221 1006
rect 178 936 181 963
rect 138 913 141 926
rect 170 923 173 936
rect 178 933 189 936
rect 178 913 181 926
rect 186 903 189 933
rect 194 913 197 936
rect 90 853 109 856
rect 74 833 85 836
rect 82 756 85 833
rect 106 776 109 853
rect 130 813 133 826
rect 162 793 165 816
rect 170 813 173 826
rect 202 803 205 826
rect 210 786 213 976
rect 226 936 229 1006
rect 234 983 237 1113
rect 218 933 229 936
rect 218 913 221 926
rect 234 846 237 966
rect 218 843 237 846
rect 218 813 221 843
rect 234 833 237 843
rect 242 836 245 1026
rect 250 1013 253 1036
rect 258 1023 261 1133
rect 266 1113 269 1126
rect 274 1123 277 1206
rect 282 1196 285 1216
rect 306 1213 309 1253
rect 354 1213 357 1336
rect 378 1323 381 1416
rect 402 1386 405 1406
rect 418 1403 421 1466
rect 426 1453 429 1586
rect 442 1573 445 1733
rect 474 1723 485 1726
rect 490 1723 493 1816
rect 498 1723 501 1853
rect 434 1443 437 1536
rect 450 1533 453 1546
rect 442 1506 445 1526
rect 442 1503 449 1506
rect 446 1406 449 1503
rect 442 1403 449 1406
rect 394 1383 405 1386
rect 394 1286 397 1383
rect 394 1283 405 1286
rect 370 1213 373 1226
rect 402 1213 405 1283
rect 282 1193 289 1196
rect 286 1126 289 1193
rect 298 1173 301 1206
rect 314 1183 317 1206
rect 282 1123 289 1126
rect 282 1013 285 1123
rect 306 1113 309 1126
rect 250 846 253 986
rect 258 973 261 1006
rect 274 993 277 1006
rect 298 966 301 1056
rect 354 1053 357 1146
rect 394 1133 397 1206
rect 410 1193 413 1206
rect 418 1026 421 1206
rect 434 1133 437 1326
rect 442 1313 445 1403
rect 458 1156 461 1596
rect 474 1583 477 1723
rect 490 1613 493 1626
rect 514 1593 517 1903
rect 522 1823 525 1936
rect 530 1903 533 1926
rect 554 1923 557 2006
rect 570 2003 573 2126
rect 582 2036 585 2133
rect 582 2033 589 2036
rect 578 1933 581 2016
rect 586 2003 589 2033
rect 594 1966 597 2166
rect 602 1986 605 2263
rect 610 2163 613 2366
rect 634 2363 637 2433
rect 642 2386 645 2596
rect 674 2576 677 2653
rect 674 2573 685 2576
rect 666 2536 669 2546
rect 658 2533 669 2536
rect 674 2533 677 2556
rect 666 2466 669 2526
rect 658 2463 669 2466
rect 650 2403 653 2446
rect 658 2413 661 2463
rect 666 2393 669 2406
rect 642 2383 649 2386
rect 626 2343 637 2346
rect 634 2313 637 2326
rect 646 2306 649 2383
rect 682 2376 685 2573
rect 698 2546 701 2653
rect 690 2543 701 2546
rect 690 2513 693 2543
rect 722 2536 725 2703
rect 738 2613 741 2806
rect 754 2783 757 3123
rect 786 3043 789 3126
rect 794 3006 797 3026
rect 802 3013 805 3126
rect 826 3023 829 3216
rect 810 3013 829 3016
rect 790 3003 797 3006
rect 810 3003 813 3013
rect 770 2973 773 2996
rect 770 2923 773 2936
rect 790 2896 793 3003
rect 818 2986 821 3006
rect 802 2983 821 2986
rect 790 2893 797 2896
rect 770 2756 773 2816
rect 794 2813 797 2893
rect 802 2803 805 2983
rect 826 2946 829 3013
rect 838 2956 841 3223
rect 838 2953 845 2956
rect 822 2943 829 2946
rect 810 2923 813 2936
rect 810 2823 813 2886
rect 822 2806 825 2943
rect 834 2813 837 2936
rect 842 2806 845 2953
rect 850 2823 853 3216
rect 858 3166 861 3303
rect 874 3226 877 3336
rect 898 3293 901 3373
rect 874 3223 901 3226
rect 882 3213 893 3216
rect 866 3186 869 3206
rect 890 3186 893 3206
rect 866 3183 893 3186
rect 858 3163 869 3166
rect 866 3046 869 3163
rect 862 3043 869 3046
rect 862 2976 865 3043
rect 874 3013 877 3026
rect 882 3013 885 3166
rect 898 2976 901 3223
rect 906 3203 909 3416
rect 922 3376 925 3423
rect 914 3373 925 3376
rect 934 3376 937 3443
rect 934 3373 941 3376
rect 946 3373 949 3596
rect 954 3496 957 3736
rect 962 3723 965 3746
rect 970 3733 973 3756
rect 970 3713 973 3726
rect 962 3613 965 3676
rect 978 3633 981 3843
rect 970 3583 973 3606
rect 978 3533 981 3616
rect 986 3593 989 3963
rect 1010 3953 1013 4223
rect 1026 4213 1029 4326
rect 1034 4203 1037 4216
rect 1018 4133 1021 4146
rect 1026 4133 1029 4146
rect 1034 4063 1037 4116
rect 1042 4026 1045 4406
rect 1050 4403 1053 4416
rect 1058 4403 1061 4433
rect 1066 4413 1069 4526
rect 1082 4463 1085 4526
rect 1090 4523 1093 4536
rect 1162 4533 1165 4616
rect 1178 4556 1181 4623
rect 1170 4553 1181 4556
rect 1114 4513 1117 4526
rect 1138 4513 1141 4526
rect 1090 4423 1093 4476
rect 1074 4403 1085 4406
rect 1090 4403 1093 4416
rect 1098 4383 1101 4426
rect 1106 4413 1109 4436
rect 1114 4413 1117 4426
rect 1154 4416 1157 4526
rect 1162 4493 1165 4526
rect 1170 4523 1173 4553
rect 1186 4526 1189 4536
rect 1178 4523 1189 4526
rect 1154 4413 1165 4416
rect 1178 4413 1181 4523
rect 1186 4496 1189 4516
rect 1194 4513 1197 4536
rect 1210 4523 1213 4536
rect 1226 4523 1229 4616
rect 1258 4526 1261 4606
rect 1266 4533 1269 4556
rect 1250 4523 1261 4526
rect 1186 4493 1197 4496
rect 1194 4436 1197 4493
rect 1186 4433 1197 4436
rect 1186 4413 1189 4433
rect 1058 4296 1061 4326
rect 1074 4323 1077 4336
rect 1082 4313 1085 4346
rect 1090 4333 1093 4366
rect 1106 4343 1125 4346
rect 1058 4293 1069 4296
rect 1066 4236 1069 4293
rect 1058 4233 1069 4236
rect 1098 4236 1101 4336
rect 1106 4323 1109 4343
rect 1114 4303 1117 4336
rect 1122 4333 1125 4343
rect 1130 4303 1133 4406
rect 1138 4393 1141 4406
rect 1098 4233 1117 4236
rect 1058 4216 1061 4233
rect 1058 4213 1069 4216
rect 1066 4156 1069 4213
rect 1066 4153 1077 4156
rect 1050 4116 1053 4136
rect 1050 4113 1061 4116
rect 1058 4046 1061 4113
rect 1074 4083 1077 4153
rect 1082 4133 1085 4206
rect 1090 4183 1093 4216
rect 1098 4193 1101 4226
rect 1106 4213 1109 4226
rect 1098 4136 1101 4156
rect 1026 4023 1045 4026
rect 1050 4043 1061 4046
rect 1026 3953 1029 4023
rect 1034 4013 1045 4016
rect 994 3896 997 3946
rect 994 3893 1001 3896
rect 998 3836 1001 3893
rect 1010 3863 1013 3936
rect 1034 3923 1037 4006
rect 1042 3983 1045 4006
rect 1050 3996 1053 4043
rect 1058 4013 1061 4026
rect 1050 3993 1057 3996
rect 1074 3993 1077 4016
rect 1082 4013 1085 4056
rect 994 3833 1001 3836
rect 994 3813 997 3833
rect 994 3716 997 3806
rect 1002 3763 1013 3766
rect 1002 3733 1005 3746
rect 1010 3743 1013 3763
rect 994 3713 1001 3716
rect 998 3636 1001 3713
rect 994 3633 1001 3636
rect 994 3543 997 3633
rect 962 3513 965 3526
rect 1002 3523 1005 3616
rect 954 3493 965 3496
rect 962 3426 965 3493
rect 1010 3476 1013 3636
rect 1018 3613 1021 3646
rect 954 3423 965 3426
rect 1002 3473 1013 3476
rect 914 3186 917 3373
rect 922 3313 925 3326
rect 910 3183 917 3186
rect 910 3106 913 3183
rect 922 3163 925 3296
rect 922 3113 925 3126
rect 910 3103 917 3106
rect 906 3003 909 3026
rect 858 2973 865 2976
rect 874 2973 901 2976
rect 818 2803 825 2806
rect 834 2803 845 2806
rect 754 2753 773 2756
rect 746 2596 749 2676
rect 742 2593 749 2596
rect 722 2533 733 2536
rect 714 2506 717 2526
rect 706 2503 717 2506
rect 706 2456 709 2503
rect 730 2466 733 2533
rect 742 2516 745 2593
rect 754 2523 757 2753
rect 762 2743 781 2746
rect 762 2733 765 2743
rect 770 2723 773 2736
rect 778 2723 781 2743
rect 742 2513 749 2516
rect 726 2463 733 2466
rect 706 2453 717 2456
rect 714 2413 717 2453
rect 726 2406 729 2463
rect 746 2456 749 2513
rect 746 2453 753 2456
rect 722 2403 729 2406
rect 682 2373 693 2376
rect 642 2303 649 2306
rect 610 2046 613 2136
rect 618 2133 621 2236
rect 642 2213 645 2303
rect 642 2193 645 2206
rect 658 2176 661 2356
rect 650 2173 661 2176
rect 610 2043 621 2046
rect 610 2003 613 2036
rect 602 1983 609 1986
rect 586 1963 597 1966
rect 562 1873 565 1926
rect 578 1913 581 1926
rect 586 1873 589 1963
rect 594 1943 597 1956
rect 606 1916 609 1983
rect 618 1933 621 2043
rect 634 1916 637 2156
rect 650 1936 653 2173
rect 666 2156 669 2336
rect 674 2323 677 2346
rect 674 2286 677 2306
rect 674 2283 681 2286
rect 678 2176 681 2283
rect 690 2223 693 2373
rect 722 2336 725 2403
rect 750 2396 753 2453
rect 762 2406 765 2416
rect 770 2413 773 2716
rect 794 2683 797 2756
rect 818 2736 821 2803
rect 802 2716 805 2736
rect 818 2733 829 2736
rect 802 2713 813 2716
rect 810 2636 813 2713
rect 794 2633 813 2636
rect 786 2603 789 2626
rect 762 2403 773 2406
rect 746 2393 753 2396
rect 746 2376 749 2393
rect 738 2373 749 2376
rect 722 2333 729 2336
rect 714 2213 717 2326
rect 726 2216 729 2333
rect 722 2213 729 2216
rect 690 2193 693 2206
rect 722 2196 725 2213
rect 714 2193 725 2196
rect 662 2153 669 2156
rect 674 2173 681 2176
rect 674 2153 677 2173
rect 662 2036 665 2153
rect 674 2123 677 2146
rect 714 2136 717 2193
rect 738 2146 741 2373
rect 786 2306 789 2326
rect 778 2303 789 2306
rect 778 2246 781 2303
rect 794 2283 797 2633
rect 826 2613 829 2733
rect 834 2716 837 2803
rect 850 2733 853 2806
rect 834 2713 845 2716
rect 842 2626 845 2713
rect 838 2623 845 2626
rect 802 2543 821 2546
rect 802 2533 805 2543
rect 810 2403 813 2536
rect 818 2523 821 2543
rect 826 2533 829 2576
rect 838 2546 841 2623
rect 834 2543 841 2546
rect 834 2433 837 2543
rect 850 2526 853 2606
rect 858 2596 861 2973
rect 874 2956 877 2973
rect 866 2943 869 2956
rect 874 2953 893 2956
rect 866 2813 869 2906
rect 890 2846 893 2953
rect 874 2843 893 2846
rect 874 2723 877 2843
rect 914 2826 917 3103
rect 938 3036 941 3373
rect 954 3336 957 3423
rect 978 3346 981 3406
rect 1002 3346 1005 3473
rect 1018 3456 1021 3546
rect 1014 3453 1021 3456
rect 1026 3453 1029 3806
rect 1034 3803 1037 3816
rect 1034 3693 1037 3716
rect 1034 3603 1037 3626
rect 1014 3396 1017 3453
rect 1026 3403 1029 3416
rect 1034 3403 1037 3476
rect 1014 3393 1021 3396
rect 978 3343 985 3346
rect 1002 3343 1009 3346
rect 954 3333 973 3336
rect 946 3323 957 3326
rect 962 3313 965 3326
rect 970 3306 973 3333
rect 954 3303 973 3306
rect 946 3103 949 3116
rect 934 3033 941 3036
rect 922 2993 925 3006
rect 934 2976 937 3033
rect 946 3013 949 3026
rect 930 2973 937 2976
rect 930 2846 933 2973
rect 930 2843 937 2846
rect 866 2613 869 2636
rect 882 2613 885 2686
rect 890 2613 893 2626
rect 858 2593 865 2596
rect 846 2523 853 2526
rect 846 2446 849 2523
rect 862 2516 865 2593
rect 858 2513 865 2516
rect 858 2456 861 2513
rect 858 2453 865 2456
rect 846 2443 853 2446
rect 818 2413 829 2416
rect 826 2396 829 2413
rect 842 2403 845 2426
rect 826 2393 837 2396
rect 802 2366 805 2386
rect 802 2363 813 2366
rect 810 2306 813 2363
rect 834 2323 837 2393
rect 850 2353 853 2443
rect 862 2396 865 2453
rect 858 2393 865 2396
rect 850 2333 853 2346
rect 858 2306 861 2393
rect 874 2383 877 2606
rect 882 2593 885 2606
rect 866 2323 869 2376
rect 874 2306 877 2336
rect 802 2303 813 2306
rect 850 2303 861 2306
rect 870 2303 877 2306
rect 778 2243 789 2246
rect 754 2156 757 2216
rect 754 2153 761 2156
rect 738 2143 749 2146
rect 706 2133 717 2136
rect 730 2133 741 2136
rect 662 2033 669 2036
rect 674 2033 677 2116
rect 706 2066 709 2133
rect 722 2076 725 2126
rect 730 2123 733 2133
rect 746 2116 749 2143
rect 742 2113 749 2116
rect 722 2073 733 2076
rect 706 2063 717 2066
rect 666 2013 669 2033
rect 690 2016 693 2046
rect 682 2013 693 2016
rect 714 2013 717 2063
rect 730 2026 733 2073
rect 722 2023 733 2026
rect 650 1933 657 1936
rect 666 1933 669 2006
rect 606 1913 613 1916
rect 610 1866 613 1913
rect 602 1863 613 1866
rect 626 1913 637 1916
rect 602 1826 605 1863
rect 602 1823 613 1826
rect 538 1723 541 1806
rect 554 1713 557 1736
rect 522 1603 525 1616
rect 530 1613 533 1626
rect 538 1613 541 1646
rect 474 1463 477 1576
rect 554 1546 557 1696
rect 562 1673 565 1726
rect 570 1696 573 1806
rect 594 1733 597 1816
rect 610 1756 613 1823
rect 602 1753 613 1756
rect 578 1713 581 1726
rect 602 1716 605 1753
rect 626 1746 629 1913
rect 642 1763 645 1916
rect 654 1846 657 1933
rect 690 1913 693 1926
rect 654 1843 661 1846
rect 650 1803 653 1826
rect 626 1743 637 1746
rect 594 1713 605 1716
rect 570 1693 581 1696
rect 570 1603 573 1626
rect 578 1566 581 1693
rect 594 1646 597 1713
rect 594 1643 605 1646
rect 586 1613 589 1626
rect 586 1603 597 1606
rect 578 1563 589 1566
rect 546 1543 557 1546
rect 514 1483 517 1526
rect 466 1413 469 1426
rect 482 1296 485 1476
rect 490 1376 493 1466
rect 498 1393 501 1416
rect 490 1373 497 1376
rect 474 1293 485 1296
rect 474 1213 477 1293
rect 494 1286 497 1373
rect 506 1323 509 1416
rect 514 1413 517 1426
rect 530 1413 533 1486
rect 546 1456 549 1543
rect 546 1453 557 1456
rect 514 1363 517 1406
rect 538 1403 541 1426
rect 554 1413 557 1453
rect 554 1333 557 1346
rect 546 1313 549 1326
rect 554 1303 557 1326
rect 490 1283 497 1286
rect 442 1153 461 1156
rect 442 1116 445 1153
rect 458 1133 461 1146
rect 434 1113 445 1116
rect 434 1046 437 1113
rect 434 1043 441 1046
rect 346 1003 349 1016
rect 378 1006 381 1016
rect 386 1013 389 1026
rect 418 1023 429 1026
rect 394 1006 397 1016
rect 378 1003 397 1006
rect 402 976 405 1016
rect 418 1013 421 1023
rect 410 983 413 1006
rect 402 973 413 976
rect 298 963 325 966
rect 290 923 293 936
rect 322 896 325 963
rect 338 913 341 926
rect 314 893 325 896
rect 250 843 277 846
rect 242 833 253 836
rect 226 813 237 816
rect 242 813 245 826
rect 250 813 253 833
rect 74 753 85 756
rect 90 773 109 776
rect 194 783 213 786
rect 74 656 77 753
rect 90 656 93 773
rect 138 713 141 726
rect 170 723 173 736
rect 178 713 181 726
rect 74 653 85 656
rect 90 653 125 656
rect 82 503 85 653
rect 98 533 101 546
rect 106 523 109 616
rect 122 556 125 653
rect 162 593 165 616
rect 114 553 125 556
rect 82 193 85 406
rect 114 393 117 553
rect 130 516 133 536
rect 130 513 141 516
rect 138 466 141 513
rect 130 463 141 466
rect 130 413 133 463
rect 162 413 165 536
rect 170 533 173 616
rect 170 486 173 526
rect 186 523 189 606
rect 194 513 197 783
rect 202 613 205 626
rect 202 533 205 606
rect 202 493 205 526
rect 210 523 213 726
rect 218 683 221 736
rect 226 733 229 806
rect 234 623 237 813
rect 250 766 253 806
rect 258 803 261 816
rect 266 813 269 836
rect 274 803 277 843
rect 314 786 317 893
rect 242 763 253 766
rect 298 783 317 786
rect 242 716 245 763
rect 250 733 253 756
rect 258 733 269 736
rect 242 713 249 716
rect 246 626 249 713
rect 242 623 249 626
rect 218 543 221 616
rect 234 586 237 616
rect 242 603 245 623
rect 226 583 237 586
rect 170 483 189 486
rect 130 323 133 336
rect 170 333 173 416
rect 178 323 181 416
rect 186 413 189 483
rect 186 396 189 406
rect 194 403 197 416
rect 202 396 205 416
rect 186 393 205 396
rect 210 376 213 516
rect 226 493 229 583
rect 258 576 261 726
rect 266 716 269 733
rect 266 713 277 716
rect 274 626 277 713
rect 266 623 277 626
rect 266 603 269 623
rect 290 613 293 626
rect 234 533 237 576
rect 242 573 261 576
rect 242 513 245 573
rect 250 523 253 536
rect 202 373 213 376
rect 202 256 205 373
rect 202 253 213 256
rect 130 213 133 226
rect 162 213 165 236
rect 170 213 173 226
rect 186 213 189 226
rect 186 196 189 206
rect 194 203 197 236
rect 202 196 205 216
rect 210 203 213 253
rect 218 213 221 256
rect 226 213 229 426
rect 250 333 253 506
rect 266 393 269 536
rect 282 286 285 416
rect 298 413 301 783
rect 322 736 325 806
rect 362 766 365 816
rect 370 803 373 926
rect 378 913 381 926
rect 402 813 405 936
rect 410 933 413 973
rect 418 923 421 1006
rect 438 966 441 1043
rect 450 1033 453 1126
rect 466 1103 469 1126
rect 450 983 453 1006
rect 458 966 461 1016
rect 474 1013 477 1136
rect 490 1046 493 1283
rect 562 1226 565 1536
rect 570 1496 573 1536
rect 578 1523 581 1546
rect 586 1533 589 1563
rect 602 1533 605 1643
rect 610 1603 613 1736
rect 610 1533 613 1546
rect 586 1513 589 1526
rect 570 1493 581 1496
rect 570 1403 573 1416
rect 570 1323 573 1366
rect 578 1343 581 1493
rect 594 1413 597 1426
rect 602 1413 605 1526
rect 618 1486 621 1726
rect 626 1703 629 1726
rect 610 1483 621 1486
rect 610 1416 613 1483
rect 634 1473 637 1743
rect 650 1733 653 1756
rect 658 1733 661 1843
rect 666 1813 669 1906
rect 698 1886 701 1946
rect 706 1933 709 2006
rect 722 1933 725 2023
rect 722 1893 725 1926
rect 698 1883 717 1886
rect 666 1793 669 1806
rect 674 1726 677 1806
rect 642 1723 677 1726
rect 658 1576 661 1716
rect 674 1706 677 1723
rect 670 1703 677 1706
rect 670 1596 673 1703
rect 670 1593 677 1596
rect 650 1573 661 1576
rect 674 1573 677 1593
rect 650 1516 653 1573
rect 682 1566 685 1816
rect 714 1803 717 1883
rect 722 1803 725 1886
rect 730 1866 733 2006
rect 742 1956 745 2113
rect 758 2106 761 2153
rect 754 2103 761 2106
rect 754 1966 757 2103
rect 770 2003 773 2226
rect 778 2183 781 2216
rect 786 2203 789 2243
rect 802 2233 805 2303
rect 794 2193 797 2216
rect 802 2213 813 2216
rect 802 2176 805 2213
rect 818 2206 821 2286
rect 850 2236 853 2303
rect 798 2173 805 2176
rect 810 2203 821 2206
rect 798 2126 801 2173
rect 810 2133 813 2203
rect 826 2186 829 2236
rect 850 2233 861 2236
rect 858 2213 861 2233
rect 822 2183 829 2186
rect 786 2083 789 2126
rect 798 2123 805 2126
rect 802 2026 805 2123
rect 822 2116 825 2183
rect 818 2113 825 2116
rect 802 2023 809 2026
rect 754 1963 765 1966
rect 742 1953 749 1956
rect 746 1936 749 1953
rect 746 1933 753 1936
rect 738 1883 741 1926
rect 750 1886 753 1933
rect 746 1883 753 1886
rect 730 1863 737 1866
rect 734 1796 737 1863
rect 746 1843 749 1883
rect 762 1866 765 1963
rect 786 1933 789 1946
rect 794 1923 797 2016
rect 806 1936 809 2023
rect 802 1933 809 1936
rect 802 1916 805 1933
rect 758 1863 765 1866
rect 794 1913 805 1916
rect 730 1793 737 1796
rect 690 1713 693 1736
rect 706 1733 709 1746
rect 730 1676 733 1793
rect 722 1673 733 1676
rect 722 1606 725 1673
rect 738 1613 741 1726
rect 746 1723 749 1816
rect 758 1776 761 1863
rect 754 1773 761 1776
rect 754 1703 757 1773
rect 770 1636 773 1736
rect 754 1633 773 1636
rect 722 1603 733 1606
rect 666 1563 685 1566
rect 666 1523 669 1563
rect 674 1533 677 1556
rect 690 1526 693 1576
rect 682 1523 693 1526
rect 650 1513 661 1516
rect 658 1426 661 1513
rect 658 1423 665 1426
rect 610 1413 629 1416
rect 610 1393 613 1406
rect 578 1313 581 1336
rect 602 1246 605 1346
rect 610 1313 613 1326
rect 618 1323 621 1406
rect 626 1313 629 1413
rect 634 1303 637 1416
rect 642 1393 645 1406
rect 642 1333 645 1386
rect 602 1243 621 1246
rect 538 1213 541 1226
rect 558 1223 565 1226
rect 558 1176 561 1223
rect 570 1183 573 1216
rect 578 1213 581 1226
rect 558 1173 565 1176
rect 490 1043 501 1046
rect 474 966 477 1006
rect 498 993 501 1043
rect 514 1013 517 1126
rect 562 1016 565 1173
rect 586 1163 589 1216
rect 602 1136 605 1243
rect 610 1196 613 1206
rect 618 1203 621 1243
rect 626 1196 629 1216
rect 610 1193 629 1196
rect 634 1183 637 1206
rect 642 1136 645 1316
rect 650 1283 653 1416
rect 662 1356 665 1423
rect 682 1416 685 1523
rect 722 1513 725 1526
rect 730 1426 733 1603
rect 754 1566 757 1633
rect 762 1603 765 1626
rect 754 1563 761 1566
rect 758 1486 761 1563
rect 770 1523 773 1616
rect 722 1423 733 1426
rect 754 1483 761 1486
rect 658 1353 665 1356
rect 594 1133 605 1136
rect 634 1133 645 1136
rect 594 1026 597 1133
rect 554 1013 565 1016
rect 586 1023 597 1026
rect 438 963 445 966
rect 458 963 469 966
rect 474 963 485 966
rect 442 886 445 963
rect 466 923 469 963
rect 482 916 485 963
rect 554 946 557 1013
rect 554 943 565 946
rect 474 913 485 916
rect 554 913 557 926
rect 442 883 453 886
rect 362 763 369 766
rect 322 733 333 736
rect 306 613 309 686
rect 314 603 317 616
rect 322 613 325 733
rect 346 713 349 726
rect 366 686 369 763
rect 378 703 381 726
rect 386 713 389 726
rect 362 683 369 686
rect 330 596 333 616
rect 314 593 333 596
rect 338 593 341 606
rect 314 523 317 593
rect 346 523 349 616
rect 354 456 357 526
rect 346 453 357 456
rect 298 393 301 406
rect 322 396 325 416
rect 346 413 349 453
rect 362 423 365 683
rect 386 596 389 606
rect 394 603 397 616
rect 402 596 405 616
rect 386 593 405 596
rect 370 516 373 556
rect 386 543 405 546
rect 386 533 389 543
rect 370 513 381 516
rect 378 426 381 513
rect 370 423 381 426
rect 314 393 325 396
rect 298 313 301 326
rect 282 283 309 286
rect 146 133 149 196
rect 186 193 205 196
rect 218 193 221 206
rect 194 113 197 126
rect 226 123 229 206
rect 242 133 245 216
rect 266 213 269 276
rect 250 193 253 206
rect 274 193 277 206
rect 282 133 285 216
rect 290 203 293 216
rect 298 213 301 226
rect 306 213 309 283
rect 298 193 301 206
rect 314 133 317 393
rect 322 333 341 336
rect 322 213 325 333
rect 330 203 333 326
rect 338 313 341 326
rect 354 303 357 336
rect 362 296 365 416
rect 370 383 373 423
rect 394 413 397 536
rect 402 523 405 543
rect 410 533 413 806
rect 434 776 437 836
rect 450 803 453 883
rect 474 846 477 913
rect 474 843 485 846
rect 482 796 485 843
rect 498 813 501 826
rect 530 803 533 816
rect 538 813 541 826
rect 474 793 485 796
rect 434 773 461 776
rect 426 743 445 746
rect 426 733 429 743
rect 418 613 421 626
rect 426 413 429 726
rect 434 703 437 736
rect 442 723 445 743
rect 450 716 453 746
rect 458 733 461 773
rect 474 763 477 793
rect 442 613 445 716
rect 450 713 457 716
rect 466 713 469 736
rect 454 646 457 713
rect 450 643 457 646
rect 434 593 437 606
rect 434 503 437 526
rect 442 523 445 536
rect 378 403 389 406
rect 434 403 437 416
rect 378 336 381 403
rect 442 396 445 416
rect 450 403 453 643
rect 458 613 461 626
rect 514 613 517 726
rect 522 713 525 736
rect 530 716 533 766
rect 546 756 549 806
rect 554 803 557 826
rect 546 753 557 756
rect 546 733 549 746
rect 554 723 557 753
rect 530 713 541 716
rect 538 656 541 713
rect 534 653 541 656
rect 534 606 537 653
rect 562 626 565 943
rect 570 903 573 926
rect 578 906 581 1006
rect 586 1003 589 1023
rect 610 1016 613 1026
rect 594 993 597 1016
rect 602 1013 613 1016
rect 618 1013 621 1126
rect 626 993 629 1006
rect 586 923 589 986
rect 594 913 597 936
rect 578 903 597 906
rect 570 733 573 806
rect 578 733 581 816
rect 586 813 589 836
rect 594 806 597 903
rect 602 813 605 826
rect 586 803 597 806
rect 586 733 589 803
rect 558 623 565 626
rect 466 533 469 566
rect 490 553 493 606
rect 534 603 541 606
rect 458 513 461 526
rect 474 523 477 536
rect 458 413 461 506
rect 482 413 485 536
rect 490 533 493 546
rect 498 493 501 526
rect 506 523 509 536
rect 514 503 517 536
rect 522 533 525 596
rect 538 436 541 603
rect 558 566 561 623
rect 570 593 573 616
rect 578 603 581 616
rect 602 576 605 736
rect 618 706 621 926
rect 634 923 637 1133
rect 650 923 653 1226
rect 658 1196 661 1353
rect 674 1343 677 1416
rect 682 1413 693 1416
rect 682 1403 693 1406
rect 666 1306 669 1336
rect 674 1323 677 1336
rect 690 1326 693 1346
rect 698 1333 701 1406
rect 690 1323 701 1326
rect 666 1303 677 1306
rect 674 1236 677 1303
rect 666 1233 677 1236
rect 666 1213 669 1233
rect 658 1193 665 1196
rect 662 1056 665 1193
rect 690 1156 693 1306
rect 698 1213 701 1323
rect 722 1246 725 1423
rect 738 1323 741 1416
rect 754 1363 757 1483
rect 778 1446 781 1846
rect 786 1733 789 1856
rect 794 1793 797 1913
rect 818 1853 821 2113
rect 834 2003 837 2206
rect 842 1976 845 2126
rect 850 2106 853 2146
rect 858 2123 861 2196
rect 870 2186 873 2303
rect 882 2196 885 2576
rect 890 2243 893 2536
rect 898 2476 901 2826
rect 914 2823 925 2826
rect 906 2723 909 2816
rect 922 2776 925 2823
rect 914 2773 925 2776
rect 934 2776 937 2843
rect 934 2773 941 2776
rect 914 2716 917 2773
rect 910 2713 917 2716
rect 910 2546 913 2713
rect 922 2563 925 2726
rect 938 2683 941 2773
rect 930 2606 933 2626
rect 946 2623 949 3006
rect 954 2996 957 3303
rect 982 3296 985 3343
rect 978 3293 985 3296
rect 962 3203 965 3216
rect 962 3116 965 3136
rect 962 3113 969 3116
rect 966 3036 969 3113
rect 962 3033 969 3036
rect 962 3016 965 3033
rect 962 3013 973 3016
rect 954 2993 965 2996
rect 962 2826 965 2993
rect 954 2823 965 2826
rect 938 2613 949 2616
rect 930 2603 941 2606
rect 906 2543 913 2546
rect 906 2523 909 2543
rect 922 2503 925 2526
rect 930 2486 933 2536
rect 926 2483 933 2486
rect 898 2473 917 2476
rect 898 2283 901 2436
rect 914 2396 917 2473
rect 926 2416 929 2483
rect 926 2413 933 2416
rect 914 2393 921 2396
rect 906 2313 909 2386
rect 918 2306 921 2393
rect 930 2346 933 2413
rect 938 2353 941 2603
rect 946 2573 949 2606
rect 954 2596 957 2823
rect 962 2723 965 2806
rect 970 2743 973 2766
rect 978 2716 981 3293
rect 994 3223 997 3326
rect 1006 3246 1009 3343
rect 1006 3243 1013 3246
rect 1002 3213 1005 3226
rect 994 3173 997 3196
rect 994 3133 997 3156
rect 986 3123 997 3126
rect 994 3106 997 3123
rect 990 3103 997 3106
rect 990 3006 993 3103
rect 1002 3013 1005 3126
rect 990 3003 997 3006
rect 994 2833 997 3003
rect 1002 2923 1005 2946
rect 1002 2816 1005 2846
rect 1010 2823 1013 3243
rect 1018 3133 1021 3393
rect 1026 3313 1029 3336
rect 1026 3126 1029 3236
rect 1034 3186 1037 3376
rect 1042 3193 1045 3956
rect 1054 3876 1057 3993
rect 1074 3966 1077 3986
rect 1074 3963 1081 3966
rect 1078 3886 1081 3963
rect 1090 3923 1093 4136
rect 1098 4133 1105 4136
rect 1102 4026 1105 4133
rect 1098 4023 1105 4026
rect 1074 3883 1081 3886
rect 1054 3873 1061 3876
rect 1058 3786 1061 3873
rect 1050 3783 1061 3786
rect 1050 3763 1053 3783
rect 1050 3716 1053 3736
rect 1050 3713 1061 3716
rect 1058 3646 1061 3713
rect 1050 3643 1061 3646
rect 1050 3253 1053 3643
rect 1074 3626 1077 3883
rect 1082 3813 1085 3826
rect 1090 3803 1093 3816
rect 1098 3766 1101 4023
rect 1106 3983 1109 4006
rect 1114 4003 1117 4233
rect 1122 4196 1125 4216
rect 1130 4203 1133 4236
rect 1138 4213 1141 4326
rect 1146 4306 1149 4406
rect 1162 4356 1165 4413
rect 1154 4353 1165 4356
rect 1234 4353 1237 4516
rect 1250 4506 1253 4523
rect 1246 4503 1253 4506
rect 1246 4396 1249 4503
rect 1258 4403 1261 4516
rect 1274 4473 1277 4536
rect 1306 4533 1309 4546
rect 1314 4533 1317 4616
rect 1370 4603 1373 4616
rect 1346 4526 1349 4596
rect 1394 4593 1397 4606
rect 1282 4523 1301 4526
rect 1282 4503 1285 4516
rect 1290 4456 1293 4523
rect 1306 4513 1309 4526
rect 1338 4523 1349 4526
rect 1362 4523 1365 4546
rect 1418 4533 1421 4616
rect 1426 4523 1429 4536
rect 1442 4533 1445 4606
rect 1506 4596 1509 4616
rect 1506 4593 1517 4596
rect 1530 4593 1533 4606
rect 1490 4533 1493 4566
rect 1282 4453 1293 4456
rect 1266 4423 1269 4436
rect 1282 4416 1285 4453
rect 1266 4413 1285 4416
rect 1246 4393 1253 4396
rect 1154 4323 1157 4353
rect 1162 4323 1165 4336
rect 1146 4303 1157 4306
rect 1170 4303 1173 4326
rect 1202 4323 1205 4336
rect 1250 4333 1253 4393
rect 1266 4373 1269 4406
rect 1266 4333 1269 4346
rect 1154 4236 1157 4303
rect 1146 4233 1157 4236
rect 1138 4196 1141 4206
rect 1122 4193 1141 4196
rect 1146 4146 1149 4233
rect 1138 4143 1149 4146
rect 1130 4033 1133 4136
rect 1138 4023 1141 4143
rect 1130 4003 1133 4016
rect 1146 4013 1149 4136
rect 1154 4096 1157 4216
rect 1170 4203 1173 4216
rect 1178 4213 1181 4236
rect 1210 4203 1213 4216
rect 1274 4213 1277 4356
rect 1282 4326 1285 4413
rect 1290 4403 1293 4436
rect 1298 4423 1301 4446
rect 1298 4383 1301 4406
rect 1282 4323 1293 4326
rect 1258 4166 1261 4206
rect 1274 4193 1277 4206
rect 1258 4163 1269 4166
rect 1162 4113 1165 4146
rect 1178 4123 1181 4136
rect 1186 4123 1197 4126
rect 1218 4123 1221 4136
rect 1154 4093 1165 4096
rect 1162 3993 1165 4093
rect 1170 3996 1173 4016
rect 1170 3993 1177 3996
rect 1106 3906 1109 3926
rect 1106 3903 1117 3906
rect 1114 3846 1117 3903
rect 1106 3843 1117 3846
rect 1106 3786 1109 3843
rect 1114 3803 1117 3826
rect 1106 3783 1117 3786
rect 1090 3763 1101 3766
rect 1090 3706 1093 3763
rect 1098 3713 1101 3756
rect 1090 3703 1101 3706
rect 1066 3613 1069 3626
rect 1074 3623 1085 3626
rect 1058 3473 1061 3606
rect 1074 3593 1077 3623
rect 1082 3463 1085 3606
rect 1090 3603 1093 3636
rect 1098 3603 1101 3703
rect 1114 3636 1117 3783
rect 1130 3733 1133 3926
rect 1154 3823 1157 3906
rect 1174 3886 1177 3993
rect 1170 3883 1177 3886
rect 1170 3816 1173 3883
rect 1186 3866 1189 4026
rect 1194 4003 1197 4123
rect 1234 3943 1237 4006
rect 1242 3993 1245 4026
rect 1250 4003 1253 4066
rect 1258 3936 1261 4036
rect 1266 3963 1269 4163
rect 1282 4133 1285 4146
rect 1290 4126 1293 4323
rect 1306 4313 1309 4426
rect 1314 4403 1317 4416
rect 1322 4403 1325 4426
rect 1338 4366 1341 4523
rect 1434 4513 1437 4526
rect 1386 4393 1389 4416
rect 1434 4413 1437 4426
rect 1330 4363 1341 4366
rect 1314 4323 1317 4336
rect 1330 4303 1333 4363
rect 1378 4323 1381 4346
rect 1466 4336 1469 4526
rect 1482 4513 1485 4526
rect 1498 4523 1501 4536
rect 1506 4523 1509 4546
rect 1514 4533 1517 4593
rect 1530 4533 1541 4536
rect 1482 4413 1485 4426
rect 1522 4416 1525 4526
rect 1514 4413 1525 4416
rect 1490 4393 1493 4406
rect 1458 4333 1469 4336
rect 1482 4333 1485 4346
rect 1434 4323 1445 4326
rect 1290 4123 1301 4126
rect 1162 3813 1173 3816
rect 1182 3863 1189 3866
rect 1106 3633 1117 3636
rect 1106 3473 1109 3633
rect 1130 3523 1133 3616
rect 1138 3516 1141 3616
rect 1146 3596 1149 3806
rect 1162 3713 1165 3813
rect 1170 3793 1173 3806
rect 1182 3746 1185 3863
rect 1194 3813 1197 3926
rect 1218 3923 1221 3936
rect 1234 3903 1237 3936
rect 1250 3933 1261 3936
rect 1182 3743 1189 3746
rect 1162 3613 1165 3656
rect 1178 3643 1181 3726
rect 1162 3596 1165 3606
rect 1170 3603 1173 3626
rect 1178 3596 1181 3616
rect 1146 3593 1153 3596
rect 1162 3593 1181 3596
rect 1130 3513 1141 3516
rect 1058 3413 1061 3436
rect 1066 3403 1077 3406
rect 1082 3366 1085 3406
rect 1058 3363 1085 3366
rect 1034 3183 1045 3186
rect 1018 3123 1029 3126
rect 1018 3093 1021 3123
rect 1034 3116 1037 3136
rect 1026 3113 1037 3116
rect 1026 3086 1029 3113
rect 1022 3083 1029 3086
rect 1022 2956 1025 3083
rect 1034 3013 1037 3026
rect 1018 2953 1025 2956
rect 994 2756 997 2816
rect 1002 2813 1013 2816
rect 986 2753 997 2756
rect 986 2733 989 2753
rect 962 2613 965 2696
rect 954 2593 961 2596
rect 946 2443 949 2546
rect 958 2436 961 2593
rect 954 2433 961 2436
rect 930 2343 949 2346
rect 930 2323 933 2336
rect 914 2303 921 2306
rect 898 2213 901 2236
rect 914 2213 917 2303
rect 882 2193 893 2196
rect 870 2183 877 2186
rect 874 2146 877 2183
rect 874 2143 881 2146
rect 850 2103 857 2106
rect 854 2036 857 2103
rect 850 2033 857 2036
rect 850 2013 853 2033
rect 850 1993 861 1996
rect 866 1986 869 2136
rect 826 1973 845 1976
rect 858 1983 869 1986
rect 826 1933 829 1973
rect 834 1876 837 1966
rect 826 1873 837 1876
rect 786 1713 789 1726
rect 794 1646 797 1746
rect 802 1723 805 1816
rect 810 1766 813 1796
rect 810 1763 817 1766
rect 814 1696 817 1763
rect 826 1743 829 1873
rect 842 1716 845 1816
rect 858 1813 861 1983
rect 878 1976 881 2143
rect 874 1973 881 1976
rect 874 1846 877 1973
rect 870 1843 877 1846
rect 870 1766 873 1843
rect 890 1836 893 2193
rect 906 2186 909 2206
rect 882 1833 893 1836
rect 902 2183 909 2186
rect 870 1763 877 1766
rect 850 1743 869 1746
rect 874 1743 877 1763
rect 850 1733 853 1743
rect 858 1723 861 1736
rect 866 1723 869 1743
rect 834 1696 837 1716
rect 842 1713 853 1716
rect 810 1693 817 1696
rect 826 1693 837 1696
rect 810 1673 813 1693
rect 826 1646 829 1693
rect 794 1643 801 1646
rect 826 1643 837 1646
rect 786 1613 789 1636
rect 798 1586 801 1643
rect 826 1613 829 1626
rect 810 1593 813 1606
rect 798 1583 805 1586
rect 818 1583 821 1606
rect 834 1603 837 1643
rect 778 1443 785 1446
rect 770 1413 773 1436
rect 782 1366 785 1443
rect 802 1436 805 1583
rect 818 1513 821 1536
rect 794 1433 805 1436
rect 794 1386 797 1433
rect 810 1413 813 1426
rect 810 1396 813 1406
rect 818 1403 821 1416
rect 826 1396 829 1416
rect 810 1393 829 1396
rect 834 1393 837 1406
rect 794 1383 805 1386
rect 782 1363 789 1366
rect 722 1243 733 1246
rect 730 1223 733 1243
rect 738 1213 741 1286
rect 762 1236 765 1346
rect 778 1343 781 1356
rect 786 1306 789 1363
rect 794 1326 797 1366
rect 802 1343 805 1383
rect 842 1326 845 1706
rect 850 1696 853 1713
rect 850 1693 861 1696
rect 858 1646 861 1693
rect 850 1643 861 1646
rect 850 1613 853 1643
rect 874 1626 877 1736
rect 882 1733 885 1833
rect 902 1816 905 2183
rect 898 1813 905 1816
rect 890 1743 893 1756
rect 866 1623 877 1626
rect 858 1523 861 1596
rect 850 1393 853 1446
rect 794 1323 805 1326
rect 754 1233 765 1236
rect 770 1303 789 1306
rect 698 1183 701 1206
rect 730 1203 741 1206
rect 682 1153 693 1156
rect 658 1053 665 1056
rect 658 1003 661 1053
rect 658 933 661 956
rect 666 903 669 1036
rect 674 1003 677 1136
rect 682 1083 685 1153
rect 698 1096 701 1166
rect 754 1163 757 1233
rect 746 1103 749 1126
rect 694 1093 701 1096
rect 694 1036 697 1093
rect 706 1046 709 1086
rect 706 1043 717 1046
rect 682 1013 685 1036
rect 694 1033 701 1036
rect 634 793 637 806
rect 642 803 645 816
rect 650 813 653 826
rect 658 803 661 816
rect 634 733 637 766
rect 658 723 661 736
rect 618 703 637 706
rect 674 703 677 806
rect 682 783 685 1006
rect 698 983 701 1033
rect 714 976 717 1043
rect 730 993 733 1016
rect 706 973 717 976
rect 706 826 709 973
rect 714 933 717 946
rect 730 933 733 986
rect 762 976 765 1226
rect 770 1003 773 1303
rect 778 1213 781 1296
rect 802 1256 805 1323
rect 794 1253 805 1256
rect 834 1323 845 1326
rect 794 1236 797 1253
rect 790 1233 797 1236
rect 778 1093 781 1206
rect 790 1186 793 1233
rect 802 1193 805 1206
rect 810 1196 813 1216
rect 818 1203 821 1236
rect 826 1196 829 1206
rect 810 1193 829 1196
rect 834 1186 837 1323
rect 866 1216 869 1623
rect 874 1533 877 1616
rect 874 1503 877 1526
rect 882 1406 885 1706
rect 890 1673 893 1726
rect 890 1593 893 1606
rect 890 1543 893 1556
rect 898 1526 901 1813
rect 894 1523 901 1526
rect 894 1416 897 1523
rect 894 1413 901 1416
rect 878 1403 885 1406
rect 878 1356 881 1403
rect 890 1383 893 1396
rect 898 1366 901 1413
rect 906 1403 909 1746
rect 914 1533 917 2206
rect 922 2106 925 2246
rect 930 2123 933 2316
rect 938 2213 941 2336
rect 922 2103 929 2106
rect 926 1646 929 2103
rect 922 1643 929 1646
rect 922 1526 925 1643
rect 938 1613 941 2206
rect 946 2153 949 2343
rect 954 2333 957 2433
rect 970 2366 973 2716
rect 978 2713 985 2716
rect 982 2606 985 2713
rect 994 2703 997 2726
rect 994 2613 997 2646
rect 982 2603 989 2606
rect 966 2363 973 2366
rect 966 2316 969 2363
rect 978 2316 981 2356
rect 986 2333 989 2603
rect 1002 2596 1005 2806
rect 998 2593 1005 2596
rect 998 2546 1001 2593
rect 1010 2556 1013 2806
rect 1018 2643 1021 2953
rect 1026 2906 1029 2936
rect 1034 2923 1037 2966
rect 1026 2903 1033 2906
rect 1030 2756 1033 2903
rect 1042 2813 1045 3183
rect 1050 2863 1053 3226
rect 1058 3153 1061 3363
rect 1066 3313 1069 3326
rect 1074 3323 1077 3336
rect 1066 3213 1069 3226
rect 1058 3013 1061 3136
rect 1058 2906 1061 2936
rect 1066 2923 1069 3196
rect 1074 3063 1077 3256
rect 1082 3233 1085 3346
rect 1098 3216 1101 3236
rect 1090 3213 1101 3216
rect 1106 3213 1109 3466
rect 1122 3413 1125 3426
rect 1130 3413 1133 3513
rect 1150 3506 1153 3593
rect 1186 3576 1189 3743
rect 1194 3723 1197 3796
rect 1194 3613 1197 3646
rect 1202 3623 1205 3736
rect 1210 3733 1213 3786
rect 1178 3573 1189 3576
rect 1178 3516 1181 3573
rect 1194 3523 1197 3606
rect 1178 3513 1189 3516
rect 1146 3503 1153 3506
rect 1146 3433 1149 3503
rect 1146 3396 1149 3416
rect 1154 3403 1157 3446
rect 1162 3396 1165 3406
rect 1146 3393 1165 3396
rect 1170 3343 1173 3416
rect 1186 3393 1189 3513
rect 1194 3376 1197 3436
rect 1190 3373 1197 3376
rect 1178 3343 1181 3366
rect 1154 3306 1157 3326
rect 1138 3303 1157 3306
rect 1138 3206 1141 3303
rect 1162 3286 1165 3336
rect 1170 3316 1173 3336
rect 1170 3313 1181 3316
rect 1154 3283 1165 3286
rect 1154 3236 1157 3283
rect 1178 3246 1181 3313
rect 1190 3306 1193 3373
rect 1202 3333 1205 3536
rect 1210 3533 1213 3546
rect 1210 3373 1213 3456
rect 1202 3313 1205 3326
rect 1190 3303 1197 3306
rect 1170 3243 1181 3246
rect 1154 3233 1165 3236
rect 1162 3213 1165 3233
rect 1170 3223 1173 3243
rect 1194 3216 1197 3303
rect 1186 3213 1197 3216
rect 1210 3213 1213 3336
rect 1218 3316 1221 3766
rect 1226 3733 1229 3746
rect 1234 3623 1237 3806
rect 1250 3723 1253 3933
rect 1274 3886 1277 4016
rect 1282 4003 1285 4066
rect 1290 4023 1293 4116
rect 1298 4016 1301 4123
rect 1306 4113 1309 4216
rect 1338 4193 1341 4206
rect 1330 4123 1333 4136
rect 1338 4133 1341 4156
rect 1346 4133 1349 4216
rect 1402 4183 1405 4216
rect 1378 4146 1381 4166
rect 1370 4143 1381 4146
rect 1338 4063 1341 4126
rect 1290 4013 1309 4016
rect 1290 3993 1293 4006
rect 1266 3883 1277 3886
rect 1258 3693 1261 3736
rect 1266 3723 1269 3883
rect 1290 3846 1293 3866
rect 1282 3843 1293 3846
rect 1282 3776 1285 3843
rect 1298 3786 1301 3926
rect 1322 3913 1325 3936
rect 1330 3923 1333 4006
rect 1370 3986 1373 4143
rect 1394 3996 1397 4136
rect 1402 4106 1405 4166
rect 1426 4133 1429 4306
rect 1442 4193 1445 4216
rect 1434 4133 1437 4186
rect 1458 4163 1461 4333
rect 1466 4323 1477 4326
rect 1506 4263 1509 4336
rect 1458 4126 1461 4136
rect 1410 4123 1429 4126
rect 1450 4123 1461 4126
rect 1450 4106 1453 4123
rect 1466 4106 1469 4136
rect 1402 4103 1413 4106
rect 1410 4036 1413 4103
rect 1402 4033 1413 4036
rect 1442 4103 1453 4106
rect 1462 4103 1469 4106
rect 1442 4036 1445 4103
rect 1462 4036 1465 4103
rect 1474 4096 1477 4256
rect 1482 4133 1485 4186
rect 1474 4093 1485 4096
rect 1442 4033 1453 4036
rect 1462 4033 1469 4036
rect 1402 4003 1405 4033
rect 1418 4013 1437 4016
rect 1450 4013 1453 4033
rect 1466 4016 1469 4033
rect 1466 4013 1473 4016
rect 1394 3993 1413 3996
rect 1370 3983 1381 3986
rect 1346 3946 1349 3966
rect 1342 3943 1349 3946
rect 1342 3886 1345 3943
rect 1370 3906 1373 3926
rect 1366 3903 1373 3906
rect 1342 3883 1349 3886
rect 1346 3846 1349 3883
rect 1346 3843 1353 3846
rect 1306 3803 1309 3816
rect 1298 3783 1317 3786
rect 1282 3773 1293 3776
rect 1290 3756 1293 3773
rect 1290 3753 1297 3756
rect 1234 3523 1237 3606
rect 1266 3593 1269 3606
rect 1274 3576 1277 3616
rect 1270 3573 1277 3576
rect 1226 3333 1229 3446
rect 1234 3413 1237 3426
rect 1250 3416 1253 3446
rect 1242 3413 1253 3416
rect 1258 3413 1261 3536
rect 1270 3506 1273 3573
rect 1270 3503 1277 3506
rect 1282 3503 1285 3726
rect 1274 3486 1277 3503
rect 1274 3483 1285 3486
rect 1274 3413 1277 3426
rect 1218 3313 1225 3316
rect 1222 3236 1225 3313
rect 1218 3233 1225 3236
rect 1082 3056 1085 3206
rect 1114 3186 1117 3206
rect 1138 3203 1157 3206
rect 1114 3183 1133 3186
rect 1090 3136 1093 3156
rect 1090 3133 1097 3136
rect 1074 3053 1085 3056
rect 1058 2903 1065 2906
rect 1062 2856 1065 2903
rect 1058 2853 1065 2856
rect 1026 2753 1033 2756
rect 1026 2613 1029 2753
rect 1034 2683 1037 2736
rect 1042 2716 1045 2766
rect 1050 2723 1053 2746
rect 1058 2733 1061 2853
rect 1066 2733 1069 2776
rect 1074 2763 1077 3053
rect 1094 3046 1097 3133
rect 1106 3123 1109 3136
rect 1130 3066 1133 3183
rect 1154 3133 1157 3203
rect 1162 3186 1165 3206
rect 1162 3183 1173 3186
rect 1170 3126 1173 3183
rect 1090 3043 1097 3046
rect 1082 2773 1085 2936
rect 1090 2933 1093 3043
rect 1098 3013 1101 3026
rect 1090 2913 1093 2926
rect 1042 2713 1049 2716
rect 1058 2713 1061 2726
rect 1066 2723 1077 2726
rect 1046 2656 1049 2713
rect 1082 2703 1085 2736
rect 1058 2666 1061 2686
rect 1058 2663 1065 2666
rect 1046 2653 1053 2656
rect 1026 2586 1029 2606
rect 1018 2583 1029 2586
rect 1018 2563 1021 2583
rect 1042 2576 1045 2596
rect 1026 2573 1045 2576
rect 1010 2553 1021 2556
rect 998 2543 1005 2546
rect 1002 2506 1005 2543
rect 998 2503 1005 2506
rect 998 2326 1001 2503
rect 994 2323 1001 2326
rect 954 2296 957 2316
rect 966 2313 973 2316
rect 978 2313 985 2316
rect 954 2293 961 2296
rect 946 2133 949 2146
rect 958 2126 961 2293
rect 954 2123 961 2126
rect 954 2016 957 2123
rect 970 2106 973 2313
rect 982 2236 985 2313
rect 978 2233 985 2236
rect 978 2213 981 2233
rect 966 2103 973 2106
rect 966 2026 969 2103
rect 978 2036 981 2156
rect 994 2136 997 2323
rect 1010 2313 1013 2496
rect 1018 2476 1021 2553
rect 1026 2496 1029 2573
rect 1034 2523 1037 2536
rect 1050 2513 1053 2653
rect 1062 2586 1065 2663
rect 1074 2613 1077 2626
rect 1058 2583 1065 2586
rect 1058 2516 1061 2583
rect 1066 2523 1069 2566
rect 1074 2533 1077 2606
rect 1058 2513 1065 2516
rect 1026 2493 1037 2496
rect 1018 2473 1025 2476
rect 1022 2396 1025 2473
rect 1018 2393 1025 2396
rect 1002 2213 1005 2296
rect 1018 2213 1021 2393
rect 1034 2376 1037 2493
rect 1062 2456 1065 2513
rect 1062 2453 1069 2456
rect 1026 2373 1037 2376
rect 1026 2296 1029 2373
rect 1026 2293 1033 2296
rect 1030 2226 1033 2293
rect 1030 2223 1037 2226
rect 1026 2193 1029 2216
rect 1034 2146 1037 2223
rect 1042 2183 1045 2346
rect 1058 2343 1061 2436
rect 1034 2143 1045 2146
rect 994 2133 1001 2136
rect 986 2083 989 2126
rect 998 2036 1001 2133
rect 978 2033 989 2036
rect 998 2033 1005 2036
rect 966 2023 973 2026
rect 950 2013 957 2016
rect 950 1916 953 2013
rect 962 1923 965 2006
rect 950 1913 957 1916
rect 954 1813 957 1913
rect 970 1906 973 2023
rect 978 1993 981 2026
rect 986 1906 989 2033
rect 994 2013 997 2026
rect 1002 1996 1005 2033
rect 1010 2023 1013 2136
rect 1034 2116 1037 2136
rect 1026 2113 1037 2116
rect 1026 2036 1029 2113
rect 1026 2033 1037 2036
rect 1034 2013 1037 2033
rect 966 1903 973 1906
rect 978 1903 989 1906
rect 998 1993 1005 1996
rect 966 1826 969 1903
rect 966 1823 973 1826
rect 954 1793 957 1806
rect 962 1733 965 1806
rect 970 1776 973 1823
rect 978 1796 981 1903
rect 986 1813 989 1886
rect 978 1793 989 1796
rect 970 1773 977 1776
rect 930 1543 933 1566
rect 914 1396 917 1526
rect 922 1523 929 1526
rect 926 1436 929 1523
rect 894 1363 901 1366
rect 906 1393 917 1396
rect 922 1433 929 1436
rect 878 1353 885 1356
rect 882 1333 885 1353
rect 894 1256 897 1363
rect 894 1253 901 1256
rect 790 1183 797 1186
rect 786 1103 789 1126
rect 794 1123 797 1183
rect 826 1183 837 1186
rect 858 1213 869 1216
rect 882 1213 885 1226
rect 890 1213 893 1236
rect 826 1103 829 1183
rect 834 1143 853 1146
rect 834 1133 837 1143
rect 786 1013 789 1026
rect 826 1013 829 1026
rect 810 983 813 1006
rect 834 983 837 1126
rect 842 1093 845 1136
rect 850 1123 853 1143
rect 858 1133 861 1213
rect 898 1196 901 1253
rect 890 1193 901 1196
rect 866 1113 869 1156
rect 890 1146 893 1193
rect 874 1133 877 1146
rect 890 1143 901 1146
rect 898 1123 901 1143
rect 906 1136 909 1393
rect 922 1206 925 1433
rect 930 1373 933 1416
rect 938 1273 941 1606
rect 962 1566 965 1726
rect 974 1686 977 1773
rect 954 1563 965 1566
rect 970 1683 977 1686
rect 954 1496 957 1563
rect 970 1503 973 1683
rect 986 1666 989 1793
rect 998 1746 1001 1993
rect 1010 1813 1013 2006
rect 1010 1756 1013 1806
rect 1026 1803 1029 1936
rect 1034 1903 1037 1926
rect 1042 1886 1045 2143
rect 1050 2046 1053 2206
rect 1066 2203 1069 2453
rect 1074 2296 1077 2516
rect 1082 2476 1085 2556
rect 1090 2533 1093 2906
rect 1098 2553 1101 2806
rect 1106 2643 1109 3066
rect 1114 3063 1133 3066
rect 1162 3123 1173 3126
rect 1114 2966 1117 3063
rect 1162 3006 1165 3123
rect 1194 3106 1197 3126
rect 1186 3103 1197 3106
rect 1186 3056 1189 3103
rect 1202 3086 1205 3206
rect 1210 3103 1213 3136
rect 1202 3083 1209 3086
rect 1186 3053 1197 3056
rect 1114 2963 1125 2966
rect 1122 2836 1125 2963
rect 1114 2833 1125 2836
rect 1114 2786 1117 2833
rect 1130 2803 1133 2816
rect 1114 2783 1125 2786
rect 1122 2696 1125 2783
rect 1138 2773 1141 3006
rect 1154 3003 1165 3006
rect 1146 2913 1149 2926
rect 1146 2813 1149 2826
rect 1114 2693 1125 2696
rect 1114 2673 1117 2693
rect 1138 2673 1141 2726
rect 1154 2716 1157 3003
rect 1162 2983 1165 2996
rect 1178 2983 1181 3036
rect 1194 3013 1197 3053
rect 1206 3006 1209 3083
rect 1202 3003 1209 3006
rect 1170 2813 1173 2926
rect 1186 2903 1189 2926
rect 1194 2813 1197 2826
rect 1170 2773 1173 2806
rect 1170 2733 1173 2746
rect 1154 2713 1165 2716
rect 1162 2646 1165 2713
rect 1186 2703 1189 2776
rect 1194 2713 1197 2726
rect 1202 2686 1205 3003
rect 1218 2986 1221 3233
rect 1226 3203 1229 3216
rect 1226 3096 1229 3176
rect 1234 3163 1237 3396
rect 1242 3356 1245 3376
rect 1242 3353 1249 3356
rect 1246 3246 1249 3353
rect 1258 3323 1261 3346
rect 1282 3323 1285 3483
rect 1294 3366 1297 3753
rect 1306 3603 1309 3746
rect 1314 3696 1317 3783
rect 1322 3773 1325 3806
rect 1350 3766 1353 3843
rect 1366 3836 1369 3903
rect 1378 3863 1381 3983
rect 1386 3923 1389 3936
rect 1410 3876 1413 3993
rect 1426 3933 1429 4006
rect 1442 3933 1445 4006
rect 1458 3906 1461 4006
rect 1470 3966 1473 4013
rect 1402 3873 1413 3876
rect 1450 3903 1461 3906
rect 1466 3963 1473 3966
rect 1366 3833 1373 3836
rect 1362 3793 1365 3816
rect 1350 3763 1361 3766
rect 1322 3723 1325 3736
rect 1330 3723 1333 3746
rect 1338 3713 1341 3736
rect 1346 3733 1349 3756
rect 1346 3703 1349 3716
rect 1314 3693 1325 3696
rect 1322 3596 1325 3693
rect 1358 3676 1361 3763
rect 1370 3686 1373 3833
rect 1402 3796 1405 3873
rect 1402 3793 1413 3796
rect 1410 3773 1413 3793
rect 1418 3756 1421 3866
rect 1450 3836 1453 3903
rect 1450 3833 1461 3836
rect 1434 3813 1445 3816
rect 1410 3753 1421 3756
rect 1386 3713 1389 3726
rect 1410 3706 1413 3753
rect 1426 3713 1429 3736
rect 1410 3703 1421 3706
rect 1370 3683 1377 3686
rect 1358 3673 1365 3676
rect 1314 3593 1325 3596
rect 1314 3546 1317 3593
rect 1346 3576 1349 3626
rect 1342 3573 1349 3576
rect 1306 3533 1309 3546
rect 1314 3543 1325 3546
rect 1314 3523 1317 3536
rect 1322 3526 1325 3543
rect 1322 3523 1333 3526
rect 1314 3503 1317 3516
rect 1342 3496 1345 3573
rect 1342 3493 1349 3496
rect 1290 3363 1297 3366
rect 1290 3256 1293 3363
rect 1322 3353 1325 3406
rect 1338 3403 1341 3476
rect 1346 3376 1349 3493
rect 1338 3373 1349 3376
rect 1298 3333 1301 3346
rect 1306 3323 1309 3336
rect 1290 3253 1297 3256
rect 1242 3243 1249 3246
rect 1242 3206 1245 3243
rect 1250 3223 1261 3226
rect 1242 3203 1249 3206
rect 1234 3113 1237 3146
rect 1246 3106 1249 3203
rect 1258 3113 1261 3223
rect 1274 3196 1277 3216
rect 1282 3203 1285 3246
rect 1274 3193 1285 3196
rect 1242 3103 1249 3106
rect 1226 3093 1233 3096
rect 1214 2983 1221 2986
rect 1214 2916 1217 2983
rect 1230 2976 1233 3093
rect 1226 2973 1233 2976
rect 1226 2923 1229 2973
rect 1242 2956 1245 3103
rect 1258 3013 1261 3086
rect 1274 3013 1277 3166
rect 1282 3123 1285 3193
rect 1294 3096 1297 3253
rect 1306 3113 1309 3316
rect 1322 3203 1325 3326
rect 1338 3186 1341 3373
rect 1338 3183 1349 3186
rect 1346 3163 1349 3183
rect 1314 3133 1317 3156
rect 1354 3146 1357 3656
rect 1362 3323 1365 3673
rect 1374 3636 1377 3683
rect 1370 3633 1377 3636
rect 1370 3533 1373 3633
rect 1418 3626 1421 3703
rect 1442 3686 1445 3806
rect 1458 3753 1461 3833
rect 1442 3683 1461 3686
rect 1414 3623 1421 3626
rect 1378 3546 1381 3616
rect 1378 3543 1389 3546
rect 1386 3533 1389 3543
rect 1414 3536 1417 3623
rect 1426 3543 1429 3616
rect 1458 3603 1461 3683
rect 1466 3636 1469 3963
rect 1482 3946 1485 4093
rect 1498 4063 1501 4206
rect 1506 4203 1509 4236
rect 1514 4213 1517 4413
rect 1522 4333 1525 4356
rect 1530 4316 1533 4406
rect 1546 4373 1549 4596
rect 1570 4446 1573 4646
rect 1586 4593 1589 4606
rect 1586 4533 1597 4536
rect 1602 4523 1605 4536
rect 1610 4523 1613 4556
rect 1618 4533 1621 4616
rect 1658 4576 1661 4653
rect 1858 4653 1869 4656
rect 1650 4573 1661 4576
rect 1570 4443 1581 4446
rect 1578 4396 1581 4443
rect 1626 4423 1629 4526
rect 1570 4393 1581 4396
rect 1594 4393 1597 4416
rect 1522 4313 1533 4316
rect 1522 4253 1525 4313
rect 1514 4163 1517 4206
rect 1522 4193 1525 4216
rect 1530 4203 1533 4306
rect 1538 4233 1541 4326
rect 1538 4213 1549 4216
rect 1538 4133 1541 4213
rect 1554 4203 1557 4256
rect 1562 4153 1565 4216
rect 1546 4123 1549 4146
rect 1522 3956 1525 4016
rect 1514 3953 1525 3956
rect 1482 3943 1493 3946
rect 1490 3836 1493 3943
rect 1514 3906 1517 3953
rect 1514 3903 1525 3906
rect 1482 3833 1493 3836
rect 1482 3816 1485 3833
rect 1474 3813 1485 3816
rect 1498 3813 1509 3816
rect 1522 3813 1525 3903
rect 1474 3683 1477 3813
rect 1466 3633 1477 3636
rect 1414 3533 1421 3536
rect 1370 3523 1381 3526
rect 1370 3306 1373 3516
rect 1378 3506 1381 3523
rect 1378 3503 1389 3506
rect 1386 3446 1389 3503
rect 1378 3443 1389 3446
rect 1418 3446 1421 3533
rect 1442 3503 1445 3526
rect 1474 3496 1477 3633
rect 1482 3603 1485 3806
rect 1514 3793 1517 3806
rect 1506 3736 1509 3756
rect 1506 3733 1513 3736
rect 1490 3603 1493 3726
rect 1498 3586 1501 3686
rect 1510 3626 1513 3733
rect 1490 3583 1501 3586
rect 1506 3623 1513 3626
rect 1490 3516 1493 3583
rect 1506 3516 1509 3623
rect 1522 3613 1525 3726
rect 1538 3613 1541 3816
rect 1546 3803 1549 4066
rect 1570 4046 1573 4393
rect 1618 4333 1621 4376
rect 1578 4303 1581 4326
rect 1634 4296 1637 4536
rect 1650 4533 1653 4573
rect 1642 4413 1645 4436
rect 1650 4403 1653 4526
rect 1658 4523 1661 4556
rect 1674 4533 1677 4616
rect 1802 4613 1805 4626
rect 1842 4613 1845 4626
rect 1794 4593 1797 4606
rect 1690 4496 1693 4546
rect 1818 4543 1821 4606
rect 1738 4513 1741 4526
rect 1674 4493 1693 4496
rect 1658 4466 1661 4486
rect 1658 4463 1665 4466
rect 1662 4376 1665 4463
rect 1658 4373 1665 4376
rect 1658 4356 1661 4373
rect 1650 4353 1661 4356
rect 1650 4306 1653 4353
rect 1650 4303 1661 4306
rect 1626 4293 1637 4296
rect 1626 4236 1629 4293
rect 1658 4286 1661 4303
rect 1642 4283 1661 4286
rect 1674 4283 1677 4493
rect 1690 4413 1693 4436
rect 1706 4413 1709 4426
rect 1698 4393 1701 4406
rect 1722 4403 1725 4416
rect 1746 4413 1749 4426
rect 1770 4423 1773 4526
rect 1778 4513 1781 4526
rect 1794 4483 1797 4526
rect 1754 4406 1757 4416
rect 1738 4403 1757 4406
rect 1802 4393 1805 4416
rect 1722 4323 1725 4336
rect 1754 4323 1757 4346
rect 1762 4323 1765 4336
rect 1778 4323 1781 4356
rect 1810 4326 1813 4436
rect 1818 4413 1821 4536
rect 1834 4433 1837 4546
rect 1842 4523 1845 4596
rect 1858 4586 1861 4653
rect 2018 4626 2021 4686
rect 2010 4623 2021 4626
rect 1858 4583 1869 4586
rect 1826 4403 1829 4426
rect 1826 4343 1845 4346
rect 1826 4333 1829 4343
rect 1834 4326 1837 4336
rect 1810 4323 1837 4326
rect 1842 4323 1845 4343
rect 1850 4333 1853 4346
rect 1858 4323 1861 4526
rect 1866 4523 1869 4583
rect 1898 4546 1901 4616
rect 1930 4583 1933 4606
rect 1882 4543 1901 4546
rect 1882 4533 1885 4543
rect 1890 4463 1893 4536
rect 1906 4533 1909 4546
rect 1906 4513 1909 4526
rect 1922 4523 1925 4536
rect 1938 4533 1941 4546
rect 1954 4523 1957 4616
rect 2010 4546 2013 4623
rect 2010 4543 2021 4546
rect 1962 4523 1965 4536
rect 1970 4523 1973 4536
rect 2010 4503 2013 4526
rect 1810 4303 1813 4316
rect 1626 4233 1637 4236
rect 1578 4123 1581 4206
rect 1586 4133 1589 4206
rect 1610 4133 1613 4216
rect 1634 4163 1637 4233
rect 1642 4206 1645 4283
rect 1650 4213 1653 4266
rect 1642 4203 1653 4206
rect 1658 4203 1661 4276
rect 1666 4193 1669 4216
rect 1674 4183 1677 4216
rect 1682 4173 1685 4206
rect 1730 4186 1733 4286
rect 1778 4213 1781 4236
rect 1802 4213 1813 4216
rect 1706 4183 1733 4186
rect 1570 4043 1581 4046
rect 1578 3996 1581 4043
rect 1570 3993 1581 3996
rect 1594 3993 1597 4016
rect 1618 4006 1621 4136
rect 1626 4123 1629 4156
rect 1634 4133 1637 4146
rect 1642 4123 1645 4136
rect 1682 4106 1685 4126
rect 1674 4103 1685 4106
rect 1674 4036 1677 4103
rect 1674 4033 1685 4036
rect 1618 4003 1637 4006
rect 1570 3946 1573 3993
rect 1570 3943 1577 3946
rect 1574 3896 1577 3943
rect 1618 3936 1621 4003
rect 1614 3933 1621 3936
rect 1650 3933 1653 4016
rect 1570 3893 1577 3896
rect 1570 3816 1573 3893
rect 1562 3813 1573 3816
rect 1562 3766 1565 3813
rect 1578 3776 1581 3806
rect 1586 3793 1589 3926
rect 1614 3876 1617 3933
rect 1626 3896 1629 3926
rect 1634 3913 1637 3926
rect 1666 3923 1669 4016
rect 1682 4013 1685 4033
rect 1690 4013 1693 4136
rect 1706 4053 1709 4183
rect 1746 4166 1749 4186
rect 1742 4163 1749 4166
rect 1742 4086 1745 4163
rect 1754 4123 1757 4136
rect 1770 4106 1773 4166
rect 1786 4123 1789 4146
rect 1794 4123 1797 4136
rect 1810 4123 1813 4176
rect 1770 4103 1781 4106
rect 1738 4083 1745 4086
rect 1674 3993 1677 4006
rect 1690 3946 1693 4006
rect 1706 4003 1709 4046
rect 1690 3943 1701 3946
rect 1674 3923 1677 3936
rect 1698 3913 1701 3943
rect 1738 3936 1741 4083
rect 1762 4036 1765 4056
rect 1778 4036 1781 4103
rect 1818 4036 1821 4323
rect 1826 4213 1829 4276
rect 1858 4193 1861 4216
rect 1866 4203 1869 4216
rect 1874 4213 1877 4326
rect 1890 4323 1893 4416
rect 1906 4413 1933 4416
rect 1898 4403 1909 4406
rect 1906 4353 1909 4403
rect 1922 4333 1925 4376
rect 1882 4213 1885 4236
rect 1858 4126 1861 4136
rect 1866 4133 1869 4156
rect 1882 4133 1885 4146
rect 1858 4123 1877 4126
rect 1890 4123 1893 4206
rect 1906 4153 1909 4326
rect 1930 4276 1933 4413
rect 1986 4403 1989 4416
rect 1994 4403 1997 4426
rect 1970 4333 1973 4346
rect 1978 4306 1981 4336
rect 1994 4333 1997 4366
rect 2002 4336 2005 4416
rect 2010 4363 2013 4406
rect 2018 4393 2021 4543
rect 2026 4523 2029 4546
rect 2026 4413 2029 4426
rect 2002 4333 2013 4336
rect 1930 4273 1941 4276
rect 1922 4213 1925 4256
rect 1922 4193 1925 4206
rect 1930 4203 1933 4226
rect 1906 4126 1909 4146
rect 1754 4033 1765 4036
rect 1770 4033 1781 4036
rect 1810 4033 1821 4036
rect 1754 3956 1757 4033
rect 1754 3953 1761 3956
rect 1714 3923 1717 3936
rect 1738 3933 1749 3936
rect 1626 3893 1637 3896
rect 1610 3873 1617 3876
rect 1578 3773 1589 3776
rect 1562 3763 1573 3766
rect 1562 3733 1565 3746
rect 1546 3723 1557 3726
rect 1570 3706 1573 3763
rect 1562 3703 1573 3706
rect 1562 3636 1565 3703
rect 1586 3676 1589 3773
rect 1610 3733 1613 3873
rect 1634 3826 1637 3893
rect 1626 3823 1637 3826
rect 1618 3713 1621 3816
rect 1626 3803 1629 3823
rect 1626 3733 1629 3796
rect 1634 3773 1637 3806
rect 1698 3803 1709 3806
rect 1634 3703 1637 3726
rect 1666 3713 1669 3736
rect 1698 3733 1701 3746
rect 1578 3673 1589 3676
rect 1562 3633 1573 3636
rect 1514 3523 1517 3606
rect 1522 3603 1533 3606
rect 1546 3533 1549 3546
rect 1490 3513 1501 3516
rect 1506 3513 1525 3516
rect 1474 3493 1485 3496
rect 1418 3443 1429 3446
rect 1378 3413 1381 3443
rect 1386 3366 1389 3416
rect 1402 3393 1405 3406
rect 1426 3373 1429 3443
rect 1450 3376 1453 3416
rect 1450 3373 1469 3376
rect 1386 3363 1405 3366
rect 1366 3303 1373 3306
rect 1378 3306 1381 3326
rect 1378 3303 1389 3306
rect 1366 3236 1369 3303
rect 1386 3256 1389 3303
rect 1378 3253 1389 3256
rect 1366 3233 1373 3236
rect 1322 3133 1325 3146
rect 1350 3143 1357 3146
rect 1294 3093 1301 3096
rect 1238 2953 1245 2956
rect 1214 2913 1221 2916
rect 1210 2766 1213 2856
rect 1218 2773 1221 2913
rect 1210 2763 1221 2766
rect 1218 2733 1221 2763
rect 1238 2756 1241 2953
rect 1250 2766 1253 3006
rect 1258 2916 1261 2936
rect 1258 2913 1265 2916
rect 1262 2836 1265 2913
rect 1258 2833 1265 2836
rect 1258 2813 1261 2833
rect 1250 2763 1257 2766
rect 1274 2763 1277 3006
rect 1282 3003 1285 3016
rect 1298 2966 1301 3093
rect 1290 2963 1301 2966
rect 1290 2866 1293 2963
rect 1306 2933 1309 2946
rect 1314 2883 1317 2936
rect 1322 2903 1325 2916
rect 1338 2913 1341 3116
rect 1350 2916 1353 3143
rect 1362 2923 1365 3216
rect 1370 3196 1373 3233
rect 1378 3213 1381 3253
rect 1402 3236 1405 3363
rect 1450 3313 1453 3336
rect 1458 3333 1461 3366
rect 1466 3336 1469 3373
rect 1482 3363 1485 3493
rect 1498 3473 1501 3513
rect 1522 3486 1525 3513
rect 1538 3503 1541 3526
rect 1554 3523 1557 3616
rect 1570 3596 1573 3633
rect 1578 3613 1581 3673
rect 1602 3603 1605 3656
rect 1570 3593 1581 3596
rect 1578 3516 1581 3593
rect 1610 3546 1613 3616
rect 1618 3603 1621 3686
rect 1634 3603 1637 3646
rect 1722 3643 1725 3826
rect 1610 3543 1621 3546
rect 1570 3513 1581 3516
rect 1514 3483 1525 3486
rect 1514 3436 1517 3483
rect 1514 3433 1525 3436
rect 1466 3333 1477 3336
rect 1498 3326 1501 3416
rect 1386 3233 1405 3236
rect 1370 3193 1377 3196
rect 1374 2956 1377 3193
rect 1386 3106 1389 3233
rect 1410 3213 1437 3216
rect 1458 3213 1461 3326
rect 1474 3306 1477 3326
rect 1470 3303 1477 3306
rect 1482 3323 1501 3326
rect 1470 3246 1473 3303
rect 1470 3243 1477 3246
rect 1482 3243 1485 3323
rect 1506 3306 1509 3346
rect 1514 3333 1517 3416
rect 1522 3346 1525 3433
rect 1530 3366 1533 3476
rect 1562 3396 1565 3416
rect 1554 3393 1565 3396
rect 1530 3363 1541 3366
rect 1522 3343 1529 3346
rect 1498 3303 1509 3306
rect 1474 3226 1477 3243
rect 1474 3223 1485 3226
rect 1410 3123 1413 3213
rect 1418 3183 1421 3206
rect 1426 3143 1429 3206
rect 1386 3103 1397 3106
rect 1394 3026 1397 3103
rect 1370 2953 1377 2956
rect 1386 3023 1397 3026
rect 1350 2913 1357 2916
rect 1290 2863 1301 2866
rect 1298 2786 1301 2863
rect 1354 2836 1357 2913
rect 1354 2833 1361 2836
rect 1346 2806 1349 2826
rect 1290 2783 1301 2786
rect 1338 2803 1349 2806
rect 1238 2753 1245 2756
rect 1138 2626 1141 2646
rect 1154 2643 1165 2646
rect 1194 2683 1205 2686
rect 1106 2533 1109 2616
rect 1114 2613 1117 2626
rect 1138 2623 1145 2626
rect 1114 2566 1117 2606
rect 1114 2563 1125 2566
rect 1090 2523 1101 2526
rect 1090 2496 1093 2516
rect 1090 2493 1101 2496
rect 1082 2473 1089 2476
rect 1086 2396 1089 2473
rect 1082 2393 1089 2396
rect 1082 2353 1085 2393
rect 1098 2376 1101 2493
rect 1114 2436 1117 2556
rect 1122 2523 1125 2563
rect 1130 2543 1133 2596
rect 1142 2536 1145 2623
rect 1090 2373 1101 2376
rect 1110 2433 1117 2436
rect 1082 2313 1085 2326
rect 1074 2293 1081 2296
rect 1058 2113 1061 2126
rect 1066 2113 1069 2196
rect 1078 2156 1081 2293
rect 1074 2153 1081 2156
rect 1074 2096 1077 2153
rect 1090 2136 1093 2373
rect 1110 2276 1113 2433
rect 1122 2363 1125 2426
rect 1130 2343 1133 2536
rect 1138 2533 1145 2536
rect 1138 2513 1141 2533
rect 1154 2436 1157 2643
rect 1170 2613 1173 2626
rect 1170 2523 1173 2606
rect 1178 2593 1181 2606
rect 1194 2576 1197 2683
rect 1194 2573 1205 2576
rect 1186 2463 1189 2536
rect 1194 2523 1197 2556
rect 1150 2433 1157 2436
rect 1138 2366 1141 2406
rect 1150 2386 1153 2433
rect 1162 2413 1165 2426
rect 1178 2403 1181 2436
rect 1150 2383 1157 2386
rect 1138 2363 1149 2366
rect 1138 2333 1141 2356
rect 1146 2346 1149 2363
rect 1154 2353 1157 2383
rect 1146 2343 1157 2346
rect 1122 2286 1125 2326
rect 1130 2303 1133 2326
rect 1122 2283 1133 2286
rect 1110 2273 1117 2276
rect 1070 2093 1077 2096
rect 1082 2133 1093 2136
rect 1050 2043 1061 2046
rect 1050 2013 1053 2036
rect 1058 1946 1061 2043
rect 1070 1966 1073 2093
rect 1070 1963 1077 1966
rect 1058 1943 1065 1946
rect 1038 1883 1045 1886
rect 1018 1773 1021 1796
rect 1010 1753 1021 1756
rect 998 1743 1005 1746
rect 978 1663 989 1666
rect 954 1493 965 1496
rect 946 1393 949 1406
rect 962 1403 965 1493
rect 946 1366 949 1386
rect 978 1383 981 1663
rect 986 1613 989 1626
rect 986 1523 989 1556
rect 1002 1426 1005 1743
rect 1018 1656 1021 1753
rect 1038 1746 1041 1883
rect 1038 1743 1045 1746
rect 1010 1653 1021 1656
rect 1010 1533 1013 1653
rect 1018 1613 1021 1636
rect 1026 1613 1029 1626
rect 1034 1596 1037 1726
rect 1026 1593 1037 1596
rect 1002 1423 1013 1426
rect 994 1383 997 1416
rect 1010 1376 1013 1423
rect 1002 1373 1013 1376
rect 946 1363 957 1366
rect 954 1296 957 1363
rect 1002 1336 1005 1373
rect 1026 1346 1029 1593
rect 1026 1343 1037 1346
rect 946 1293 957 1296
rect 994 1333 1005 1336
rect 946 1246 949 1293
rect 994 1286 997 1333
rect 1018 1293 1021 1326
rect 994 1283 1005 1286
rect 942 1243 949 1246
rect 930 1213 933 1226
rect 922 1203 933 1206
rect 914 1143 925 1146
rect 906 1133 925 1136
rect 930 1133 933 1203
rect 942 1196 945 1243
rect 942 1193 949 1196
rect 946 1133 949 1193
rect 906 1106 909 1126
rect 850 1013 853 1106
rect 898 1103 909 1106
rect 898 1036 901 1103
rect 898 1033 909 1036
rect 754 973 765 976
rect 754 946 757 973
rect 754 943 765 946
rect 706 823 733 826
rect 706 813 709 823
rect 714 806 717 816
rect 690 803 717 806
rect 722 723 725 806
rect 730 706 733 823
rect 738 803 741 886
rect 746 773 749 856
rect 762 836 765 943
rect 778 913 781 926
rect 754 833 765 836
rect 726 703 733 706
rect 634 616 637 703
rect 618 596 621 616
rect 626 603 629 616
rect 634 613 645 616
rect 634 596 637 606
rect 618 593 637 596
rect 602 573 609 576
rect 558 563 565 566
rect 562 546 565 563
rect 562 543 573 546
rect 570 496 573 543
rect 586 523 589 536
rect 606 506 609 573
rect 642 556 645 613
rect 626 553 645 556
rect 618 523 621 546
rect 554 493 573 496
rect 602 503 609 506
rect 626 506 629 553
rect 634 533 637 546
rect 650 533 653 596
rect 658 533 661 626
rect 674 613 677 626
rect 714 613 717 626
rect 690 583 693 606
rect 726 556 729 703
rect 746 696 749 736
rect 706 553 729 556
rect 738 693 749 696
rect 642 513 645 526
rect 666 523 669 536
rect 682 513 685 536
rect 706 523 709 553
rect 626 503 645 506
rect 538 433 545 436
rect 490 413 493 426
rect 530 413 533 426
rect 458 396 461 406
rect 442 393 461 396
rect 506 383 509 406
rect 354 293 365 296
rect 374 333 381 336
rect 394 333 397 356
rect 410 333 413 346
rect 338 213 341 246
rect 346 213 349 256
rect 338 193 341 206
rect 354 203 357 293
rect 374 266 377 333
rect 386 296 389 326
rect 386 293 397 296
rect 374 263 381 266
rect 362 213 365 226
rect 378 213 381 263
rect 378 193 381 206
rect 386 136 389 216
rect 394 213 397 293
rect 402 286 405 326
rect 402 283 413 286
rect 402 203 405 266
rect 410 203 413 283
rect 426 213 429 246
rect 418 183 421 206
rect 386 133 397 136
rect 234 113 237 126
rect 298 113 301 126
rect 338 113 341 126
rect 394 123 397 133
rect 426 123 429 206
rect 442 203 445 336
rect 466 323 469 336
rect 514 313 517 326
rect 450 203 453 216
rect 458 203 461 236
rect 466 203 469 226
rect 474 123 477 216
rect 530 173 533 406
rect 542 366 545 433
rect 554 403 557 493
rect 602 486 605 503
rect 594 483 605 486
rect 578 413 589 416
rect 538 363 545 366
rect 538 323 541 363
rect 546 323 549 346
rect 594 326 597 483
rect 602 413 605 436
rect 642 416 645 503
rect 722 436 725 536
rect 730 533 733 546
rect 730 513 733 526
rect 738 523 741 693
rect 746 496 749 516
rect 754 503 757 833
rect 802 816 805 906
rect 810 896 813 926
rect 818 913 821 926
rect 810 893 817 896
rect 814 826 817 893
rect 814 823 821 826
rect 762 733 765 816
rect 770 813 813 816
rect 770 786 773 813
rect 778 793 781 806
rect 786 803 797 806
rect 802 803 813 806
rect 818 793 821 823
rect 770 783 797 786
rect 770 716 773 736
rect 766 713 773 716
rect 766 636 769 713
rect 766 633 773 636
rect 770 616 773 633
rect 762 613 773 616
rect 778 606 781 776
rect 786 733 789 766
rect 762 603 781 606
rect 786 603 789 616
rect 742 493 749 496
rect 722 433 733 436
rect 626 396 629 416
rect 634 403 637 416
rect 642 413 653 416
rect 642 396 645 406
rect 626 393 645 396
rect 650 386 653 413
rect 634 383 653 386
rect 602 343 621 346
rect 602 333 605 343
rect 610 326 613 336
rect 554 313 557 326
rect 570 306 573 326
rect 566 303 573 306
rect 566 246 569 303
rect 578 253 581 326
rect 594 323 613 326
rect 618 323 621 343
rect 626 333 629 346
rect 566 243 573 246
rect 570 226 573 243
rect 546 203 549 226
rect 570 223 581 226
rect 610 223 613 323
rect 506 133 509 146
rect 554 136 557 216
rect 578 176 581 223
rect 634 213 637 383
rect 658 323 661 336
rect 682 323 685 416
rect 722 403 725 416
rect 730 413 733 433
rect 742 426 745 493
rect 742 423 749 426
rect 730 403 741 406
rect 746 403 749 423
rect 754 413 757 496
rect 762 486 765 603
rect 770 533 773 556
rect 794 526 797 783
rect 802 696 805 786
rect 826 743 829 906
rect 850 813 853 936
rect 858 933 861 946
rect 866 903 869 1016
rect 874 1003 877 1016
rect 890 1013 901 1016
rect 882 993 885 1006
rect 890 976 893 1006
rect 906 1003 909 1033
rect 914 1013 917 1046
rect 886 973 893 976
rect 874 826 877 946
rect 886 846 889 973
rect 886 843 893 846
rect 858 823 877 826
rect 834 783 837 806
rect 842 793 845 806
rect 858 803 861 823
rect 866 796 869 806
rect 850 793 869 796
rect 810 713 813 726
rect 826 703 829 736
rect 802 693 813 696
rect 834 693 837 726
rect 810 626 813 693
rect 806 623 813 626
rect 806 566 809 623
rect 778 523 797 526
rect 802 563 809 566
rect 778 493 781 523
rect 762 483 781 486
rect 738 323 741 403
rect 746 333 749 346
rect 642 196 645 206
rect 650 203 653 216
rect 658 196 661 216
rect 666 203 669 226
rect 690 213 693 276
rect 674 196 677 206
rect 642 193 653 196
rect 658 193 677 196
rect 538 133 557 136
rect 570 173 581 176
rect 570 133 573 173
rect 554 113 557 126
rect 594 113 597 126
rect 650 123 653 193
rect 682 133 685 146
rect 706 123 709 216
rect 714 213 717 246
rect 714 193 717 206
rect 730 193 733 206
rect 738 203 741 216
rect 746 113 749 206
rect 754 136 757 216
rect 762 213 765 426
rect 770 333 773 366
rect 778 306 781 483
rect 794 433 797 516
rect 794 413 797 426
rect 802 413 805 563
rect 810 533 813 546
rect 794 343 797 356
rect 778 303 789 306
rect 786 236 789 303
rect 778 233 789 236
rect 810 236 813 486
rect 818 453 821 606
rect 834 556 837 616
rect 842 603 845 736
rect 850 723 853 793
rect 858 713 861 786
rect 866 706 869 746
rect 874 736 877 823
rect 882 813 885 826
rect 890 793 893 843
rect 874 733 885 736
rect 874 723 877 733
rect 850 613 853 636
rect 858 603 861 706
rect 866 703 873 706
rect 870 636 873 703
rect 866 633 873 636
rect 866 556 869 633
rect 882 623 885 726
rect 890 633 893 736
rect 898 676 901 986
rect 922 963 925 1133
rect 938 1106 941 1126
rect 934 1103 941 1106
rect 934 1036 937 1103
rect 934 1033 941 1036
rect 938 1013 941 1033
rect 906 906 909 936
rect 930 933 933 1006
rect 914 913 917 926
rect 906 903 917 906
rect 906 733 909 816
rect 914 813 917 903
rect 930 893 933 926
rect 946 856 949 1126
rect 954 1073 957 1126
rect 970 1056 973 1276
rect 1002 1236 1005 1283
rect 986 1233 1005 1236
rect 986 1186 989 1233
rect 1026 1213 1029 1326
rect 1002 1193 1005 1206
rect 986 1183 997 1186
rect 994 1083 997 1183
rect 962 1053 973 1056
rect 962 993 965 1053
rect 962 946 965 966
rect 958 943 965 946
rect 958 876 961 943
rect 958 873 965 876
rect 946 853 953 856
rect 950 776 953 853
rect 946 773 953 776
rect 906 713 909 726
rect 938 723 941 736
rect 946 716 949 773
rect 962 746 965 873
rect 970 813 973 926
rect 978 913 981 936
rect 994 766 997 996
rect 1002 976 1005 1136
rect 1018 1103 1021 1126
rect 1010 1013 1013 1026
rect 1002 973 1021 976
rect 1010 943 1013 956
rect 1018 926 1021 973
rect 1010 923 1021 926
rect 1010 846 1013 923
rect 1026 856 1029 1086
rect 1034 933 1037 1343
rect 1042 986 1045 1743
rect 1050 1403 1053 1936
rect 1062 1746 1065 1943
rect 1074 1906 1077 1963
rect 1082 1923 1085 2133
rect 1090 2083 1093 2126
rect 1098 1993 1101 2106
rect 1106 1976 1109 2206
rect 1114 2116 1117 2273
rect 1130 2226 1133 2283
rect 1122 2223 1133 2226
rect 1122 2133 1125 2223
rect 1146 2203 1149 2336
rect 1154 2323 1157 2343
rect 1162 2333 1165 2376
rect 1154 2186 1157 2226
rect 1146 2183 1157 2186
rect 1114 2113 1121 2116
rect 1098 1973 1109 1976
rect 1074 1903 1085 1906
rect 1082 1826 1085 1903
rect 1058 1743 1065 1746
rect 1074 1823 1085 1826
rect 1098 1826 1101 1973
rect 1118 1966 1121 2113
rect 1146 2106 1149 2183
rect 1162 2106 1165 2256
rect 1170 2213 1173 2346
rect 1178 2313 1181 2326
rect 1194 2306 1197 2326
rect 1190 2303 1197 2306
rect 1190 2236 1193 2303
rect 1190 2233 1197 2236
rect 1178 2123 1181 2216
rect 1194 2213 1197 2233
rect 1202 2213 1205 2573
rect 1210 2523 1213 2706
rect 1242 2686 1245 2753
rect 1238 2683 1245 2686
rect 1226 2523 1229 2676
rect 1238 2466 1241 2683
rect 1254 2676 1257 2763
rect 1266 2723 1269 2736
rect 1250 2673 1257 2676
rect 1210 2413 1213 2426
rect 1210 2223 1213 2356
rect 1218 2306 1221 2466
rect 1238 2463 1245 2466
rect 1226 2323 1229 2336
rect 1218 2303 1225 2306
rect 1222 2236 1225 2303
rect 1218 2233 1225 2236
rect 1194 2203 1205 2206
rect 1202 2186 1205 2203
rect 1210 2193 1213 2206
rect 1202 2183 1213 2186
rect 1146 2103 1157 2106
rect 1162 2103 1181 2106
rect 1130 2003 1133 2086
rect 1114 1963 1121 1966
rect 1114 1946 1117 1963
rect 1110 1943 1117 1946
rect 1110 1896 1113 1943
rect 1122 1906 1125 1936
rect 1138 1923 1141 2006
rect 1122 1903 1133 1906
rect 1110 1893 1117 1896
rect 1098 1823 1109 1826
rect 1058 1696 1061 1743
rect 1074 1733 1077 1823
rect 1082 1733 1085 1756
rect 1066 1713 1069 1726
rect 1058 1693 1065 1696
rect 1062 1546 1065 1693
rect 1074 1673 1077 1726
rect 1090 1723 1093 1806
rect 1106 1743 1109 1823
rect 1098 1706 1101 1736
rect 1090 1703 1101 1706
rect 1090 1636 1093 1703
rect 1058 1543 1065 1546
rect 1074 1633 1093 1636
rect 1058 1496 1061 1543
rect 1066 1513 1069 1526
rect 1058 1493 1065 1496
rect 1062 1396 1065 1493
rect 1058 1393 1065 1396
rect 1058 1356 1061 1393
rect 1058 1353 1065 1356
rect 1050 1203 1053 1346
rect 1062 1256 1065 1353
rect 1062 1253 1069 1256
rect 1050 1123 1053 1146
rect 1066 1133 1069 1253
rect 1050 1006 1053 1096
rect 1058 1023 1061 1126
rect 1066 1103 1069 1126
rect 1050 1003 1061 1006
rect 1042 983 1049 986
rect 1046 926 1049 983
rect 1042 923 1049 926
rect 1026 853 1033 856
rect 1010 843 1021 846
rect 1010 793 1013 806
rect 938 713 949 716
rect 958 743 965 746
rect 986 763 997 766
rect 898 673 917 676
rect 914 566 917 673
rect 938 656 941 713
rect 958 696 961 743
rect 986 706 989 763
rect 1010 743 1013 756
rect 1018 726 1021 843
rect 1030 786 1033 853
rect 1026 783 1033 786
rect 1026 733 1029 783
rect 1034 743 1037 766
rect 1018 723 1029 726
rect 986 703 1005 706
rect 958 693 965 696
rect 930 653 941 656
rect 930 576 933 653
rect 954 613 957 626
rect 962 583 965 693
rect 930 573 949 576
rect 898 563 917 566
rect 834 553 861 556
rect 866 553 877 556
rect 826 543 845 546
rect 826 523 829 543
rect 818 333 821 346
rect 810 233 821 236
rect 770 183 773 206
rect 778 203 781 233
rect 810 203 813 216
rect 818 203 821 233
rect 826 203 829 506
rect 834 423 837 536
rect 842 533 845 543
rect 842 503 845 526
rect 834 333 837 416
rect 786 193 797 196
rect 826 183 829 196
rect 754 133 765 136
rect 762 123 765 133
rect 770 123 773 176
rect 802 133 805 146
rect 810 143 829 146
rect 842 143 845 456
rect 850 413 853 526
rect 858 493 861 553
rect 866 533 869 546
rect 866 503 869 526
rect 874 523 877 553
rect 890 413 893 536
rect 898 483 901 563
rect 922 543 941 546
rect 922 523 925 543
rect 874 393 877 406
rect 858 283 861 326
rect 866 243 869 326
rect 882 313 885 326
rect 850 213 853 226
rect 882 213 885 236
rect 890 213 893 346
rect 898 296 901 326
rect 906 313 909 336
rect 914 323 917 506
rect 930 453 933 536
rect 938 533 941 543
rect 946 333 949 573
rect 954 523 957 536
rect 962 413 965 526
rect 978 523 981 546
rect 1002 516 1005 703
rect 1026 646 1029 723
rect 1026 643 1033 646
rect 986 513 1005 516
rect 898 293 909 296
rect 906 226 909 293
rect 898 223 909 226
rect 794 93 797 126
rect 810 123 813 143
rect 818 113 821 136
rect 826 133 829 143
rect 842 123 845 136
rect 898 133 901 223
rect 946 213 949 326
rect 954 263 957 346
rect 970 333 973 346
rect 986 326 989 513
rect 1002 363 1005 396
rect 1010 333 1013 586
rect 1018 573 1021 596
rect 1030 576 1033 643
rect 1030 573 1037 576
rect 1018 533 1021 546
rect 1026 543 1029 556
rect 1034 536 1037 573
rect 1042 543 1045 923
rect 1058 836 1061 1003
rect 1050 833 1061 836
rect 1050 803 1053 833
rect 1050 723 1053 746
rect 1050 603 1053 716
rect 1058 653 1061 816
rect 1066 803 1069 816
rect 1066 733 1069 796
rect 1074 713 1077 1633
rect 1082 1386 1085 1506
rect 1090 1433 1093 1626
rect 1106 1583 1109 1726
rect 1114 1476 1117 1893
rect 1130 1836 1133 1903
rect 1122 1833 1133 1836
rect 1122 1756 1125 1833
rect 1130 1803 1133 1816
rect 1146 1813 1149 1836
rect 1130 1776 1133 1796
rect 1130 1773 1141 1776
rect 1122 1753 1129 1756
rect 1126 1676 1129 1753
rect 1122 1673 1129 1676
rect 1122 1586 1125 1673
rect 1138 1656 1141 1773
rect 1130 1653 1141 1656
rect 1130 1623 1133 1653
rect 1130 1596 1133 1606
rect 1138 1603 1141 1636
rect 1146 1596 1149 1616
rect 1154 1613 1157 2103
rect 1178 1946 1181 2103
rect 1162 1943 1181 1946
rect 1162 1926 1165 1943
rect 1202 1926 1205 2176
rect 1210 2153 1213 2183
rect 1218 2136 1221 2233
rect 1214 2133 1221 2136
rect 1214 1956 1217 2133
rect 1226 1966 1229 2216
rect 1234 2123 1237 2336
rect 1242 2106 1245 2463
rect 1250 2356 1253 2673
rect 1258 2603 1261 2626
rect 1266 2593 1269 2626
rect 1282 2613 1285 2626
rect 1282 2543 1285 2606
rect 1258 2373 1261 2536
rect 1282 2513 1285 2526
rect 1250 2353 1257 2356
rect 1254 2236 1257 2353
rect 1266 2256 1269 2506
rect 1290 2483 1293 2783
rect 1298 2746 1301 2766
rect 1338 2756 1341 2803
rect 1338 2753 1349 2756
rect 1298 2743 1309 2746
rect 1306 2586 1309 2743
rect 1338 2723 1341 2736
rect 1346 2723 1349 2753
rect 1358 2716 1361 2833
rect 1354 2713 1361 2716
rect 1322 2603 1325 2646
rect 1330 2613 1333 2626
rect 1346 2613 1349 2626
rect 1330 2593 1333 2606
rect 1298 2583 1309 2586
rect 1298 2466 1301 2583
rect 1354 2576 1357 2713
rect 1346 2573 1357 2576
rect 1306 2513 1309 2546
rect 1314 2533 1317 2566
rect 1294 2463 1301 2466
rect 1274 2383 1277 2406
rect 1266 2253 1277 2256
rect 1254 2233 1261 2236
rect 1258 2166 1261 2233
rect 1274 2173 1277 2253
rect 1282 2223 1285 2426
rect 1294 2266 1297 2463
rect 1294 2263 1301 2266
rect 1238 2103 1245 2106
rect 1250 2163 1261 2166
rect 1282 2163 1285 2216
rect 1238 1986 1241 2103
rect 1250 1996 1253 2163
rect 1258 2133 1261 2146
rect 1258 2013 1261 2026
rect 1266 2003 1269 2126
rect 1274 2116 1277 2156
rect 1282 2133 1285 2146
rect 1274 2113 1281 2116
rect 1278 2006 1281 2113
rect 1274 2003 1281 2006
rect 1250 1993 1257 1996
rect 1238 1983 1245 1986
rect 1226 1963 1233 1966
rect 1214 1953 1221 1956
rect 1162 1923 1173 1926
rect 1194 1923 1205 1926
rect 1194 1866 1197 1923
rect 1194 1863 1205 1866
rect 1170 1793 1173 1846
rect 1194 1813 1197 1836
rect 1162 1613 1165 1646
rect 1130 1593 1149 1596
rect 1122 1583 1137 1586
rect 1106 1473 1117 1476
rect 1090 1403 1093 1416
rect 1106 1406 1109 1473
rect 1122 1413 1125 1526
rect 1134 1446 1137 1583
rect 1154 1576 1157 1596
rect 1154 1573 1161 1576
rect 1134 1443 1141 1446
rect 1130 1413 1133 1426
rect 1106 1403 1117 1406
rect 1082 1383 1093 1386
rect 1090 1216 1093 1383
rect 1114 1216 1117 1403
rect 1138 1396 1141 1443
rect 1130 1393 1141 1396
rect 1130 1246 1133 1393
rect 1130 1243 1141 1246
rect 1082 1213 1093 1216
rect 1106 1213 1117 1216
rect 1130 1213 1133 1226
rect 1082 1103 1085 1213
rect 1090 1173 1093 1196
rect 1106 1156 1109 1213
rect 1106 1153 1117 1156
rect 1090 1133 1109 1136
rect 1082 993 1085 1016
rect 1090 1013 1093 1046
rect 1098 903 1101 1126
rect 1106 1013 1109 1133
rect 1114 1093 1117 1153
rect 1122 1113 1125 1206
rect 1138 1203 1141 1243
rect 1146 1196 1149 1486
rect 1158 1446 1161 1573
rect 1154 1443 1161 1446
rect 1154 1393 1157 1443
rect 1162 1403 1165 1426
rect 1162 1326 1165 1396
rect 1138 1193 1149 1196
rect 1158 1323 1165 1326
rect 1122 993 1125 1006
rect 1138 1003 1141 1193
rect 1158 1156 1161 1323
rect 1158 1153 1165 1156
rect 1162 1136 1165 1153
rect 1146 1123 1149 1136
rect 1154 1133 1165 1136
rect 1170 1133 1173 1746
rect 1178 1706 1181 1736
rect 1186 1723 1189 1796
rect 1194 1733 1197 1746
rect 1202 1723 1205 1863
rect 1178 1703 1189 1706
rect 1186 1506 1189 1703
rect 1210 1656 1213 1936
rect 1218 1733 1221 1953
rect 1230 1856 1233 1963
rect 1242 1923 1245 1983
rect 1254 1916 1257 1993
rect 1274 1983 1277 2003
rect 1290 1966 1293 2246
rect 1298 2226 1301 2263
rect 1306 2243 1309 2486
rect 1322 2306 1325 2526
rect 1346 2326 1349 2573
rect 1362 2533 1365 2546
rect 1362 2333 1365 2356
rect 1346 2323 1357 2326
rect 1322 2303 1333 2306
rect 1330 2246 1333 2303
rect 1354 2276 1357 2323
rect 1322 2243 1333 2246
rect 1346 2273 1357 2276
rect 1370 2276 1373 2953
rect 1386 2946 1389 3023
rect 1418 3013 1421 3136
rect 1410 3003 1421 3006
rect 1426 2986 1429 3046
rect 1418 2983 1429 2986
rect 1386 2943 1397 2946
rect 1378 2823 1381 2936
rect 1386 2896 1389 2936
rect 1394 2923 1397 2943
rect 1402 2903 1405 2936
rect 1386 2893 1393 2896
rect 1390 2816 1393 2893
rect 1386 2813 1393 2816
rect 1386 2716 1389 2813
rect 1402 2773 1405 2896
rect 1418 2886 1421 2983
rect 1434 2966 1437 3166
rect 1442 3076 1445 3206
rect 1450 3123 1453 3156
rect 1466 3076 1469 3196
rect 1442 3073 1453 3076
rect 1450 3013 1453 3073
rect 1462 3073 1469 3076
rect 1462 2996 1465 3073
rect 1482 3066 1485 3223
rect 1498 3166 1501 3303
rect 1514 3286 1517 3326
rect 1510 3283 1517 3286
rect 1510 3186 1513 3283
rect 1526 3276 1529 3343
rect 1522 3273 1529 3276
rect 1510 3183 1517 3186
rect 1498 3163 1509 3166
rect 1506 3093 1509 3163
rect 1430 2963 1437 2966
rect 1458 2993 1465 2996
rect 1474 3063 1485 3066
rect 1430 2906 1433 2963
rect 1442 2906 1445 2956
rect 1458 2926 1461 2993
rect 1458 2923 1469 2926
rect 1430 2903 1437 2906
rect 1442 2903 1453 2906
rect 1418 2883 1429 2886
rect 1378 2713 1389 2716
rect 1386 2626 1389 2713
rect 1402 2626 1405 2726
rect 1378 2623 1389 2626
rect 1386 2413 1389 2623
rect 1394 2623 1405 2626
rect 1394 2613 1397 2623
rect 1402 2523 1405 2623
rect 1410 2596 1413 2866
rect 1418 2733 1421 2836
rect 1418 2613 1421 2706
rect 1426 2686 1429 2883
rect 1434 2706 1437 2903
rect 1450 2846 1453 2903
rect 1466 2863 1469 2923
rect 1442 2843 1453 2846
rect 1442 2723 1445 2843
rect 1458 2813 1461 2826
rect 1450 2723 1453 2806
rect 1466 2786 1469 2806
rect 1458 2783 1469 2786
rect 1458 2733 1461 2783
rect 1466 2706 1469 2776
rect 1434 2703 1445 2706
rect 1426 2683 1433 2686
rect 1430 2606 1433 2683
rect 1426 2603 1433 2606
rect 1410 2593 1417 2596
rect 1414 2516 1417 2593
rect 1410 2513 1417 2516
rect 1402 2413 1405 2436
rect 1378 2383 1381 2406
rect 1386 2363 1389 2406
rect 1410 2346 1413 2513
rect 1410 2343 1417 2346
rect 1386 2323 1389 2336
rect 1414 2296 1417 2343
rect 1410 2293 1417 2296
rect 1370 2273 1381 2276
rect 1298 2223 1309 2226
rect 1306 2146 1309 2223
rect 1322 2213 1325 2243
rect 1346 2216 1349 2273
rect 1362 2223 1365 2266
rect 1346 2213 1357 2216
rect 1298 2143 1309 2146
rect 1298 2056 1301 2143
rect 1306 2073 1309 2126
rect 1298 2053 1309 2056
rect 1306 1966 1309 2053
rect 1282 1963 1293 1966
rect 1298 1963 1309 1966
rect 1250 1913 1257 1916
rect 1230 1853 1237 1856
rect 1234 1836 1237 1853
rect 1234 1833 1241 1836
rect 1238 1776 1241 1833
rect 1234 1773 1241 1776
rect 1226 1733 1229 1766
rect 1218 1723 1229 1726
rect 1226 1703 1229 1723
rect 1234 1686 1237 1773
rect 1202 1653 1213 1656
rect 1230 1683 1237 1686
rect 1202 1606 1205 1653
rect 1202 1603 1213 1606
rect 1202 1523 1205 1586
rect 1178 1503 1189 1506
rect 1210 1503 1213 1603
rect 1218 1536 1221 1646
rect 1230 1586 1233 1683
rect 1242 1643 1245 1756
rect 1250 1726 1253 1913
rect 1266 1826 1269 1936
rect 1282 1866 1285 1963
rect 1282 1863 1293 1866
rect 1290 1843 1293 1863
rect 1298 1826 1301 1963
rect 1330 1933 1333 2186
rect 1354 2026 1357 2213
rect 1378 2186 1381 2273
rect 1402 2193 1405 2206
rect 1346 2023 1357 2026
rect 1370 2183 1381 2186
rect 1346 1976 1349 2023
rect 1346 1973 1357 1976
rect 1266 1823 1273 1826
rect 1258 1743 1261 1816
rect 1270 1776 1273 1823
rect 1294 1823 1301 1826
rect 1266 1773 1273 1776
rect 1266 1753 1269 1773
rect 1250 1723 1257 1726
rect 1254 1636 1257 1723
rect 1242 1603 1245 1636
rect 1250 1633 1257 1636
rect 1230 1583 1237 1586
rect 1234 1563 1237 1583
rect 1250 1573 1253 1633
rect 1258 1603 1261 1616
rect 1266 1603 1269 1716
rect 1218 1533 1229 1536
rect 1234 1533 1237 1546
rect 1242 1533 1253 1536
rect 1258 1533 1261 1546
rect 1226 1526 1229 1533
rect 1178 1483 1181 1503
rect 1178 1333 1181 1416
rect 1186 1413 1189 1446
rect 1194 1413 1205 1416
rect 1218 1413 1221 1526
rect 1226 1523 1237 1526
rect 1186 1296 1189 1316
rect 1182 1293 1189 1296
rect 1182 1226 1185 1293
rect 1182 1223 1189 1226
rect 1178 1133 1181 1206
rect 1162 1123 1173 1126
rect 1154 1036 1157 1116
rect 1178 1086 1181 1106
rect 1174 1083 1181 1086
rect 1154 1033 1165 1036
rect 1106 913 1109 926
rect 1114 893 1117 986
rect 1130 973 1133 996
rect 1082 813 1085 826
rect 1122 813 1125 826
rect 1130 813 1133 926
rect 1146 893 1149 1026
rect 1162 956 1165 1033
rect 1154 953 1165 956
rect 1154 886 1157 953
rect 1162 923 1165 936
rect 1146 883 1157 886
rect 1162 883 1165 916
rect 1146 866 1149 883
rect 1174 866 1177 1083
rect 1186 1023 1189 1223
rect 1194 1146 1197 1396
rect 1202 1166 1205 1356
rect 1210 1223 1213 1406
rect 1218 1316 1221 1366
rect 1226 1333 1229 1506
rect 1234 1333 1237 1523
rect 1242 1423 1245 1526
rect 1250 1523 1261 1526
rect 1242 1353 1245 1416
rect 1258 1343 1261 1436
rect 1266 1363 1269 1566
rect 1282 1416 1285 1776
rect 1294 1696 1297 1823
rect 1306 1813 1317 1816
rect 1306 1773 1309 1813
rect 1322 1803 1325 1896
rect 1338 1766 1341 1846
rect 1346 1783 1349 1816
rect 1354 1793 1357 1973
rect 1362 1923 1365 2016
rect 1370 1906 1373 2183
rect 1410 2176 1413 2293
rect 1406 2173 1413 2176
rect 1378 2046 1381 2166
rect 1386 2103 1389 2136
rect 1394 2063 1397 2126
rect 1406 2046 1409 2173
rect 1418 2113 1421 2206
rect 1378 2043 1389 2046
rect 1386 1976 1389 2043
rect 1366 1903 1373 1906
rect 1378 1973 1389 1976
rect 1402 2043 1409 2046
rect 1366 1776 1369 1903
rect 1362 1773 1369 1776
rect 1338 1763 1349 1766
rect 1322 1736 1325 1756
rect 1322 1733 1333 1736
rect 1306 1703 1309 1726
rect 1294 1693 1301 1696
rect 1290 1523 1293 1546
rect 1298 1506 1301 1693
rect 1322 1683 1325 1726
rect 1346 1676 1349 1763
rect 1362 1706 1365 1773
rect 1362 1703 1373 1706
rect 1370 1683 1373 1703
rect 1338 1673 1349 1676
rect 1322 1603 1325 1616
rect 1330 1603 1333 1616
rect 1322 1533 1325 1556
rect 1306 1523 1317 1526
rect 1338 1523 1341 1673
rect 1346 1613 1349 1626
rect 1354 1613 1357 1636
rect 1354 1596 1357 1606
rect 1362 1603 1365 1616
rect 1370 1596 1373 1616
rect 1354 1593 1373 1596
rect 1378 1576 1381 1973
rect 1402 1916 1405 2043
rect 1418 2026 1421 2106
rect 1414 2023 1421 2026
rect 1414 1946 1417 2023
rect 1414 1943 1421 1946
rect 1418 1923 1421 1943
rect 1402 1913 1413 1916
rect 1394 1776 1397 1806
rect 1394 1773 1405 1776
rect 1394 1733 1397 1746
rect 1402 1733 1405 1773
rect 1410 1726 1413 1913
rect 1426 1866 1429 2603
rect 1442 2566 1445 2703
rect 1434 2563 1445 2566
rect 1458 2703 1469 2706
rect 1458 2566 1461 2703
rect 1458 2563 1465 2566
rect 1434 2463 1437 2563
rect 1450 2533 1453 2546
rect 1462 2476 1465 2563
rect 1474 2483 1477 3063
rect 1482 2896 1485 2996
rect 1498 2976 1501 3016
rect 1514 3003 1517 3183
rect 1522 3106 1525 3273
rect 1538 3226 1541 3363
rect 1554 3346 1557 3393
rect 1554 3343 1565 3346
rect 1554 3306 1557 3326
rect 1550 3303 1557 3306
rect 1550 3236 1553 3303
rect 1550 3233 1557 3236
rect 1530 3223 1541 3226
rect 1530 3163 1533 3223
rect 1538 3133 1541 3206
rect 1546 3176 1549 3206
rect 1554 3183 1557 3233
rect 1562 3203 1565 3343
rect 1570 3323 1573 3513
rect 1602 3473 1605 3536
rect 1610 3503 1613 3536
rect 1594 3393 1597 3406
rect 1578 3333 1581 3346
rect 1594 3316 1597 3376
rect 1594 3313 1601 3316
rect 1578 3213 1581 3296
rect 1578 3183 1581 3206
rect 1586 3203 1589 3306
rect 1598 3236 1601 3313
rect 1594 3233 1601 3236
rect 1546 3173 1557 3176
rect 1546 3133 1549 3156
rect 1554 3133 1557 3173
rect 1578 3136 1581 3146
rect 1570 3133 1581 3136
rect 1586 3133 1589 3166
rect 1546 3123 1565 3126
rect 1522 3103 1533 3106
rect 1530 3036 1533 3103
rect 1522 3033 1533 3036
rect 1522 2993 1525 3033
rect 1498 2973 1509 2976
rect 1490 2933 1493 2946
rect 1506 2933 1509 2973
rect 1482 2893 1493 2896
rect 1490 2826 1493 2893
rect 1482 2823 1493 2826
rect 1482 2803 1485 2823
rect 1506 2816 1509 2926
rect 1506 2813 1525 2816
rect 1546 2813 1549 3016
rect 1562 3013 1565 3026
rect 1578 3023 1581 3126
rect 1594 3116 1597 3233
rect 1602 3123 1605 3216
rect 1590 3113 1597 3116
rect 1590 3036 1593 3113
rect 1610 3103 1613 3366
rect 1618 3183 1621 3543
rect 1626 3533 1629 3546
rect 1658 3543 1661 3616
rect 1634 3523 1637 3536
rect 1642 3526 1645 3536
rect 1642 3523 1653 3526
rect 1626 3276 1629 3396
rect 1634 3313 1637 3426
rect 1642 3333 1645 3406
rect 1658 3393 1661 3406
rect 1682 3403 1685 3416
rect 1666 3336 1669 3366
rect 1690 3363 1693 3576
rect 1722 3533 1725 3576
rect 1714 3456 1717 3526
rect 1714 3453 1725 3456
rect 1698 3346 1701 3406
rect 1690 3343 1701 3346
rect 1666 3333 1677 3336
rect 1650 3293 1653 3326
rect 1674 3286 1677 3333
rect 1666 3283 1677 3286
rect 1626 3273 1637 3276
rect 1634 3176 1637 3273
rect 1626 3173 1637 3176
rect 1590 3033 1597 3036
rect 1554 2923 1557 2936
rect 1578 2933 1581 3006
rect 1586 2943 1589 3016
rect 1594 2926 1597 3033
rect 1590 2923 1597 2926
rect 1590 2856 1593 2923
rect 1590 2853 1597 2856
rect 1482 2703 1485 2726
rect 1490 2623 1493 2736
rect 1498 2723 1501 2806
rect 1522 2716 1525 2813
rect 1570 2726 1573 2806
rect 1594 2786 1597 2853
rect 1590 2783 1597 2786
rect 1506 2713 1525 2716
rect 1562 2723 1573 2726
rect 1506 2666 1509 2713
rect 1498 2663 1509 2666
rect 1562 2666 1565 2723
rect 1578 2676 1581 2726
rect 1590 2716 1593 2783
rect 1602 2723 1605 3096
rect 1610 2996 1613 3016
rect 1626 3013 1629 3173
rect 1650 3123 1653 3146
rect 1610 2993 1617 2996
rect 1614 2846 1617 2993
rect 1626 2923 1629 2946
rect 1610 2843 1617 2846
rect 1610 2743 1613 2843
rect 1618 2813 1621 2826
rect 1626 2733 1629 2776
rect 1642 2756 1645 3036
rect 1666 3033 1669 3283
rect 1690 3276 1693 3343
rect 1706 3286 1709 3446
rect 1722 3403 1725 3453
rect 1714 3333 1717 3346
rect 1706 3283 1713 3286
rect 1690 3273 1701 3276
rect 1690 3203 1693 3256
rect 1658 2813 1661 2936
rect 1666 2923 1669 3016
rect 1682 3013 1685 3026
rect 1674 2823 1677 3006
rect 1682 2933 1685 2976
rect 1638 2753 1645 2756
rect 1590 2713 1597 2716
rect 1578 2673 1585 2676
rect 1562 2663 1573 2666
rect 1462 2473 1469 2476
rect 1434 2323 1437 2346
rect 1434 2173 1437 2226
rect 1434 2116 1437 2136
rect 1434 2113 1441 2116
rect 1438 2046 1441 2113
rect 1450 2083 1453 2436
rect 1466 2186 1469 2473
rect 1482 2403 1485 2526
rect 1490 2306 1493 2326
rect 1482 2303 1493 2306
rect 1482 2246 1485 2303
rect 1498 2256 1501 2663
rect 1570 2636 1573 2663
rect 1562 2633 1573 2636
rect 1514 2613 1517 2626
rect 1562 2576 1565 2633
rect 1582 2626 1585 2673
rect 1578 2623 1585 2626
rect 1578 2603 1581 2623
rect 1562 2573 1573 2576
rect 1514 2426 1517 2486
rect 1510 2423 1517 2426
rect 1510 2276 1513 2423
rect 1522 2413 1541 2416
rect 1510 2273 1517 2276
rect 1498 2253 1505 2256
rect 1482 2243 1493 2246
rect 1482 2203 1485 2226
rect 1490 2203 1493 2243
rect 1502 2196 1505 2253
rect 1498 2193 1505 2196
rect 1466 2183 1477 2186
rect 1474 2076 1477 2183
rect 1434 2043 1441 2046
rect 1466 2073 1477 2076
rect 1434 2023 1437 2043
rect 1434 1923 1437 1986
rect 1466 1946 1469 2073
rect 1498 2016 1501 2193
rect 1514 2133 1517 2273
rect 1522 2116 1525 2366
rect 1530 2203 1533 2406
rect 1546 2403 1549 2526
rect 1570 2433 1573 2573
rect 1586 2466 1589 2536
rect 1578 2463 1589 2466
rect 1538 2213 1541 2386
rect 1546 2333 1549 2346
rect 1554 2323 1557 2416
rect 1578 2373 1581 2463
rect 1586 2403 1589 2456
rect 1594 2336 1597 2713
rect 1610 2613 1613 2646
rect 1602 2533 1605 2606
rect 1610 2526 1613 2576
rect 1618 2543 1621 2606
rect 1626 2533 1629 2726
rect 1638 2696 1641 2753
rect 1658 2733 1661 2746
rect 1682 2723 1685 2806
rect 1690 2706 1693 3186
rect 1698 3106 1701 3273
rect 1710 3236 1713 3283
rect 1706 3233 1713 3236
rect 1706 3183 1709 3233
rect 1714 3196 1717 3216
rect 1722 3213 1725 3326
rect 1714 3193 1721 3196
rect 1706 3123 1709 3156
rect 1718 3116 1721 3193
rect 1714 3113 1721 3116
rect 1698 3103 1705 3106
rect 1702 2986 1705 3103
rect 1714 3013 1717 3113
rect 1722 3003 1725 3076
rect 1730 2986 1733 3916
rect 1746 3836 1749 3933
rect 1758 3876 1761 3953
rect 1770 3886 1773 4033
rect 1786 3903 1789 4016
rect 1794 3993 1797 4006
rect 1802 3923 1805 3956
rect 1770 3883 1781 3886
rect 1758 3873 1765 3876
rect 1738 3833 1749 3836
rect 1738 3706 1741 3833
rect 1746 3813 1749 3826
rect 1754 3806 1757 3816
rect 1746 3803 1757 3806
rect 1746 3723 1749 3803
rect 1762 3743 1765 3873
rect 1778 3816 1781 3883
rect 1810 3846 1813 4033
rect 1818 4013 1821 4026
rect 1834 4003 1837 4056
rect 1858 4013 1861 4026
rect 1818 3923 1821 3996
rect 1818 3896 1821 3916
rect 1818 3893 1825 3896
rect 1806 3843 1813 3846
rect 1770 3813 1781 3816
rect 1770 3773 1773 3813
rect 1778 3723 1781 3796
rect 1794 3733 1797 3816
rect 1806 3746 1809 3843
rect 1822 3836 1825 3893
rect 1818 3833 1825 3836
rect 1806 3743 1813 3746
rect 1786 3713 1789 3726
rect 1738 3703 1745 3706
rect 1742 3636 1745 3703
rect 1738 3633 1745 3636
rect 1738 3506 1741 3633
rect 1794 3626 1797 3646
rect 1790 3623 1797 3626
rect 1746 3523 1749 3616
rect 1762 3533 1765 3586
rect 1738 3503 1745 3506
rect 1742 3436 1745 3503
rect 1754 3493 1757 3526
rect 1770 3443 1773 3616
rect 1790 3576 1793 3623
rect 1802 3583 1805 3726
rect 1810 3663 1813 3743
rect 1818 3603 1821 3833
rect 1826 3796 1829 3806
rect 1834 3803 1837 3866
rect 1850 3816 1853 3926
rect 1842 3796 1845 3816
rect 1850 3813 1861 3816
rect 1826 3793 1845 3796
rect 1850 3793 1853 3806
rect 1866 3796 1869 4066
rect 1882 4016 1885 4036
rect 1878 4013 1885 4016
rect 1878 3936 1881 4013
rect 1898 3956 1901 4126
rect 1906 4123 1917 4126
rect 1914 4036 1917 4123
rect 1890 3953 1901 3956
rect 1906 4033 1917 4036
rect 1878 3933 1885 3936
rect 1882 3913 1885 3933
rect 1890 3923 1893 3953
rect 1898 3933 1901 3946
rect 1906 3906 1909 4033
rect 1938 4026 1941 4273
rect 1946 4213 1949 4306
rect 1978 4303 1989 4306
rect 1994 4303 1997 4326
rect 1986 4213 1989 4303
rect 1978 4193 1981 4206
rect 1954 4063 1957 4156
rect 1978 4133 1981 4146
rect 1986 4123 1989 4166
rect 2002 4036 2005 4326
rect 2018 4203 2021 4346
rect 2026 4323 2029 4406
rect 2034 4393 2037 4616
rect 2050 4583 2053 4606
rect 2050 4533 2061 4536
rect 2042 4513 2045 4526
rect 2066 4523 2069 4536
rect 2074 4523 2077 4616
rect 2082 4463 2085 4526
rect 2130 4523 2133 4536
rect 2138 4533 2141 4616
rect 2170 4613 2173 4626
rect 2210 4613 2213 4626
rect 2162 4543 2165 4606
rect 2186 4593 2189 4606
rect 2162 4533 2181 4536
rect 2146 4513 2149 4526
rect 2154 4483 2157 4526
rect 2162 4523 2173 4526
rect 2034 4306 2037 4366
rect 2042 4323 2045 4406
rect 2066 4403 2069 4416
rect 2114 4386 2117 4406
rect 2138 4386 2141 4406
rect 2114 4383 2141 4386
rect 2050 4323 2053 4346
rect 2034 4303 2045 4306
rect 2082 4303 2085 4326
rect 2042 4226 2045 4303
rect 2034 4223 2045 4226
rect 2034 4193 2037 4223
rect 2130 4216 2133 4383
rect 2162 4323 2165 4416
rect 2170 4306 2173 4486
rect 2178 4363 2181 4533
rect 2194 4523 2197 4536
rect 2226 4533 2229 4546
rect 2234 4533 2237 4566
rect 2210 4426 2213 4526
rect 2242 4446 2245 4526
rect 2162 4303 2173 4306
rect 2162 4236 2165 4303
rect 2162 4233 2173 4236
rect 2170 4216 2173 4233
rect 2122 4213 2133 4216
rect 2042 4133 2045 4156
rect 2050 4123 2053 4206
rect 1930 4023 1941 4026
rect 1994 4033 2005 4036
rect 1914 3943 1917 4016
rect 1930 3956 1933 4023
rect 1930 3953 1941 3956
rect 1922 3933 1933 3936
rect 1898 3903 1909 3906
rect 1898 3836 1901 3903
rect 1914 3883 1917 3926
rect 1898 3833 1909 3836
rect 1862 3793 1869 3796
rect 1826 3756 1829 3776
rect 1826 3753 1837 3756
rect 1834 3696 1837 3753
rect 1826 3693 1837 3696
rect 1778 3533 1781 3576
rect 1790 3573 1797 3576
rect 1778 3523 1789 3526
rect 1794 3516 1797 3573
rect 1786 3513 1797 3516
rect 1738 3433 1745 3436
rect 1738 3386 1741 3433
rect 1746 3406 1749 3416
rect 1754 3413 1757 3426
rect 1746 3403 1765 3406
rect 1770 3386 1773 3416
rect 1738 3383 1749 3386
rect 1746 3296 1749 3383
rect 1762 3383 1773 3386
rect 1762 3306 1765 3383
rect 1778 3313 1781 3496
rect 1786 3403 1789 3513
rect 1802 3496 1805 3526
rect 1798 3493 1805 3496
rect 1798 3436 1801 3493
rect 1798 3433 1805 3436
rect 1794 3366 1797 3416
rect 1786 3363 1797 3366
rect 1762 3303 1773 3306
rect 1738 3293 1749 3296
rect 1738 3186 1741 3293
rect 1746 3203 1749 3276
rect 1770 3256 1773 3303
rect 1762 3253 1773 3256
rect 1738 3183 1749 3186
rect 1746 3036 1749 3183
rect 1702 2983 1709 2986
rect 1706 2856 1709 2983
rect 1686 2703 1693 2706
rect 1698 2853 1709 2856
rect 1722 2983 1733 2986
rect 1738 3033 1749 3036
rect 1638 2693 1645 2696
rect 1642 2676 1645 2693
rect 1642 2673 1653 2676
rect 1634 2613 1637 2646
rect 1634 2593 1637 2606
rect 1650 2596 1653 2673
rect 1686 2626 1689 2703
rect 1686 2623 1693 2626
rect 1650 2593 1661 2596
rect 1658 2576 1661 2593
rect 1650 2573 1661 2576
rect 1602 2413 1605 2526
rect 1610 2523 1617 2526
rect 1614 2446 1617 2523
rect 1650 2516 1653 2573
rect 1674 2523 1677 2606
rect 1650 2513 1661 2516
rect 1610 2443 1617 2446
rect 1610 2383 1613 2443
rect 1626 2403 1629 2436
rect 1658 2426 1661 2513
rect 1682 2493 1685 2606
rect 1690 2563 1693 2623
rect 1698 2546 1701 2853
rect 1722 2836 1725 2983
rect 1738 2966 1741 3033
rect 1762 3016 1765 3253
rect 1770 3213 1773 3246
rect 1786 3243 1789 3363
rect 1802 3356 1805 3433
rect 1810 3373 1813 3526
rect 1794 3353 1805 3356
rect 1794 3253 1797 3353
rect 1802 3303 1805 3336
rect 1810 3313 1813 3326
rect 1818 3216 1821 3526
rect 1826 3343 1829 3693
rect 1862 3686 1865 3793
rect 1858 3683 1865 3686
rect 1834 3606 1837 3676
rect 1858 3646 1861 3683
rect 1842 3613 1845 3646
rect 1854 3643 1861 3646
rect 1874 3643 1877 3726
rect 1834 3603 1845 3606
rect 1842 3536 1845 3603
rect 1854 3596 1857 3643
rect 1882 3636 1885 3816
rect 1890 3763 1893 3816
rect 1906 3756 1909 3833
rect 1922 3796 1925 3866
rect 1930 3803 1933 3926
rect 1938 3863 1941 3953
rect 1946 3933 1949 4016
rect 1922 3793 1933 3796
rect 1906 3753 1925 3756
rect 1906 3733 1909 3746
rect 1866 3633 1885 3636
rect 1866 3613 1869 3633
rect 1866 3596 1869 3606
rect 1874 3603 1877 3626
rect 1882 3596 1885 3616
rect 1890 3603 1893 3666
rect 1898 3613 1901 3686
rect 1922 3636 1925 3753
rect 1930 3706 1933 3793
rect 1938 3723 1941 3816
rect 1946 3723 1949 3886
rect 1930 3703 1941 3706
rect 1970 3703 1973 3946
rect 1986 3783 1989 3886
rect 1994 3883 1997 4033
rect 2002 4013 2005 4026
rect 2018 3923 2021 3966
rect 2026 3943 2029 4066
rect 2042 4013 2045 4026
rect 2042 3963 2045 4006
rect 2026 3906 2029 3936
rect 2018 3903 2029 3906
rect 2018 3846 2021 3903
rect 2034 3853 2037 3956
rect 2058 3933 2061 4196
rect 2066 4133 2069 4176
rect 2122 4156 2125 4213
rect 2146 4186 2149 4206
rect 2154 4196 2157 4216
rect 2170 4213 2177 4216
rect 2154 4193 2165 4196
rect 2142 4183 2149 4186
rect 2074 4123 2077 4156
rect 2122 4153 2133 4156
rect 2114 4133 2125 4136
rect 2130 4116 2133 4153
rect 2122 4113 2133 4116
rect 2122 4036 2125 4113
rect 2142 4086 2145 4183
rect 2162 4123 2165 4193
rect 2174 4116 2177 4213
rect 2170 4113 2177 4116
rect 2142 4083 2149 4086
rect 2122 4033 2133 4036
rect 2082 4003 2085 4016
rect 2018 3843 2029 3846
rect 2026 3826 2029 3843
rect 2010 3823 2029 3826
rect 2002 3803 2005 3816
rect 1986 3726 1989 3736
rect 1994 3733 1997 3796
rect 2002 3733 2005 3776
rect 1914 3633 1925 3636
rect 1854 3593 1861 3596
rect 1866 3593 1885 3596
rect 1858 3576 1861 3593
rect 1858 3573 1869 3576
rect 1834 3516 1837 3536
rect 1842 3533 1853 3536
rect 1842 3523 1845 3533
rect 1850 3516 1853 3526
rect 1834 3513 1853 3516
rect 1866 3506 1869 3573
rect 1914 3566 1917 3633
rect 1938 3626 1941 3703
rect 1906 3563 1917 3566
rect 1930 3623 1941 3626
rect 1906 3546 1909 3563
rect 1890 3523 1893 3546
rect 1902 3543 1909 3546
rect 1858 3503 1869 3506
rect 1734 2963 1741 2966
rect 1734 2856 1737 2963
rect 1734 2853 1741 2856
rect 1746 2853 1749 3016
rect 1754 3013 1765 3016
rect 1754 2863 1757 3013
rect 1762 2983 1765 3006
rect 1770 2993 1773 3006
rect 1778 2983 1781 3126
rect 1786 3123 1789 3146
rect 1794 3046 1797 3216
rect 1810 3203 1813 3216
rect 1818 3213 1829 3216
rect 1794 3043 1805 3046
rect 1802 3026 1805 3043
rect 1794 3023 1805 3026
rect 1794 2956 1797 3023
rect 1794 2953 1805 2956
rect 1770 2856 1773 2936
rect 1754 2853 1773 2856
rect 1706 2813 1709 2836
rect 1722 2833 1733 2836
rect 1714 2766 1717 2806
rect 1706 2763 1717 2766
rect 1706 2723 1709 2763
rect 1722 2703 1725 2816
rect 1730 2776 1733 2833
rect 1738 2803 1741 2853
rect 1730 2773 1741 2776
rect 1706 2573 1709 2606
rect 1722 2603 1725 2686
rect 1738 2586 1741 2773
rect 1754 2626 1757 2853
rect 1778 2803 1781 2866
rect 1778 2766 1781 2796
rect 1770 2763 1781 2766
rect 1770 2636 1773 2763
rect 1786 2746 1789 2856
rect 1782 2743 1789 2746
rect 1782 2656 1785 2743
rect 1782 2653 1789 2656
rect 1770 2633 1777 2636
rect 1730 2583 1741 2586
rect 1750 2623 1757 2626
rect 1694 2543 1701 2546
rect 1694 2486 1697 2543
rect 1714 2523 1717 2546
rect 1694 2483 1701 2486
rect 1654 2423 1661 2426
rect 1642 2366 1645 2386
rect 1546 2283 1549 2306
rect 1578 2273 1581 2336
rect 1590 2333 1597 2336
rect 1634 2363 1645 2366
rect 1590 2226 1593 2333
rect 1590 2223 1597 2226
rect 1578 2163 1581 2216
rect 1514 2113 1525 2116
rect 1514 2056 1517 2113
rect 1530 2066 1533 2136
rect 1554 2083 1557 2136
rect 1586 2123 1589 2206
rect 1594 2196 1597 2223
rect 1602 2213 1605 2326
rect 1594 2193 1601 2196
rect 1598 2116 1601 2193
rect 1594 2113 1601 2116
rect 1530 2063 1541 2066
rect 1514 2053 1525 2056
rect 1490 2013 1501 2016
rect 1490 1966 1493 2013
rect 1490 1963 1501 1966
rect 1458 1943 1469 1946
rect 1498 1943 1501 1963
rect 1458 1886 1461 1943
rect 1506 1936 1509 2006
rect 1458 1883 1469 1886
rect 1426 1863 1433 1866
rect 1418 1743 1421 1856
rect 1430 1766 1433 1863
rect 1442 1803 1445 1836
rect 1426 1763 1433 1766
rect 1386 1703 1389 1726
rect 1298 1503 1309 1506
rect 1306 1436 1309 1503
rect 1298 1433 1309 1436
rect 1218 1313 1225 1316
rect 1222 1246 1225 1313
rect 1218 1243 1225 1246
rect 1218 1183 1221 1243
rect 1226 1213 1229 1226
rect 1234 1193 1237 1326
rect 1242 1283 1245 1326
rect 1258 1306 1261 1326
rect 1254 1303 1261 1306
rect 1242 1216 1245 1246
rect 1254 1236 1257 1303
rect 1254 1233 1261 1236
rect 1242 1213 1253 1216
rect 1258 1213 1261 1233
rect 1258 1193 1261 1206
rect 1202 1163 1221 1166
rect 1194 1143 1205 1146
rect 1202 1056 1205 1143
rect 1194 1053 1205 1056
rect 1186 993 1189 1006
rect 1194 986 1197 1053
rect 1218 1036 1221 1163
rect 1250 1156 1253 1176
rect 1186 983 1197 986
rect 1206 1033 1221 1036
rect 1242 1153 1253 1156
rect 1242 1036 1245 1153
rect 1266 1136 1269 1356
rect 1274 1313 1277 1416
rect 1282 1413 1293 1416
rect 1298 1413 1301 1433
rect 1282 1243 1285 1413
rect 1290 1403 1301 1406
rect 1306 1353 1309 1416
rect 1290 1313 1293 1336
rect 1298 1276 1301 1346
rect 1314 1333 1317 1346
rect 1298 1273 1309 1276
rect 1274 1193 1277 1206
rect 1282 1203 1285 1216
rect 1306 1196 1309 1273
rect 1338 1213 1341 1326
rect 1298 1193 1309 1196
rect 1330 1193 1333 1206
rect 1258 1133 1269 1136
rect 1258 1056 1261 1133
rect 1258 1053 1269 1056
rect 1266 1036 1269 1053
rect 1242 1033 1253 1036
rect 1186 933 1189 983
rect 1206 946 1209 1033
rect 1218 963 1221 1016
rect 1234 946 1237 1016
rect 1242 1003 1245 1016
rect 1250 986 1253 1033
rect 1202 943 1209 946
rect 1226 943 1237 946
rect 1246 983 1253 986
rect 1258 1033 1269 1036
rect 1142 863 1149 866
rect 1170 863 1177 866
rect 1058 603 1061 616
rect 1026 533 1037 536
rect 1058 533 1061 586
rect 1074 576 1077 616
rect 1098 613 1101 806
rect 1142 776 1145 863
rect 1142 773 1149 776
rect 1114 706 1117 726
rect 1110 703 1117 706
rect 1110 616 1113 703
rect 1110 613 1117 616
rect 1122 613 1125 726
rect 1114 593 1117 613
rect 1146 583 1149 773
rect 1170 746 1173 863
rect 1170 743 1181 746
rect 1178 693 1181 743
rect 1154 613 1157 626
rect 1074 573 1085 576
rect 1026 506 1029 533
rect 1034 523 1045 526
rect 1066 523 1069 556
rect 1026 503 1037 506
rect 1034 446 1037 503
rect 1026 443 1037 446
rect 1026 403 1029 443
rect 1042 403 1045 416
rect 978 323 989 326
rect 1018 323 1021 356
rect 1058 336 1061 416
rect 1082 413 1085 573
rect 1130 523 1133 536
rect 1162 533 1165 616
rect 1170 543 1173 616
rect 1178 596 1181 606
rect 1186 603 1189 906
rect 1194 813 1197 936
rect 1194 596 1197 616
rect 1202 613 1205 943
rect 1210 903 1213 926
rect 1210 813 1213 836
rect 1226 826 1229 943
rect 1234 913 1237 936
rect 1246 926 1249 983
rect 1246 923 1253 926
rect 1258 923 1261 1033
rect 1250 906 1253 923
rect 1250 903 1261 906
rect 1226 823 1237 826
rect 1226 756 1229 816
rect 1234 783 1237 823
rect 1242 763 1245 896
rect 1258 826 1261 903
rect 1250 823 1261 826
rect 1226 753 1245 756
rect 1210 743 1229 746
rect 1210 733 1213 743
rect 1218 723 1221 736
rect 1226 723 1229 743
rect 1178 593 1197 596
rect 1202 556 1205 606
rect 1186 553 1205 556
rect 1178 513 1181 546
rect 1186 523 1189 553
rect 1202 543 1205 553
rect 1210 543 1213 566
rect 1218 526 1221 616
rect 1210 523 1221 526
rect 1210 466 1213 523
rect 1058 333 1069 336
rect 938 133 941 146
rect 962 133 965 146
rect 978 143 981 323
rect 850 113 853 126
rect 858 103 861 126
rect 890 113 893 126
rect 994 123 997 216
rect 1002 203 1005 216
rect 1010 196 1013 206
rect 1018 203 1021 216
rect 1026 196 1029 216
rect 1042 213 1045 256
rect 1010 193 1029 196
rect 1034 193 1037 206
rect 1042 123 1045 206
rect 1066 166 1069 333
rect 1082 303 1085 326
rect 1090 213 1093 326
rect 1106 323 1109 416
rect 1154 393 1157 416
rect 1162 413 1165 466
rect 1210 463 1221 466
rect 1122 323 1125 336
rect 1162 266 1165 406
rect 1178 333 1181 416
rect 1186 393 1189 406
rect 1194 346 1197 416
rect 1218 413 1221 463
rect 1202 383 1205 406
rect 1194 343 1201 346
rect 1162 263 1173 266
rect 1154 193 1157 216
rect 1162 213 1165 246
rect 1170 206 1173 263
rect 1178 213 1181 326
rect 1162 203 1173 206
rect 1058 163 1069 166
rect 1058 133 1061 163
rect 1162 156 1165 203
rect 1186 193 1189 336
rect 1198 236 1201 343
rect 1218 333 1221 406
rect 1226 403 1229 646
rect 1234 633 1237 736
rect 1242 733 1245 753
rect 1234 533 1237 616
rect 1242 613 1245 726
rect 1250 533 1253 823
rect 1258 793 1261 806
rect 1266 793 1269 806
rect 1274 803 1277 1186
rect 1298 1176 1301 1193
rect 1290 1173 1301 1176
rect 1290 1126 1293 1173
rect 1346 1146 1349 1216
rect 1354 1173 1357 1576
rect 1370 1573 1381 1576
rect 1370 1496 1373 1573
rect 1370 1493 1381 1496
rect 1378 1473 1381 1493
rect 1386 1466 1389 1686
rect 1402 1636 1405 1726
rect 1410 1723 1417 1726
rect 1414 1636 1417 1723
rect 1370 1463 1389 1466
rect 1394 1633 1405 1636
rect 1410 1633 1417 1636
rect 1370 1376 1373 1463
rect 1394 1416 1397 1633
rect 1402 1533 1405 1546
rect 1410 1533 1413 1633
rect 1418 1593 1421 1616
rect 1418 1533 1421 1556
rect 1402 1516 1405 1526
rect 1410 1523 1421 1526
rect 1402 1513 1413 1516
rect 1386 1413 1397 1416
rect 1402 1413 1405 1426
rect 1370 1373 1381 1376
rect 1378 1286 1381 1373
rect 1370 1283 1381 1286
rect 1362 1196 1365 1216
rect 1370 1203 1373 1283
rect 1378 1196 1381 1206
rect 1386 1203 1389 1413
rect 1394 1393 1397 1406
rect 1410 1396 1413 1513
rect 1406 1393 1413 1396
rect 1394 1313 1397 1326
rect 1362 1193 1381 1196
rect 1306 1133 1309 1146
rect 1338 1143 1349 1146
rect 1290 1123 1301 1126
rect 1282 933 1285 956
rect 1298 943 1301 1123
rect 1298 873 1301 936
rect 1322 923 1325 1126
rect 1338 1123 1341 1143
rect 1346 1003 1349 1136
rect 1354 1123 1357 1146
rect 1362 1043 1365 1136
rect 1378 1116 1381 1126
rect 1386 1123 1389 1196
rect 1394 1116 1397 1216
rect 1406 1206 1409 1393
rect 1418 1213 1421 1416
rect 1426 1386 1429 1763
rect 1434 1673 1437 1746
rect 1450 1733 1453 1816
rect 1458 1763 1461 1866
rect 1466 1736 1469 1883
rect 1474 1863 1477 1926
rect 1482 1833 1485 1936
rect 1490 1816 1493 1936
rect 1486 1813 1493 1816
rect 1498 1933 1509 1936
rect 1486 1746 1489 1813
rect 1498 1766 1501 1933
rect 1506 1813 1509 1926
rect 1522 1893 1525 2053
rect 1538 1916 1541 2063
rect 1562 2006 1565 2016
rect 1570 2013 1573 2026
rect 1562 2003 1589 2006
rect 1586 1993 1589 2003
rect 1594 1963 1597 2113
rect 1602 1973 1605 2026
rect 1634 2016 1637 2363
rect 1654 2356 1657 2423
rect 1654 2353 1661 2356
rect 1650 2313 1653 2336
rect 1658 2296 1661 2353
rect 1666 2333 1669 2416
rect 1674 2323 1677 2356
rect 1682 2296 1685 2376
rect 1650 2293 1661 2296
rect 1666 2293 1685 2296
rect 1650 2226 1653 2293
rect 1650 2223 1661 2226
rect 1650 2186 1653 2206
rect 1646 2183 1653 2186
rect 1646 2096 1649 2183
rect 1658 2106 1661 2223
rect 1666 2176 1669 2293
rect 1674 2213 1677 2226
rect 1690 2213 1693 2246
rect 1698 2236 1701 2483
rect 1722 2476 1725 2566
rect 1714 2473 1725 2476
rect 1714 2286 1717 2473
rect 1730 2426 1733 2583
rect 1750 2566 1753 2623
rect 1738 2563 1753 2566
rect 1762 2563 1765 2616
rect 1774 2566 1777 2633
rect 1774 2563 1781 2566
rect 1738 2496 1741 2563
rect 1738 2493 1749 2496
rect 1726 2423 1733 2426
rect 1746 2426 1749 2493
rect 1746 2423 1753 2426
rect 1726 2306 1729 2423
rect 1738 2353 1741 2416
rect 1750 2376 1753 2423
rect 1762 2383 1765 2536
rect 1778 2483 1781 2563
rect 1778 2416 1781 2436
rect 1774 2413 1781 2416
rect 1746 2373 1753 2376
rect 1726 2303 1733 2306
rect 1714 2283 1725 2286
rect 1722 2263 1725 2283
rect 1698 2233 1717 2236
rect 1682 2193 1685 2206
rect 1706 2196 1709 2226
rect 1698 2193 1709 2196
rect 1666 2173 1685 2176
rect 1674 2123 1677 2166
rect 1682 2123 1685 2173
rect 1658 2103 1669 2106
rect 1646 2093 1653 2096
rect 1634 2013 1645 2016
rect 1530 1913 1541 1916
rect 1530 1766 1533 1913
rect 1546 1786 1549 1896
rect 1554 1856 1557 1876
rect 1554 1853 1561 1856
rect 1498 1763 1509 1766
rect 1458 1733 1469 1736
rect 1474 1733 1477 1746
rect 1486 1743 1493 1746
rect 1458 1656 1461 1733
rect 1466 1723 1477 1726
rect 1458 1653 1469 1656
rect 1434 1613 1445 1616
rect 1434 1523 1437 1536
rect 1434 1403 1437 1446
rect 1442 1413 1445 1596
rect 1450 1566 1453 1646
rect 1450 1563 1457 1566
rect 1454 1466 1457 1563
rect 1466 1506 1469 1653
rect 1474 1613 1477 1626
rect 1482 1593 1485 1726
rect 1490 1723 1493 1743
rect 1506 1666 1509 1763
rect 1522 1763 1533 1766
rect 1538 1783 1549 1786
rect 1522 1676 1525 1763
rect 1538 1686 1541 1783
rect 1558 1756 1561 1853
rect 1554 1753 1561 1756
rect 1554 1733 1557 1753
rect 1546 1703 1549 1726
rect 1578 1723 1581 1936
rect 1618 1923 1621 1996
rect 1642 1933 1645 2013
rect 1650 1973 1653 2093
rect 1666 2036 1669 2103
rect 1698 2096 1701 2193
rect 1698 2093 1709 2096
rect 1662 2033 1669 2036
rect 1662 1966 1665 2033
rect 1674 2006 1677 2016
rect 1682 2013 1685 2056
rect 1698 2006 1701 2076
rect 1706 2013 1709 2093
rect 1674 2003 1701 2006
rect 1714 1986 1717 2233
rect 1730 2153 1733 2303
rect 1746 2286 1749 2373
rect 1774 2296 1777 2413
rect 1786 2373 1789 2653
rect 1786 2303 1789 2326
rect 1774 2293 1781 2296
rect 1746 2283 1765 2286
rect 1746 2246 1749 2266
rect 1746 2243 1753 2246
rect 1658 1963 1665 1966
rect 1706 1983 1717 1986
rect 1658 1823 1661 1963
rect 1674 1923 1677 1936
rect 1682 1856 1685 1936
rect 1706 1876 1709 1983
rect 1722 1953 1725 2146
rect 1722 1923 1725 1946
rect 1730 1923 1733 2056
rect 1738 2003 1741 2216
rect 1750 2166 1753 2243
rect 1746 2163 1753 2166
rect 1746 2076 1749 2163
rect 1762 2133 1765 2283
rect 1778 2223 1781 2293
rect 1794 2236 1797 2916
rect 1802 2883 1805 2953
rect 1810 2923 1813 3016
rect 1818 2853 1821 3186
rect 1826 3093 1829 3213
rect 1834 3116 1837 3336
rect 1842 3323 1845 3416
rect 1858 3366 1861 3503
rect 1902 3486 1905 3543
rect 1922 3503 1925 3536
rect 1930 3493 1933 3623
rect 1938 3503 1941 3526
rect 1902 3483 1909 3486
rect 1858 3363 1869 3366
rect 1866 3316 1869 3363
rect 1858 3313 1869 3316
rect 1842 3123 1845 3216
rect 1858 3213 1861 3313
rect 1834 3113 1841 3116
rect 1838 3036 1841 3113
rect 1850 3046 1853 3096
rect 1850 3043 1857 3046
rect 1838 3033 1845 3036
rect 1826 2983 1829 3006
rect 1834 2993 1837 3016
rect 1842 3003 1845 3033
rect 1854 2996 1857 3043
rect 1866 3013 1869 3256
rect 1890 3253 1893 3406
rect 1874 3153 1877 3206
rect 1882 3203 1885 3246
rect 1850 2993 1857 2996
rect 1802 2813 1805 2826
rect 1802 2683 1805 2806
rect 1818 2723 1821 2836
rect 1826 2716 1829 2886
rect 1834 2813 1837 2926
rect 1850 2906 1853 2993
rect 1858 2923 1861 2936
rect 1866 2923 1869 3006
rect 1874 2923 1877 3016
rect 1882 2996 1885 3016
rect 1890 3013 1893 3216
rect 1898 3203 1901 3216
rect 1906 3016 1909 3483
rect 1946 3453 1949 3606
rect 1954 3583 1957 3606
rect 1962 3563 1965 3616
rect 1978 3613 1981 3726
rect 1986 3723 2005 3726
rect 1986 3613 1989 3636
rect 1970 3543 1973 3606
rect 1986 3583 1989 3606
rect 1970 3523 1973 3536
rect 1986 3533 1989 3566
rect 1986 3503 1989 3526
rect 1994 3523 1997 3706
rect 2010 3603 2013 3823
rect 2018 3763 2021 3806
rect 2026 3803 2029 3816
rect 2034 3793 2037 3806
rect 2050 3803 2061 3806
rect 2018 3703 2021 3756
rect 2026 3733 2029 3776
rect 2058 3773 2061 3803
rect 2026 3653 2029 3726
rect 2034 3723 2037 3756
rect 2066 3753 2069 3806
rect 2050 3733 2053 3746
rect 2066 3646 2069 3676
rect 2074 3653 2077 3776
rect 2082 3673 2085 3996
rect 2090 3913 2093 3936
rect 2106 3923 2109 4016
rect 2130 4013 2133 4033
rect 2146 4023 2149 4083
rect 2114 3933 2117 3946
rect 2122 3923 2125 4006
rect 2146 3933 2149 3966
rect 2162 3933 2165 4016
rect 2154 3913 2157 3926
rect 2106 3776 2109 3886
rect 2090 3773 2109 3776
rect 2026 3543 2029 3616
rect 2042 3533 2045 3616
rect 2058 3613 2061 3646
rect 2066 3643 2077 3646
rect 2090 3606 2093 3773
rect 2122 3766 2125 3786
rect 2130 3776 2133 3816
rect 2170 3783 2173 4113
rect 2186 4016 2189 4426
rect 2206 4423 2213 4426
rect 2234 4443 2245 4446
rect 2206 4346 2209 4423
rect 2206 4343 2213 4346
rect 2218 4343 2221 4416
rect 2226 4393 2229 4406
rect 2210 4323 2213 4343
rect 2218 4323 2221 4336
rect 2226 4263 2229 4336
rect 2234 4256 2237 4443
rect 2250 4436 2253 4566
rect 2266 4536 2269 4616
rect 2242 4433 2253 4436
rect 2258 4433 2261 4536
rect 2266 4533 2277 4536
rect 2242 4403 2245 4433
rect 2250 4413 2253 4426
rect 2266 4423 2269 4526
rect 2274 4416 2277 4533
rect 2266 4413 2277 4416
rect 2266 4403 2269 4413
rect 2274 4383 2277 4406
rect 2258 4333 2261 4366
rect 2282 4333 2285 4536
rect 2290 4506 2293 4596
rect 2298 4533 2301 4616
rect 2306 4543 2325 4546
rect 2306 4523 2309 4543
rect 2290 4503 2301 4506
rect 2298 4436 2301 4503
rect 2314 4453 2317 4536
rect 2322 4533 2325 4543
rect 2322 4473 2325 4526
rect 2338 4523 2341 4616
rect 2378 4593 2381 4606
rect 2354 4533 2357 4556
rect 2378 4533 2381 4556
rect 2346 4513 2349 4526
rect 2386 4493 2389 4526
rect 2402 4523 2405 4536
rect 2410 4533 2413 4616
rect 2418 4543 2437 4546
rect 2418 4523 2421 4543
rect 2426 4453 2429 4536
rect 2434 4533 2437 4543
rect 2434 4463 2437 4526
rect 2466 4523 2469 4616
rect 2474 4523 2477 4686
rect 2538 4613 2541 4626
rect 2578 4613 2581 4626
rect 2498 4463 2501 4606
rect 2298 4433 2309 4436
rect 2290 4413 2293 4426
rect 2306 4343 2309 4433
rect 2330 4413 2333 4426
rect 2242 4323 2253 4326
rect 2266 4283 2269 4326
rect 2234 4253 2269 4256
rect 2210 4213 2213 4226
rect 2250 4213 2253 4226
rect 2266 4206 2269 4253
rect 2298 4233 2301 4326
rect 2322 4323 2325 4386
rect 2386 4346 2389 4416
rect 2418 4413 2421 4426
rect 2394 4356 2397 4406
rect 2394 4353 2405 4356
rect 2378 4343 2389 4346
rect 2330 4293 2333 4326
rect 2226 4166 2229 4206
rect 2210 4163 2229 4166
rect 2258 4203 2269 4206
rect 2210 4063 2213 4163
rect 2186 4013 2197 4016
rect 2178 3993 2181 4006
rect 2178 3893 2181 3986
rect 2194 3906 2197 4013
rect 2210 4006 2213 4016
rect 2218 4013 2221 4036
rect 2242 4013 2245 4046
rect 2210 4003 2237 4006
rect 2210 3923 2213 4003
rect 2226 3933 2229 3946
rect 2234 3933 2237 3956
rect 2250 3916 2253 4006
rect 2186 3903 2197 3906
rect 2242 3913 2253 3916
rect 2186 3883 2189 3903
rect 2202 3826 2205 3876
rect 2242 3826 2245 3913
rect 2258 3873 2261 4203
rect 2266 4013 2269 4026
rect 2274 3933 2277 3966
rect 2202 3823 2213 3826
rect 2242 3823 2253 3826
rect 2130 3773 2141 3776
rect 2118 3763 2125 3766
rect 2098 3683 2101 3726
rect 2118 3696 2121 3763
rect 2130 3706 2133 3726
rect 2138 3723 2141 3773
rect 2146 3753 2173 3756
rect 2146 3733 2149 3753
rect 2154 3733 2157 3746
rect 2130 3703 2149 3706
rect 2118 3693 2125 3696
rect 2106 3613 2109 3656
rect 2058 3503 2061 3526
rect 2066 3523 2069 3606
rect 2090 3603 2109 3606
rect 2114 3603 2117 3636
rect 2122 3613 2125 3693
rect 2138 3613 2141 3686
rect 2146 3603 2149 3703
rect 2162 3616 2165 3736
rect 2170 3723 2173 3753
rect 2178 3733 2181 3816
rect 2186 3733 2189 3816
rect 2170 3696 2173 3716
rect 2170 3693 2177 3696
rect 2174 3636 2177 3693
rect 2154 3613 2165 3616
rect 2170 3633 2177 3636
rect 2098 3503 2101 3526
rect 1922 3393 1925 3406
rect 1938 3336 1941 3356
rect 1934 3333 1941 3336
rect 1914 3183 1917 3216
rect 1922 3213 1925 3326
rect 1934 3236 1937 3333
rect 1946 3246 1949 3416
rect 1954 3296 1957 3496
rect 1962 3353 1965 3456
rect 1970 3413 1973 3426
rect 1970 3333 1973 3396
rect 2002 3336 2005 3416
rect 2010 3413 2013 3426
rect 2050 3393 2053 3406
rect 2066 3363 2069 3406
rect 2098 3366 2101 3396
rect 2090 3363 2101 3366
rect 2002 3333 2013 3336
rect 1954 3293 1965 3296
rect 1946 3243 1953 3246
rect 1934 3233 1941 3236
rect 1938 3216 1941 3233
rect 1930 3213 1941 3216
rect 1930 3166 1933 3206
rect 1914 3163 1933 3166
rect 1914 3133 1917 3163
rect 1922 3123 1925 3156
rect 1930 3056 1933 3146
rect 1938 3123 1941 3206
rect 1950 3116 1953 3243
rect 1946 3113 1953 3116
rect 1930 3053 1941 3056
rect 1898 3013 1909 3016
rect 1914 3013 1933 3016
rect 1882 2993 1889 2996
rect 1886 2916 1889 2993
rect 1898 2953 1901 3013
rect 1906 2933 1909 3006
rect 1914 2973 1917 3013
rect 1922 3003 1933 3006
rect 1938 3003 1941 3053
rect 1922 2933 1925 2986
rect 1930 2933 1933 2956
rect 1946 2936 1949 3113
rect 1962 3046 1965 3293
rect 2002 3286 2005 3326
rect 1994 3283 2005 3286
rect 1978 3203 1981 3216
rect 1994 3146 1997 3283
rect 2010 3276 2013 3333
rect 2050 3306 2053 3326
rect 2042 3303 2053 3306
rect 2010 3273 2021 3276
rect 2018 3226 2021 3273
rect 2042 3236 2045 3303
rect 2042 3233 2053 3236
rect 2010 3223 2021 3226
rect 2010 3203 2013 3223
rect 1994 3143 2005 3146
rect 1978 3113 1981 3136
rect 2002 3123 2005 3143
rect 2010 3133 2013 3186
rect 1954 3043 1965 3046
rect 2010 3043 2013 3126
rect 2018 3096 2021 3136
rect 2026 3113 2029 3126
rect 2018 3093 2025 3096
rect 1954 2993 1957 3043
rect 1970 3013 1973 3026
rect 1942 2933 1949 2936
rect 1882 2913 1889 2916
rect 1850 2903 1861 2906
rect 1858 2826 1861 2903
rect 1882 2866 1885 2913
rect 1842 2813 1845 2826
rect 1850 2823 1861 2826
rect 1874 2863 1885 2866
rect 1850 2806 1853 2823
rect 1810 2713 1829 2716
rect 1834 2803 1853 2806
rect 1802 2423 1805 2606
rect 1810 2433 1813 2713
rect 1834 2666 1837 2803
rect 1850 2733 1853 2746
rect 1874 2743 1877 2863
rect 1834 2663 1841 2666
rect 1826 2563 1829 2656
rect 1838 2546 1841 2663
rect 1834 2543 1841 2546
rect 1834 2523 1837 2543
rect 1818 2403 1821 2476
rect 1810 2316 1813 2386
rect 1826 2363 1829 2436
rect 1818 2323 1829 2326
rect 1810 2313 1829 2316
rect 1790 2233 1797 2236
rect 1778 2193 1781 2216
rect 1746 2073 1757 2076
rect 1754 1956 1757 2073
rect 1790 2036 1793 2233
rect 1790 2033 1797 2036
rect 1786 2003 1789 2016
rect 1794 1986 1797 2033
rect 1802 2013 1805 2226
rect 1826 2203 1829 2313
rect 1834 2303 1837 2326
rect 1810 2123 1813 2196
rect 1842 2193 1845 2216
rect 1850 2176 1853 2706
rect 1890 2703 1893 2856
rect 1914 2836 1917 2926
rect 1898 2833 1917 2836
rect 1898 2803 1901 2833
rect 1942 2806 1945 2933
rect 1954 2813 1957 2926
rect 1978 2923 1981 2936
rect 1986 2816 1989 3006
rect 2002 2943 2005 3006
rect 2010 2993 2013 3016
rect 2022 2996 2025 3093
rect 2034 3003 2037 3136
rect 2018 2993 2025 2996
rect 2018 2973 2021 2993
rect 2010 2943 2029 2946
rect 2010 2933 2013 2943
rect 2018 2923 2021 2936
rect 2026 2923 2029 2943
rect 2034 2933 2037 2986
rect 2042 2936 2045 3216
rect 2050 3133 2053 3233
rect 2058 3213 2061 3326
rect 2090 3296 2093 3363
rect 2106 3306 2109 3603
rect 2146 3543 2149 3586
rect 2154 3563 2157 3613
rect 2146 3523 2149 3536
rect 2162 3533 2165 3606
rect 2170 3516 2173 3633
rect 2186 3616 2189 3726
rect 2194 3713 2197 3786
rect 2210 3696 2213 3823
rect 2250 3803 2253 3823
rect 2234 3713 2237 3736
rect 2250 3733 2253 3746
rect 2178 3613 2189 3616
rect 2202 3693 2213 3696
rect 2178 3523 2181 3613
rect 2186 3576 2189 3606
rect 2202 3586 2205 3693
rect 2218 3603 2221 3676
rect 2242 3613 2245 3726
rect 2202 3583 2221 3586
rect 2186 3573 2197 3576
rect 2194 3523 2197 3573
rect 2202 3533 2205 3566
rect 2210 3533 2213 3546
rect 2170 3513 2181 3516
rect 2114 3413 2117 3426
rect 2106 3303 2113 3306
rect 2090 3293 2101 3296
rect 2058 3186 2061 3206
rect 2058 3183 2065 3186
rect 2062 3126 2065 3183
rect 2058 3123 2065 3126
rect 2074 3123 2077 3276
rect 2098 3213 2101 3293
rect 2110 3236 2113 3303
rect 2106 3233 2113 3236
rect 2106 3213 2109 3233
rect 2122 3226 2125 3356
rect 2122 3223 2129 3226
rect 2050 2996 2053 3046
rect 2058 3003 2061 3123
rect 2090 3043 2093 3206
rect 2106 3183 2109 3206
rect 2106 3076 2109 3136
rect 2114 3113 2117 3216
rect 2126 3166 2129 3223
rect 2122 3163 2129 3166
rect 2122 3116 2125 3163
rect 2130 3133 2133 3146
rect 2138 3126 2141 3216
rect 2146 3133 2149 3416
rect 2154 3413 2157 3426
rect 2154 3313 2157 3326
rect 2162 3186 2165 3376
rect 2170 3323 2173 3406
rect 2178 3393 2181 3513
rect 2178 3203 2181 3336
rect 2162 3183 2173 3186
rect 2154 3133 2157 3176
rect 2170 3126 2173 3183
rect 2130 3123 2141 3126
rect 2162 3123 2173 3126
rect 2122 3113 2129 3116
rect 2098 3073 2109 3076
rect 2050 2993 2061 2996
rect 2066 2993 2069 3016
rect 2082 3013 2085 3026
rect 2098 3016 2101 3073
rect 2126 3066 2129 3113
rect 2126 3063 2133 3066
rect 2098 3013 2117 3016
rect 2042 2933 2053 2936
rect 1986 2813 1997 2816
rect 1914 2783 1917 2806
rect 1942 2803 1949 2806
rect 1898 2723 1901 2736
rect 1930 2723 1933 2746
rect 1938 2723 1941 2736
rect 1946 2643 1949 2803
rect 2010 2783 2013 2806
rect 1890 2613 1893 2626
rect 1866 2603 1885 2606
rect 1874 2533 1877 2546
rect 1866 2386 1869 2526
rect 1882 2523 1885 2603
rect 1898 2586 1901 2616
rect 1930 2613 1933 2626
rect 1978 2603 1981 2726
rect 1890 2583 1901 2586
rect 1890 2466 1893 2583
rect 1906 2546 1909 2566
rect 1898 2533 1901 2546
rect 1906 2543 1917 2546
rect 1882 2463 1893 2466
rect 1882 2403 1885 2463
rect 1914 2436 1917 2543
rect 1978 2533 1981 2546
rect 1962 2513 1965 2526
rect 1906 2433 1917 2436
rect 1970 2433 1973 2526
rect 1986 2523 1989 2586
rect 1890 2413 1893 2426
rect 1906 2413 1909 2433
rect 1866 2383 1877 2386
rect 1866 2336 1869 2376
rect 1874 2353 1877 2383
rect 1898 2373 1901 2406
rect 1866 2333 1877 2336
rect 1842 2173 1853 2176
rect 1842 2046 1845 2173
rect 1874 2166 1877 2333
rect 1866 2163 1877 2166
rect 1866 2106 1869 2163
rect 1898 2123 1901 2136
rect 1906 2106 1909 2356
rect 1914 2323 1917 2366
rect 1930 2363 1933 2406
rect 1930 2343 1949 2346
rect 1930 2333 1933 2343
rect 1930 2213 1933 2326
rect 1938 2323 1941 2336
rect 1946 2323 1949 2343
rect 1954 2306 1957 2336
rect 1962 2333 1965 2396
rect 1954 2303 1965 2306
rect 1938 2213 1957 2216
rect 1938 2203 1941 2213
rect 1946 2136 1949 2206
rect 1962 2203 1965 2303
rect 1866 2103 1877 2106
rect 1842 2043 1853 2046
rect 1746 1953 1757 1956
rect 1778 1983 1797 1986
rect 1746 1933 1749 1953
rect 1706 1873 1717 1876
rect 1674 1853 1685 1856
rect 1714 1853 1717 1873
rect 1586 1713 1589 1736
rect 1602 1723 1605 1816
rect 1650 1766 1653 1806
rect 1642 1763 1653 1766
rect 1538 1683 1549 1686
rect 1522 1673 1533 1676
rect 1498 1663 1509 1666
rect 1498 1646 1501 1663
rect 1490 1643 1501 1646
rect 1490 1596 1493 1643
rect 1490 1593 1501 1596
rect 1514 1593 1517 1606
rect 1530 1593 1533 1673
rect 1498 1566 1501 1593
rect 1546 1586 1549 1683
rect 1618 1646 1621 1726
rect 1642 1656 1645 1763
rect 1674 1756 1677 1853
rect 1714 1813 1717 1826
rect 1666 1753 1677 1756
rect 1642 1653 1653 1656
rect 1610 1643 1621 1646
rect 1578 1603 1581 1626
rect 1610 1596 1613 1643
rect 1634 1613 1637 1636
rect 1538 1583 1549 1586
rect 1498 1563 1505 1566
rect 1482 1523 1485 1536
rect 1490 1523 1493 1546
rect 1502 1516 1505 1563
rect 1538 1553 1541 1583
rect 1522 1523 1525 1536
rect 1570 1523 1573 1596
rect 1610 1593 1621 1596
rect 1618 1533 1621 1593
rect 1634 1563 1637 1606
rect 1642 1583 1645 1616
rect 1650 1603 1653 1653
rect 1498 1513 1505 1516
rect 1466 1503 1477 1506
rect 1450 1463 1457 1466
rect 1450 1443 1453 1463
rect 1458 1403 1461 1426
rect 1426 1383 1433 1386
rect 1430 1306 1433 1383
rect 1442 1323 1445 1336
rect 1450 1333 1453 1386
rect 1474 1376 1477 1503
rect 1498 1406 1501 1513
rect 1506 1413 1509 1426
rect 1498 1403 1509 1406
rect 1466 1373 1477 1376
rect 1466 1353 1469 1373
rect 1498 1326 1501 1346
rect 1466 1313 1469 1326
rect 1490 1323 1501 1326
rect 1430 1303 1437 1306
rect 1434 1236 1437 1303
rect 1426 1233 1437 1236
rect 1406 1203 1413 1206
rect 1410 1166 1413 1203
rect 1378 1113 1397 1116
rect 1406 1163 1413 1166
rect 1378 1096 1381 1113
rect 1378 1093 1389 1096
rect 1386 1036 1389 1093
rect 1406 1086 1409 1163
rect 1406 1083 1413 1086
rect 1378 1033 1389 1036
rect 1378 1016 1381 1033
rect 1410 1026 1413 1083
rect 1370 1013 1381 1016
rect 1402 1023 1413 1026
rect 1314 813 1317 866
rect 1282 793 1285 806
rect 1258 723 1261 766
rect 1274 756 1277 776
rect 1270 753 1277 756
rect 1270 696 1273 753
rect 1282 706 1285 786
rect 1306 726 1309 806
rect 1330 773 1333 896
rect 1338 803 1341 906
rect 1346 813 1349 926
rect 1362 753 1365 946
rect 1370 903 1373 1013
rect 1378 923 1381 1006
rect 1386 983 1389 1006
rect 1402 956 1405 1023
rect 1402 953 1413 956
rect 1386 886 1389 936
rect 1378 883 1389 886
rect 1378 786 1381 883
rect 1394 813 1397 936
rect 1402 913 1405 926
rect 1410 896 1413 953
rect 1418 943 1421 1016
rect 1418 903 1421 926
rect 1426 896 1429 1233
rect 1434 1106 1437 1206
rect 1442 1123 1445 1216
rect 1450 1183 1453 1216
rect 1458 1193 1461 1286
rect 1466 1196 1469 1216
rect 1474 1203 1477 1316
rect 1490 1236 1493 1323
rect 1506 1246 1509 1403
rect 1514 1393 1517 1416
rect 1546 1413 1549 1426
rect 1538 1336 1541 1356
rect 1538 1333 1545 1336
rect 1506 1243 1517 1246
rect 1490 1233 1501 1236
rect 1482 1196 1485 1206
rect 1490 1203 1493 1216
rect 1466 1193 1485 1196
rect 1434 1103 1445 1106
rect 1442 1036 1445 1103
rect 1434 1033 1445 1036
rect 1434 1013 1437 1033
rect 1434 953 1437 1006
rect 1434 913 1437 936
rect 1442 933 1445 1016
rect 1450 933 1453 946
rect 1406 893 1413 896
rect 1418 893 1429 896
rect 1406 806 1409 893
rect 1418 876 1421 893
rect 1426 883 1437 886
rect 1418 873 1429 876
rect 1406 803 1413 806
rect 1378 783 1405 786
rect 1378 733 1381 756
rect 1290 713 1293 726
rect 1298 723 1309 726
rect 1330 713 1333 726
rect 1282 703 1293 706
rect 1270 693 1277 696
rect 1274 656 1277 693
rect 1274 653 1281 656
rect 1258 603 1261 626
rect 1266 613 1269 646
rect 1278 606 1281 653
rect 1274 603 1281 606
rect 1258 533 1261 546
rect 1242 513 1245 526
rect 1234 413 1237 496
rect 1266 473 1269 526
rect 1250 413 1253 426
rect 1258 403 1261 436
rect 1266 413 1269 446
rect 1266 393 1269 406
rect 1194 233 1201 236
rect 1194 216 1197 233
rect 1194 213 1205 216
rect 1210 213 1213 326
rect 1194 186 1197 206
rect 1154 153 1165 156
rect 1186 183 1197 186
rect 1106 113 1109 126
rect 1138 123 1141 146
rect 1146 113 1149 126
rect 1154 123 1157 153
rect 1162 143 1181 146
rect 1162 133 1165 143
rect 1162 93 1165 126
rect 1170 123 1173 136
rect 1178 123 1181 143
rect 1186 133 1189 183
rect 1202 113 1205 213
rect 1218 203 1221 226
rect 1226 213 1229 326
rect 1218 123 1221 136
rect 1234 123 1237 256
rect 1242 213 1245 346
rect 1266 316 1269 336
rect 1258 313 1269 316
rect 1258 236 1261 313
rect 1274 243 1277 603
rect 1290 566 1293 703
rect 1394 696 1397 726
rect 1390 693 1397 696
rect 1298 603 1301 656
rect 1282 563 1293 566
rect 1282 413 1285 563
rect 1290 533 1293 556
rect 1290 403 1293 516
rect 1306 513 1309 616
rect 1346 603 1349 616
rect 1354 613 1357 626
rect 1322 533 1325 546
rect 1330 433 1333 536
rect 1338 503 1341 536
rect 1346 533 1349 596
rect 1362 533 1365 606
rect 1370 593 1373 616
rect 1354 513 1357 526
rect 1378 493 1381 646
rect 1390 636 1393 693
rect 1390 633 1397 636
rect 1386 533 1389 616
rect 1394 603 1397 633
rect 1298 346 1301 416
rect 1306 403 1309 416
rect 1314 403 1317 426
rect 1338 413 1341 426
rect 1290 343 1301 346
rect 1258 233 1269 236
rect 1282 233 1285 336
rect 1290 263 1293 343
rect 1322 323 1325 336
rect 1330 313 1333 336
rect 1346 333 1349 346
rect 1338 296 1341 326
rect 1330 293 1341 296
rect 1346 293 1349 326
rect 1330 236 1333 293
rect 1354 246 1357 456
rect 1378 413 1381 426
rect 1362 313 1365 326
rect 1370 253 1373 336
rect 1378 313 1381 326
rect 1346 243 1357 246
rect 1330 233 1341 236
rect 1266 156 1269 233
rect 1338 213 1341 233
rect 1282 193 1285 206
rect 1346 173 1349 243
rect 1370 183 1373 206
rect 1386 203 1389 326
rect 1394 193 1397 326
rect 1402 213 1405 783
rect 1410 766 1413 803
rect 1410 763 1417 766
rect 1414 666 1417 763
rect 1410 663 1417 666
rect 1410 643 1413 663
rect 1410 523 1413 566
rect 1418 533 1421 636
rect 1426 326 1429 873
rect 1434 833 1437 883
rect 1442 813 1445 926
rect 1450 796 1453 906
rect 1450 793 1461 796
rect 1458 766 1461 793
rect 1458 763 1465 766
rect 1434 596 1437 616
rect 1442 603 1445 696
rect 1462 686 1465 763
rect 1474 736 1477 1156
rect 1498 1153 1501 1233
rect 1514 1176 1517 1243
rect 1530 1213 1533 1326
rect 1542 1226 1545 1333
rect 1538 1223 1545 1226
rect 1538 1196 1541 1223
rect 1554 1213 1557 1336
rect 1506 1173 1517 1176
rect 1534 1193 1541 1196
rect 1506 1056 1509 1173
rect 1534 1126 1537 1193
rect 1546 1133 1549 1206
rect 1562 1203 1565 1296
rect 1534 1123 1541 1126
rect 1538 1103 1541 1123
rect 1554 1066 1557 1126
rect 1554 1063 1573 1066
rect 1506 1053 1513 1056
rect 1510 996 1513 1053
rect 1506 993 1513 996
rect 1506 976 1509 993
rect 1498 973 1509 976
rect 1498 793 1501 973
rect 1522 923 1525 1016
rect 1554 946 1557 1056
rect 1570 1013 1573 1063
rect 1578 1053 1581 1396
rect 1594 1343 1597 1526
rect 1650 1486 1653 1526
rect 1594 1213 1597 1336
rect 1626 1256 1629 1486
rect 1642 1483 1653 1486
rect 1642 1436 1645 1483
rect 1642 1433 1653 1436
rect 1650 1413 1653 1433
rect 1634 1313 1637 1326
rect 1650 1323 1653 1336
rect 1658 1333 1661 1616
rect 1666 1393 1669 1753
rect 1674 1613 1677 1666
rect 1682 1593 1685 1606
rect 1674 1413 1677 1476
rect 1666 1333 1669 1376
rect 1674 1323 1677 1336
rect 1682 1306 1685 1576
rect 1690 1556 1693 1646
rect 1698 1636 1701 1726
rect 1706 1716 1709 1806
rect 1722 1803 1725 1916
rect 1730 1753 1733 1846
rect 1778 1826 1781 1983
rect 1802 1913 1805 1936
rect 1810 1933 1813 1946
rect 1826 1893 1829 2016
rect 1834 2013 1837 2026
rect 1850 1936 1853 2043
rect 1858 2033 1861 2096
rect 1874 2046 1877 2103
rect 1866 2043 1877 2046
rect 1890 2103 1909 2106
rect 1866 2023 1869 2043
rect 1890 1986 1893 2103
rect 1914 2086 1917 2136
rect 1906 2083 1917 2086
rect 1906 2006 1909 2083
rect 1922 2033 1925 2126
rect 1930 2103 1933 2136
rect 1938 2133 1949 2136
rect 1938 2123 1949 2126
rect 1938 2106 1941 2123
rect 1938 2103 1949 2106
rect 1946 2036 1949 2103
rect 1938 2033 1949 2036
rect 1906 2003 1917 2006
rect 1890 1983 1909 1986
rect 1850 1933 1861 1936
rect 1898 1933 1901 1966
rect 1842 1896 1845 1926
rect 1838 1893 1845 1896
rect 1738 1813 1741 1826
rect 1778 1823 1813 1826
rect 1754 1776 1757 1816
rect 1778 1793 1781 1806
rect 1786 1803 1797 1806
rect 1802 1793 1805 1816
rect 1754 1773 1765 1776
rect 1714 1743 1733 1746
rect 1714 1733 1717 1743
rect 1722 1716 1725 1736
rect 1730 1723 1733 1743
rect 1706 1713 1725 1716
rect 1738 1643 1741 1736
rect 1746 1723 1749 1766
rect 1762 1716 1765 1773
rect 1810 1746 1813 1823
rect 1754 1713 1765 1716
rect 1794 1743 1813 1746
rect 1698 1633 1717 1636
rect 1698 1613 1701 1626
rect 1714 1616 1717 1633
rect 1754 1626 1757 1713
rect 1746 1623 1757 1626
rect 1714 1613 1733 1616
rect 1706 1593 1709 1606
rect 1690 1553 1709 1556
rect 1690 1506 1693 1526
rect 1690 1503 1697 1506
rect 1694 1426 1697 1503
rect 1690 1423 1697 1426
rect 1690 1323 1693 1423
rect 1698 1396 1701 1406
rect 1706 1403 1709 1553
rect 1714 1396 1717 1416
rect 1722 1403 1725 1526
rect 1730 1506 1733 1613
rect 1746 1523 1749 1623
rect 1786 1613 1789 1636
rect 1754 1513 1757 1536
rect 1762 1523 1765 1586
rect 1730 1503 1741 1506
rect 1738 1436 1741 1503
rect 1730 1433 1741 1436
rect 1730 1413 1733 1433
rect 1698 1393 1717 1396
rect 1722 1333 1725 1346
rect 1674 1303 1685 1306
rect 1722 1303 1725 1326
rect 1626 1253 1645 1256
rect 1602 1213 1605 1236
rect 1586 1123 1589 1136
rect 1594 1123 1597 1196
rect 1602 1173 1605 1206
rect 1610 1203 1621 1206
rect 1626 1203 1629 1226
rect 1634 1213 1637 1246
rect 1642 1196 1645 1253
rect 1618 1193 1645 1196
rect 1610 1113 1613 1126
rect 1618 1123 1621 1193
rect 1626 1133 1629 1156
rect 1650 1136 1653 1236
rect 1658 1203 1661 1226
rect 1674 1203 1677 1303
rect 1730 1256 1733 1406
rect 1746 1333 1749 1346
rect 1738 1313 1741 1326
rect 1722 1253 1733 1256
rect 1634 1133 1645 1136
rect 1650 1133 1661 1136
rect 1538 943 1557 946
rect 1530 923 1533 936
rect 1474 733 1485 736
rect 1458 683 1465 686
rect 1450 596 1453 606
rect 1434 593 1453 596
rect 1434 516 1437 526
rect 1450 523 1453 586
rect 1458 563 1461 683
rect 1474 613 1477 726
rect 1482 676 1485 733
rect 1482 673 1493 676
rect 1474 583 1477 606
rect 1490 576 1493 673
rect 1506 583 1509 776
rect 1530 733 1533 796
rect 1538 773 1541 943
rect 1594 936 1597 1106
rect 1634 1096 1637 1126
rect 1626 1093 1637 1096
rect 1626 1036 1629 1093
rect 1626 1033 1637 1036
rect 1634 1013 1637 1033
rect 1642 966 1645 1126
rect 1586 933 1597 936
rect 1626 963 1645 966
rect 1586 856 1589 933
rect 1602 906 1605 926
rect 1626 923 1629 963
rect 1634 916 1637 936
rect 1642 923 1645 956
rect 1650 933 1653 966
rect 1658 923 1661 1133
rect 1666 1123 1669 1136
rect 1690 1133 1693 1146
rect 1698 1123 1701 1216
rect 1706 1133 1709 1156
rect 1674 1003 1677 1026
rect 1690 1003 1693 1076
rect 1634 913 1645 916
rect 1666 913 1669 926
rect 1602 903 1613 906
rect 1586 853 1597 856
rect 1546 813 1549 826
rect 1578 813 1581 836
rect 1586 813 1589 826
rect 1482 573 1493 576
rect 1458 533 1461 546
rect 1466 523 1469 556
rect 1474 523 1477 546
rect 1434 513 1453 516
rect 1450 496 1453 513
rect 1450 493 1461 496
rect 1434 413 1437 436
rect 1442 403 1445 466
rect 1458 436 1461 493
rect 1482 486 1485 573
rect 1522 523 1525 616
rect 1554 613 1557 726
rect 1562 603 1565 616
rect 1578 613 1581 626
rect 1570 593 1573 606
rect 1554 533 1557 586
rect 1586 573 1589 616
rect 1594 556 1597 853
rect 1610 746 1613 903
rect 1626 783 1629 816
rect 1634 796 1637 806
rect 1642 803 1645 913
rect 1674 906 1677 986
rect 1682 936 1685 956
rect 1698 953 1701 1106
rect 1714 1093 1717 1216
rect 1722 1153 1725 1253
rect 1754 1236 1757 1416
rect 1770 1413 1773 1536
rect 1778 1523 1781 1566
rect 1794 1456 1797 1743
rect 1810 1723 1813 1736
rect 1818 1733 1821 1836
rect 1838 1816 1841 1893
rect 1858 1866 1861 1933
rect 1850 1863 1861 1866
rect 1838 1813 1845 1816
rect 1834 1733 1837 1796
rect 1818 1646 1821 1706
rect 1842 1686 1845 1813
rect 1850 1786 1853 1863
rect 1858 1813 1861 1826
rect 1850 1783 1861 1786
rect 1858 1726 1861 1783
rect 1850 1723 1861 1726
rect 1850 1703 1853 1723
rect 1842 1683 1861 1686
rect 1786 1453 1797 1456
rect 1810 1643 1821 1646
rect 1786 1376 1789 1453
rect 1810 1393 1813 1643
rect 1834 1573 1837 1606
rect 1786 1373 1797 1376
rect 1762 1296 1765 1316
rect 1762 1293 1769 1296
rect 1746 1233 1757 1236
rect 1746 1216 1749 1233
rect 1766 1226 1769 1293
rect 1742 1213 1749 1216
rect 1742 1156 1745 1213
rect 1742 1153 1749 1156
rect 1730 1123 1733 1146
rect 1746 1016 1749 1153
rect 1754 1133 1757 1226
rect 1762 1223 1769 1226
rect 1762 1203 1765 1223
rect 1778 1213 1781 1316
rect 1786 1203 1789 1216
rect 1794 1186 1797 1373
rect 1818 1313 1821 1326
rect 1826 1226 1829 1556
rect 1850 1553 1853 1676
rect 1858 1666 1861 1683
rect 1858 1663 1865 1666
rect 1862 1546 1865 1663
rect 1874 1613 1877 1726
rect 1882 1676 1885 1926
rect 1906 1916 1909 1983
rect 1898 1913 1909 1916
rect 1898 1846 1901 1913
rect 1898 1843 1909 1846
rect 1898 1813 1901 1826
rect 1898 1766 1901 1806
rect 1890 1763 1901 1766
rect 1890 1723 1893 1763
rect 1898 1683 1901 1736
rect 1906 1733 1909 1843
rect 1882 1673 1893 1676
rect 1890 1576 1893 1673
rect 1906 1643 1909 1726
rect 1914 1723 1917 2003
rect 1922 1996 1925 2026
rect 1938 2013 1941 2033
rect 1922 1993 1933 1996
rect 1930 1776 1933 1993
rect 1946 1913 1949 1926
rect 1954 1923 1957 2006
rect 1970 1936 1973 2216
rect 1978 2193 1981 2346
rect 1986 2166 1989 2216
rect 2002 2213 2005 2756
rect 2010 2743 2029 2746
rect 2010 2733 2013 2743
rect 2018 2673 2021 2736
rect 2026 2723 2029 2743
rect 2034 2733 2037 2746
rect 2050 2723 2053 2933
rect 2058 2923 2061 2993
rect 2074 2983 2077 3006
rect 2066 2923 2069 2936
rect 2074 2856 2077 2976
rect 2082 2913 2085 2996
rect 2074 2853 2081 2856
rect 2058 2813 2061 2826
rect 2078 2776 2081 2853
rect 2090 2813 2093 3006
rect 2106 2933 2109 2956
rect 2114 2933 2117 3013
rect 2098 2846 2101 2926
rect 2098 2843 2109 2846
rect 2098 2813 2101 2826
rect 2106 2806 2109 2843
rect 2098 2803 2109 2806
rect 2074 2773 2081 2776
rect 2018 2613 2021 2626
rect 2010 2583 2013 2606
rect 2034 2593 2037 2616
rect 2058 2613 2061 2626
rect 2010 2513 2013 2526
rect 2066 2523 2069 2726
rect 2074 2543 2077 2773
rect 2098 2666 2101 2786
rect 2106 2733 2109 2796
rect 2082 2663 2101 2666
rect 2082 2576 2085 2663
rect 2114 2653 2117 2926
rect 2122 2873 2125 2976
rect 2106 2613 2117 2616
rect 2122 2613 2125 2806
rect 2130 2783 2133 3063
rect 2138 2973 2141 3116
rect 2162 3046 2165 3123
rect 2186 3113 2189 3326
rect 2194 3203 2197 3426
rect 2202 3323 2205 3416
rect 2210 3333 2213 3396
rect 2202 3276 2205 3296
rect 2202 3273 2209 3276
rect 2218 3273 2221 3583
rect 2242 3576 2245 3606
rect 2226 3573 2245 3576
rect 2226 3503 2229 3573
rect 2226 3323 2229 3336
rect 2206 3196 2209 3273
rect 2202 3193 2209 3196
rect 2202 3166 2205 3193
rect 2198 3163 2205 3166
rect 2198 3046 2201 3163
rect 2146 3043 2165 3046
rect 2146 2986 2149 3043
rect 2154 3013 2157 3026
rect 2178 3003 2181 3046
rect 2198 3043 2205 3046
rect 2194 3013 2197 3026
rect 2146 2983 2157 2986
rect 2138 2813 2141 2936
rect 2154 2836 2157 2983
rect 2170 2923 2173 2976
rect 2194 2973 2197 3006
rect 2146 2833 2157 2836
rect 2106 2606 2109 2613
rect 2130 2606 2133 2736
rect 2146 2706 2149 2833
rect 2170 2733 2173 2816
rect 2178 2803 2181 2956
rect 2194 2893 2197 2936
rect 2202 2923 2205 3043
rect 2186 2753 2189 2816
rect 2210 2763 2213 3156
rect 2218 2893 2221 3216
rect 2234 3153 2237 3526
rect 2250 3523 2253 3696
rect 2258 3566 2261 3726
rect 2266 3603 2269 3926
rect 2274 3723 2277 3916
rect 2258 3563 2269 3566
rect 2266 3546 2269 3563
rect 2266 3543 2277 3546
rect 2242 3486 2245 3506
rect 2274 3493 2277 3543
rect 2242 3483 2249 3486
rect 2282 3483 2285 4026
rect 2290 4003 2293 4016
rect 2290 3913 2293 3926
rect 2290 3813 2293 3826
rect 2290 3603 2293 3806
rect 2298 3706 2301 4046
rect 2306 4003 2309 4216
rect 2314 4203 2317 4216
rect 2330 4113 2333 4216
rect 2338 4186 2341 4336
rect 2378 4333 2381 4343
rect 2354 4303 2357 4326
rect 2346 4203 2349 4296
rect 2354 4213 2357 4256
rect 2362 4203 2365 4266
rect 2338 4183 2349 4186
rect 2346 4106 2349 4183
rect 2386 4166 2389 4336
rect 2402 4323 2405 4353
rect 2426 4333 2429 4416
rect 2458 4413 2461 4426
rect 2434 4333 2437 4366
rect 2506 4346 2509 4406
rect 2522 4396 2525 4536
rect 2530 4523 2533 4606
rect 2554 4436 2557 4606
rect 2570 4533 2573 4546
rect 2578 4523 2581 4536
rect 2586 4523 2589 4536
rect 2594 4513 2597 4526
rect 2602 4523 2605 4536
rect 2634 4456 2637 4616
rect 2674 4613 2677 4626
rect 2714 4613 2717 4626
rect 2642 4523 2645 4536
rect 2650 4523 2653 4606
rect 2690 4593 2693 4606
rect 2634 4453 2645 4456
rect 2554 4433 2581 4436
rect 2562 4413 2565 4426
rect 2522 4393 2533 4396
rect 2338 4103 2349 4106
rect 2378 4163 2389 4166
rect 2338 4023 2341 4103
rect 2370 4013 2373 4046
rect 2306 3913 2309 3936
rect 2314 3923 2317 3996
rect 2322 3933 2325 3956
rect 2330 3943 2349 3946
rect 2330 3923 2333 3943
rect 2338 3913 2341 3936
rect 2346 3933 2349 3943
rect 2354 3906 2357 4006
rect 2370 3993 2373 4006
rect 2378 3936 2381 4163
rect 2402 4123 2405 4256
rect 2434 4226 2437 4326
rect 2466 4253 2469 4326
rect 2474 4303 2477 4336
rect 2490 4333 2493 4346
rect 2506 4343 2517 4346
rect 2434 4223 2445 4226
rect 2410 4123 2413 4136
rect 2418 4113 2421 4216
rect 2338 3903 2357 3906
rect 2370 3933 2381 3936
rect 2394 3936 2397 4016
rect 2410 4003 2413 4106
rect 2426 4086 2429 4136
rect 2442 4126 2445 4223
rect 2482 4213 2485 4326
rect 2498 4266 2501 4336
rect 2494 4263 2501 4266
rect 2494 4156 2497 4263
rect 2514 4256 2517 4343
rect 2506 4253 2517 4256
rect 2494 4153 2501 4156
rect 2434 4123 2445 4126
rect 2434 4103 2437 4123
rect 2474 4113 2477 4136
rect 2482 4133 2493 4136
rect 2498 4116 2501 4153
rect 2490 4113 2501 4116
rect 2426 4083 2437 4086
rect 2434 4036 2437 4083
rect 2426 4033 2437 4036
rect 2490 4036 2493 4113
rect 2506 4096 2509 4253
rect 2530 4236 2533 4393
rect 2538 4376 2541 4406
rect 2538 4373 2549 4376
rect 2546 4323 2549 4373
rect 2578 4336 2581 4433
rect 2602 4413 2605 4426
rect 2642 4403 2645 4453
rect 2562 4276 2565 4336
rect 2578 4333 2589 4336
rect 2602 4333 2605 4346
rect 2618 4343 2637 4346
rect 2658 4343 2661 4416
rect 2666 4406 2669 4536
rect 2674 4533 2677 4576
rect 2674 4483 2677 4526
rect 2682 4523 2685 4546
rect 2690 4436 2693 4526
rect 2698 4523 2701 4536
rect 2706 4523 2709 4536
rect 2714 4533 2717 4546
rect 2714 4473 2717 4526
rect 2730 4523 2733 4596
rect 2778 4573 2781 4606
rect 2754 4543 2757 4556
rect 2746 4523 2749 4536
rect 2762 4533 2765 4546
rect 2778 4493 2781 4536
rect 2682 4433 2693 4436
rect 2786 4436 2789 4536
rect 2794 4533 2797 4706
rect 2810 4556 2813 4606
rect 2818 4593 2821 4606
rect 2826 4563 2829 4626
rect 2850 4613 2853 4626
rect 2802 4553 2813 4556
rect 2802 4523 2805 4553
rect 2842 4543 2845 4576
rect 2810 4523 2813 4536
rect 2826 4506 2829 4536
rect 2842 4526 2845 4536
rect 2850 4533 2853 4556
rect 2858 4533 2861 4616
rect 2874 4573 2877 4646
rect 2890 4613 2893 4626
rect 2938 4583 2941 4606
rect 2986 4593 2989 4606
rect 3034 4603 3037 4616
rect 2842 4523 2861 4526
rect 2866 4523 2869 4536
rect 2834 4513 2845 4516
rect 2826 4503 2837 4506
rect 2834 4436 2837 4503
rect 2914 4466 2917 4536
rect 2930 4486 2933 4516
rect 2938 4503 2941 4516
rect 2970 4513 2973 4536
rect 2978 4533 2981 4566
rect 3002 4533 3005 4546
rect 2978 4523 2997 4526
rect 2930 4483 2941 4486
rect 2906 4463 2917 4466
rect 2786 4433 2797 4436
rect 2834 4433 2841 4436
rect 2850 4433 2861 4436
rect 2666 4403 2677 4406
rect 2682 4403 2685 4433
rect 2698 4413 2701 4426
rect 2738 4413 2741 4426
rect 2794 4413 2797 4433
rect 2570 4283 2573 4326
rect 2562 4273 2573 4276
rect 2522 4233 2533 4236
rect 2522 4186 2525 4233
rect 2522 4183 2533 4186
rect 2514 4123 2517 4136
rect 2530 4106 2533 4183
rect 2538 4173 2541 4206
rect 2562 4133 2565 4216
rect 2538 4113 2541 4126
rect 2530 4103 2557 4106
rect 2570 4103 2573 4273
rect 2586 4266 2589 4333
rect 2578 4263 2589 4266
rect 2578 4173 2581 4263
rect 2506 4093 2517 4096
rect 2490 4033 2501 4036
rect 2426 4013 2429 4033
rect 2394 3933 2413 3936
rect 2306 3796 2309 3816
rect 2314 3803 2317 3816
rect 2322 3813 2325 3846
rect 2338 3826 2341 3903
rect 2338 3823 2345 3826
rect 2322 3796 2325 3806
rect 2306 3793 2325 3796
rect 2306 3733 2309 3746
rect 2314 3723 2317 3786
rect 2330 3733 2333 3816
rect 2342 3726 2345 3823
rect 2354 3733 2357 3816
rect 2338 3723 2345 3726
rect 2298 3703 2309 3706
rect 2306 3636 2309 3703
rect 2298 3633 2309 3636
rect 2322 3636 2325 3656
rect 2322 3633 2329 3636
rect 2290 3513 2293 3526
rect 2246 3376 2249 3483
rect 2242 3373 2249 3376
rect 2242 3353 2245 3373
rect 2258 3356 2261 3416
rect 2282 3363 2285 3406
rect 2298 3376 2301 3633
rect 2294 3373 2301 3376
rect 2258 3353 2269 3356
rect 2242 3343 2261 3346
rect 2242 3323 2245 3343
rect 2250 3203 2253 3336
rect 2258 3333 2261 3343
rect 2258 3313 2261 3326
rect 2266 3323 2269 3353
rect 2294 3286 2297 3373
rect 2306 3293 2309 3416
rect 2294 3283 2301 3286
rect 2266 3216 2269 3246
rect 2258 3213 2269 3216
rect 2274 3203 2277 3266
rect 2282 3213 2285 3276
rect 2234 3043 2237 3136
rect 2258 3076 2261 3116
rect 2250 3073 2261 3076
rect 2226 2993 2229 3036
rect 2250 2986 2253 3073
rect 2266 3013 2269 3126
rect 2258 2993 2261 3006
rect 2250 2983 2261 2986
rect 2234 2856 2237 2936
rect 2258 2933 2261 2983
rect 2258 2896 2261 2926
rect 2274 2913 2277 3016
rect 2282 3003 2285 3026
rect 2290 3003 2293 3066
rect 2298 2966 2301 3283
rect 2314 3216 2317 3616
rect 2326 3546 2329 3633
rect 2338 3613 2341 3723
rect 2354 3713 2365 3716
rect 2362 3696 2365 3713
rect 2354 3693 2365 3696
rect 2354 3636 2357 3693
rect 2354 3633 2365 3636
rect 2362 3613 2365 3633
rect 2322 3543 2329 3546
rect 2322 3523 2325 3543
rect 2330 3503 2333 3526
rect 2338 3513 2341 3526
rect 2346 3496 2349 3606
rect 2370 3556 2373 3933
rect 2378 3896 2381 3916
rect 2378 3893 2389 3896
rect 2386 3836 2389 3893
rect 2378 3833 2389 3836
rect 2378 3813 2381 3833
rect 2426 3813 2429 3926
rect 2482 3923 2485 4016
rect 2498 3946 2501 4033
rect 2506 3966 2509 4093
rect 2546 4013 2549 4046
rect 2530 3993 2533 4006
rect 2506 3963 2517 3966
rect 2490 3943 2501 3946
rect 2490 3906 2493 3943
rect 2498 3913 2501 3936
rect 2514 3906 2517 3963
rect 2482 3903 2493 3906
rect 2506 3903 2517 3906
rect 2482 3846 2485 3903
rect 2482 3843 2493 3846
rect 2458 3803 2461 3816
rect 2402 3723 2405 3736
rect 2378 3613 2381 3656
rect 2418 3613 2421 3646
rect 2426 3636 2429 3706
rect 2450 3693 2453 3736
rect 2466 3703 2469 3726
rect 2426 3633 2445 3636
rect 2426 3613 2429 3626
rect 2370 3553 2381 3556
rect 2354 3543 2373 3546
rect 2354 3533 2357 3543
rect 2322 3413 2325 3496
rect 2330 3493 2349 3496
rect 2330 3403 2333 3493
rect 2354 3483 2357 3526
rect 2346 3393 2349 3406
rect 2330 3333 2333 3366
rect 2354 3353 2357 3416
rect 2362 3403 2365 3536
rect 2370 3523 2373 3543
rect 2378 3413 2381 3553
rect 2386 3536 2389 3606
rect 2418 3563 2421 3606
rect 2434 3603 2437 3616
rect 2386 3533 2397 3536
rect 2386 3513 2389 3526
rect 2394 3523 2397 3533
rect 2402 3443 2405 3506
rect 2410 3483 2413 3556
rect 2314 3213 2325 3216
rect 2306 3126 2309 3206
rect 2322 3166 2325 3213
rect 2338 3203 2341 3226
rect 2354 3213 2357 3326
rect 2370 3316 2373 3336
rect 2362 3213 2365 3316
rect 2370 3313 2377 3316
rect 2374 3216 2377 3313
rect 2402 3283 2405 3416
rect 2418 3403 2421 3536
rect 2426 3506 2429 3576
rect 2434 3533 2437 3586
rect 2442 3573 2445 3633
rect 2450 3553 2453 3616
rect 2466 3613 2469 3626
rect 2474 3613 2477 3816
rect 2490 3796 2493 3843
rect 2498 3813 2501 3826
rect 2506 3813 2509 3903
rect 2522 3803 2525 3846
rect 2490 3793 2501 3796
rect 2498 3666 2501 3793
rect 2530 3733 2533 3936
rect 2554 3933 2557 4103
rect 2538 3893 2541 3926
rect 2546 3853 2549 3926
rect 2562 3913 2565 3926
rect 2578 3836 2581 4006
rect 2586 3896 2589 4236
rect 2610 4226 2613 4336
rect 2618 4323 2621 4343
rect 2626 4323 2629 4336
rect 2634 4333 2637 4343
rect 2642 4323 2645 4336
rect 2610 4223 2629 4226
rect 2594 4133 2597 4156
rect 2602 4116 2605 4136
rect 2598 4113 2605 4116
rect 2598 4036 2601 4113
rect 2598 4033 2605 4036
rect 2594 4003 2597 4016
rect 2602 4013 2605 4033
rect 2594 3913 2597 3936
rect 2586 3893 2597 3896
rect 2570 3833 2581 3836
rect 2538 3796 2541 3816
rect 2546 3803 2549 3816
rect 2554 3796 2557 3806
rect 2538 3793 2557 3796
rect 2546 3716 2549 3736
rect 2562 3716 2565 3736
rect 2570 3733 2573 3833
rect 2594 3826 2597 3893
rect 2610 3886 2613 4176
rect 2618 4153 2621 4216
rect 2626 4203 2629 4223
rect 2634 4213 2637 4236
rect 2658 4196 2661 4216
rect 2666 4203 2669 4216
rect 2674 4213 2677 4403
rect 2714 4366 2717 4406
rect 2802 4383 2805 4406
rect 2826 4396 2829 4426
rect 2818 4393 2829 4396
rect 2706 4363 2717 4366
rect 2690 4323 2693 4336
rect 2706 4283 2709 4363
rect 2794 4343 2797 4376
rect 2818 4336 2821 4393
rect 2838 4386 2841 4433
rect 2834 4383 2841 4386
rect 2730 4323 2733 4336
rect 2818 4333 2829 4336
rect 2778 4323 2789 4326
rect 2738 4213 2741 4226
rect 2674 4196 2677 4206
rect 2658 4193 2677 4196
rect 2754 4176 2757 4286
rect 2826 4253 2829 4333
rect 2834 4236 2837 4383
rect 2842 4293 2845 4346
rect 2850 4323 2853 4406
rect 2858 4393 2861 4433
rect 2874 4423 2877 4436
rect 2898 4403 2901 4446
rect 2906 4413 2909 4463
rect 2938 4436 2941 4483
rect 2930 4433 2941 4436
rect 2914 4413 2917 4426
rect 2930 4413 2933 4433
rect 2962 4423 2965 4476
rect 2978 4466 2981 4516
rect 2970 4463 2981 4466
rect 2970 4423 2973 4463
rect 2986 4413 2989 4523
rect 3010 4473 3013 4536
rect 3042 4523 3061 4526
rect 3018 4456 3021 4516
rect 3074 4476 3077 4536
rect 3082 4506 3085 4536
rect 3090 4513 3093 4616
rect 3098 4533 3101 4606
rect 3122 4586 3125 4736
rect 3122 4583 3133 4586
rect 3130 4533 3133 4583
rect 3098 4506 3101 4526
rect 3082 4503 3101 4506
rect 3074 4473 3093 4476
rect 2906 4403 2917 4406
rect 2858 4306 2861 4336
rect 2866 4333 2869 4376
rect 2874 4323 2877 4336
rect 2890 4323 2893 4346
rect 2922 4333 2925 4346
rect 2930 4343 2933 4356
rect 2858 4303 2869 4306
rect 2866 4256 2869 4303
rect 2826 4233 2837 4236
rect 2778 4213 2781 4226
rect 2826 4186 2829 4233
rect 2842 4213 2845 4226
rect 2842 4193 2845 4206
rect 2826 4183 2837 4186
rect 2634 4133 2637 4176
rect 2746 4173 2757 4176
rect 2722 4133 2725 4146
rect 2618 4113 2621 4126
rect 2658 4113 2661 4126
rect 2618 4003 2621 4106
rect 2626 3983 2629 4016
rect 2666 4003 2669 4026
rect 2714 4023 2717 4126
rect 2746 4116 2749 4173
rect 2834 4166 2837 4183
rect 2850 4166 2853 4256
rect 2858 4253 2869 4256
rect 2858 4233 2861 4253
rect 2826 4163 2837 4166
rect 2846 4163 2853 4166
rect 2770 4123 2773 4146
rect 2746 4113 2757 4116
rect 2674 4003 2677 4016
rect 2690 3996 2693 4016
rect 2698 4003 2701 4016
rect 2706 3996 2709 4006
rect 2714 4003 2717 4016
rect 2690 3993 2709 3996
rect 2634 3893 2637 3926
rect 2690 3913 2693 3926
rect 2610 3883 2629 3886
rect 2586 3823 2597 3826
rect 2490 3663 2501 3666
rect 2538 3713 2549 3716
rect 2558 3713 2565 3716
rect 2570 3713 2573 3726
rect 2490 3636 2493 3663
rect 2538 3646 2541 3713
rect 2538 3643 2549 3646
rect 2482 3633 2493 3636
rect 2442 3523 2445 3536
rect 2426 3503 2437 3506
rect 2434 3416 2437 3503
rect 2450 3453 2453 3526
rect 2458 3523 2461 3536
rect 2466 3523 2469 3566
rect 2474 3533 2477 3606
rect 2482 3583 2485 3633
rect 2482 3506 2485 3576
rect 2474 3503 2485 3506
rect 2426 3413 2437 3416
rect 2426 3393 2429 3413
rect 2450 3376 2453 3406
rect 2450 3373 2461 3376
rect 2394 3253 2405 3256
rect 2370 3213 2377 3216
rect 2314 3163 2325 3166
rect 2314 3136 2317 3163
rect 2314 3133 2325 3136
rect 2306 3123 2317 3126
rect 2306 3063 2309 3123
rect 2306 3016 2309 3026
rect 2306 3013 2317 3016
rect 2298 2963 2305 2966
rect 2226 2853 2237 2856
rect 2098 2603 2109 2606
rect 2114 2603 2133 2606
rect 2138 2703 2149 2706
rect 2082 2573 2093 2576
rect 2090 2506 2093 2573
rect 2082 2503 2093 2506
rect 2082 2446 2085 2503
rect 2082 2443 2093 2446
rect 2018 2353 2021 2406
rect 2058 2326 2061 2406
rect 2066 2383 2069 2416
rect 2090 2413 2093 2443
rect 2082 2383 2085 2406
rect 2098 2403 2101 2603
rect 2026 2303 2029 2326
rect 2050 2323 2061 2326
rect 2066 2303 2069 2326
rect 2114 2256 2117 2603
rect 2130 2533 2133 2566
rect 2138 2273 2141 2703
rect 2178 2613 2181 2726
rect 2202 2603 2205 2616
rect 2226 2593 2229 2853
rect 2250 2836 2253 2896
rect 2258 2893 2269 2896
rect 2242 2833 2253 2836
rect 2242 2776 2245 2833
rect 2266 2826 2269 2893
rect 2302 2886 2305 2963
rect 2262 2823 2269 2826
rect 2298 2883 2305 2886
rect 2242 2773 2249 2776
rect 2234 2733 2237 2756
rect 2246 2656 2249 2773
rect 2262 2756 2265 2823
rect 2258 2753 2265 2756
rect 2258 2723 2261 2753
rect 2266 2716 2269 2736
rect 2258 2713 2269 2716
rect 2246 2653 2253 2656
rect 2154 2523 2157 2536
rect 2162 2343 2181 2346
rect 2162 2333 2165 2343
rect 2114 2253 2125 2256
rect 2050 2213 2053 2226
rect 2002 2193 2005 2206
rect 1986 2163 1997 2166
rect 1994 2056 1997 2163
rect 1986 2053 1997 2056
rect 1962 1933 1973 1936
rect 1962 1906 1965 1933
rect 1958 1903 1965 1906
rect 1958 1826 1961 1903
rect 1946 1803 1949 1826
rect 1954 1823 1961 1826
rect 1970 1823 1973 1926
rect 1978 1886 1981 1956
rect 1986 1923 1989 2053
rect 2026 2013 2029 2026
rect 2010 1933 2013 1946
rect 1994 1906 1997 1926
rect 2018 1923 2021 2006
rect 2034 2003 2037 2136
rect 2058 2133 2061 2146
rect 2082 2133 2085 2216
rect 2090 2213 2093 2226
rect 2106 2213 2109 2246
rect 2122 2206 2125 2253
rect 2162 2213 2165 2326
rect 2170 2323 2173 2336
rect 2178 2323 2181 2343
rect 2194 2323 2197 2436
rect 2114 2203 2125 2206
rect 2050 2116 2053 2126
rect 2058 2123 2069 2126
rect 2042 2113 2053 2116
rect 2050 2093 2053 2113
rect 2042 1963 2045 2016
rect 2050 1943 2053 2006
rect 2058 1986 2061 2006
rect 2058 1983 2069 1986
rect 2050 1913 2053 1926
rect 1994 1903 2005 1906
rect 1978 1883 1989 1886
rect 1986 1836 1989 1883
rect 1978 1833 1989 1836
rect 1954 1786 1957 1823
rect 1926 1773 1933 1776
rect 1950 1783 1957 1786
rect 1926 1716 1929 1773
rect 1922 1713 1929 1716
rect 1950 1716 1953 1783
rect 1962 1723 1965 1816
rect 1978 1813 1981 1833
rect 2002 1806 2005 1903
rect 2066 1886 2069 1983
rect 2114 1956 2117 2203
rect 2170 2196 2173 2206
rect 2178 2203 2181 2216
rect 2186 2196 2189 2216
rect 2170 2193 2189 2196
rect 2162 2133 2165 2166
rect 2146 2013 2149 2126
rect 2178 2046 2181 2136
rect 2186 2093 2189 2126
rect 2202 2123 2205 2216
rect 2210 2193 2213 2336
rect 2218 2323 2221 2586
rect 2234 2446 2237 2466
rect 2230 2443 2237 2446
rect 2230 2326 2233 2443
rect 2242 2333 2245 2596
rect 2250 2583 2253 2653
rect 2258 2533 2261 2713
rect 2274 2636 2277 2806
rect 2282 2713 2285 2816
rect 2298 2766 2301 2883
rect 2294 2763 2301 2766
rect 2294 2716 2297 2763
rect 2306 2723 2309 2756
rect 2314 2733 2317 2926
rect 2322 2886 2325 3133
rect 2330 3013 2333 3036
rect 2330 2953 2333 3006
rect 2338 2903 2341 3136
rect 2346 2956 2349 3066
rect 2362 3013 2365 3126
rect 2370 3033 2373 3213
rect 2386 3203 2389 3216
rect 2394 3213 2397 3226
rect 2402 3203 2405 3253
rect 2378 3176 2381 3196
rect 2410 3186 2413 3226
rect 2418 3213 2421 3326
rect 2426 3213 2429 3276
rect 2406 3183 2413 3186
rect 2378 3173 2385 3176
rect 2382 3046 2385 3173
rect 2378 3043 2385 3046
rect 2378 3026 2381 3043
rect 2406 3036 2409 3183
rect 2406 3033 2413 3036
rect 2370 3023 2381 3026
rect 2370 3013 2373 3023
rect 2354 3003 2365 3006
rect 2370 2973 2373 3006
rect 2386 3003 2389 3016
rect 2394 2973 2397 3016
rect 2346 2953 2357 2956
rect 2354 2896 2357 2953
rect 2346 2893 2357 2896
rect 2322 2883 2333 2886
rect 2330 2756 2333 2883
rect 2322 2753 2333 2756
rect 2322 2733 2325 2753
rect 2294 2713 2301 2716
rect 2266 2633 2277 2636
rect 2266 2593 2269 2633
rect 2298 2626 2301 2713
rect 2274 2613 2277 2626
rect 2294 2623 2301 2626
rect 2294 2556 2297 2623
rect 2306 2573 2309 2616
rect 2314 2566 2317 2716
rect 2322 2683 2325 2726
rect 2346 2696 2349 2893
rect 2362 2803 2365 2816
rect 2378 2813 2381 2956
rect 2402 2866 2405 3016
rect 2410 2936 2413 3033
rect 2418 3013 2421 3206
rect 2434 3193 2437 3366
rect 2458 3306 2461 3373
rect 2450 3303 2461 3306
rect 2426 3136 2429 3156
rect 2426 3133 2433 3136
rect 2430 3046 2433 3133
rect 2442 3063 2445 3276
rect 2430 3043 2437 3046
rect 2418 2953 2421 3006
rect 2434 2946 2437 3043
rect 2426 2943 2437 2946
rect 2410 2933 2417 2936
rect 2394 2863 2405 2866
rect 2370 2753 2373 2806
rect 2338 2693 2349 2696
rect 2338 2626 2341 2693
rect 2322 2613 2325 2626
rect 2338 2623 2345 2626
rect 2306 2563 2317 2566
rect 2294 2553 2301 2556
rect 2290 2506 2293 2536
rect 2282 2503 2293 2506
rect 2250 2433 2253 2466
rect 2282 2446 2285 2503
rect 2282 2443 2293 2446
rect 2250 2386 2253 2416
rect 2274 2413 2277 2426
rect 2290 2413 2293 2443
rect 2298 2403 2301 2553
rect 2306 2523 2309 2563
rect 2314 2516 2317 2536
rect 2322 2523 2325 2606
rect 2330 2533 2333 2606
rect 2342 2556 2345 2623
rect 2342 2553 2349 2556
rect 2306 2513 2317 2516
rect 2250 2383 2261 2386
rect 2258 2336 2261 2383
rect 2282 2363 2285 2386
rect 2290 2383 2301 2386
rect 2250 2333 2261 2336
rect 2290 2333 2293 2383
rect 2306 2333 2309 2513
rect 2230 2323 2237 2326
rect 2234 2146 2237 2323
rect 2250 2283 2253 2333
rect 2314 2316 2317 2496
rect 2266 2236 2269 2316
rect 2258 2233 2269 2236
rect 2306 2313 2317 2316
rect 2306 2236 2309 2313
rect 2306 2233 2317 2236
rect 2258 2156 2261 2233
rect 2274 2203 2277 2226
rect 2258 2153 2269 2156
rect 2226 2143 2237 2146
rect 2226 2066 2229 2143
rect 2226 2063 2233 2066
rect 2178 2043 2197 2046
rect 2114 1953 2125 1956
rect 2098 1923 2101 1936
rect 2122 1906 2125 1953
rect 2162 1923 2165 2006
rect 2178 1926 2181 1986
rect 2194 1966 2197 2043
rect 2186 1963 2197 1966
rect 2186 1943 2189 1963
rect 2210 1953 2213 2016
rect 2230 1986 2233 2063
rect 2230 1983 2237 1986
rect 2178 1923 2189 1926
rect 1994 1803 2005 1806
rect 2042 1883 2069 1886
rect 2114 1903 2125 1906
rect 1950 1713 1957 1716
rect 1890 1573 1901 1576
rect 1858 1543 1865 1546
rect 1858 1443 1861 1543
rect 1874 1513 1877 1526
rect 1834 1413 1837 1426
rect 1858 1403 1861 1416
rect 1874 1413 1877 1426
rect 1842 1346 1845 1396
rect 1898 1366 1901 1573
rect 1906 1556 1909 1616
rect 1914 1563 1917 1606
rect 1922 1593 1925 1713
rect 1930 1683 1941 1686
rect 1906 1553 1925 1556
rect 1914 1513 1917 1526
rect 1922 1496 1925 1553
rect 1930 1533 1933 1616
rect 1938 1603 1941 1683
rect 1954 1676 1957 1713
rect 1954 1673 1961 1676
rect 1946 1586 1949 1666
rect 1958 1626 1961 1673
rect 1942 1583 1949 1586
rect 1954 1623 1961 1626
rect 1914 1493 1925 1496
rect 1914 1436 1917 1493
rect 1914 1433 1925 1436
rect 1922 1413 1925 1433
rect 1898 1363 1909 1366
rect 1838 1343 1845 1346
rect 1838 1296 1841 1343
rect 1866 1333 1869 1356
rect 1838 1293 1845 1296
rect 1822 1223 1829 1226
rect 1786 1183 1797 1186
rect 1754 1103 1757 1126
rect 1682 933 1689 936
rect 1666 903 1677 906
rect 1650 796 1653 816
rect 1666 813 1669 903
rect 1686 856 1689 933
rect 1698 873 1701 936
rect 1706 913 1709 936
rect 1714 906 1717 1016
rect 1746 1013 1757 1016
rect 1706 903 1717 906
rect 1686 853 1693 856
rect 1674 813 1677 846
rect 1690 806 1693 853
rect 1634 793 1653 796
rect 1602 743 1613 746
rect 1602 576 1605 743
rect 1626 733 1629 756
rect 1610 713 1613 726
rect 1618 693 1621 726
rect 1618 613 1621 626
rect 1634 613 1637 726
rect 1642 713 1645 736
rect 1650 723 1653 786
rect 1658 753 1661 806
rect 1682 803 1693 806
rect 1706 803 1709 903
rect 1722 863 1725 936
rect 1730 903 1733 926
rect 1682 713 1685 803
rect 1730 796 1733 816
rect 1738 803 1741 936
rect 1746 923 1749 1006
rect 1754 976 1757 1013
rect 1762 996 1765 1016
rect 1770 1003 1773 1156
rect 1786 1116 1789 1183
rect 1802 1123 1805 1206
rect 1822 1156 1825 1223
rect 1822 1153 1829 1156
rect 1826 1133 1829 1153
rect 1834 1123 1837 1216
rect 1842 1166 1845 1293
rect 1882 1213 1885 1326
rect 1890 1206 1893 1356
rect 1906 1266 1909 1363
rect 1930 1336 1933 1526
rect 1942 1516 1945 1583
rect 1954 1523 1957 1623
rect 1942 1513 1949 1516
rect 1946 1453 1949 1513
rect 1962 1423 1965 1606
rect 1970 1533 1973 1756
rect 1994 1733 1997 1803
rect 1994 1613 1997 1716
rect 2010 1696 2013 1746
rect 2026 1713 2029 1746
rect 2006 1693 2013 1696
rect 2006 1626 2009 1693
rect 2006 1623 2013 1626
rect 2010 1603 2013 1623
rect 2018 1603 2021 1696
rect 2042 1663 2045 1883
rect 2114 1826 2117 1903
rect 2162 1876 2165 1896
rect 2162 1873 2169 1876
rect 2050 1813 2053 1826
rect 2098 1823 2117 1826
rect 2058 1813 2069 1816
rect 2066 1733 2069 1806
rect 2098 1726 2101 1823
rect 2122 1736 2125 1816
rect 2130 1773 2133 1826
rect 2122 1733 2141 1736
rect 2146 1733 2149 1816
rect 2058 1713 2061 1726
rect 2074 1703 2077 1726
rect 2098 1723 2117 1726
rect 2114 1653 2117 1723
rect 2130 1713 2133 1726
rect 2154 1723 2157 1856
rect 2166 1716 2169 1873
rect 2186 1836 2189 1923
rect 2162 1713 2169 1716
rect 2178 1833 2189 1836
rect 2002 1483 2005 1526
rect 2018 1523 2021 1536
rect 2026 1523 2029 1646
rect 2090 1536 2093 1616
rect 2146 1603 2149 1656
rect 2162 1596 2165 1713
rect 2090 1533 2097 1536
rect 1866 1193 1869 1206
rect 1882 1203 1893 1206
rect 1898 1263 1909 1266
rect 1922 1333 1933 1336
rect 1882 1166 1885 1203
rect 1898 1176 1901 1263
rect 1922 1206 1925 1333
rect 1938 1213 1941 1326
rect 1962 1323 1965 1416
rect 1970 1396 1973 1406
rect 1978 1403 1981 1436
rect 1986 1396 1989 1416
rect 1994 1403 1997 1426
rect 2002 1413 2005 1476
rect 2034 1436 2037 1456
rect 2030 1433 2037 1436
rect 1970 1393 1989 1396
rect 1994 1343 2013 1346
rect 1994 1333 1997 1343
rect 1922 1203 1933 1206
rect 1842 1163 1853 1166
rect 1850 1116 1853 1163
rect 1786 1113 1813 1116
rect 1778 1013 1781 1056
rect 1810 1026 1813 1113
rect 1842 1113 1853 1116
rect 1874 1163 1885 1166
rect 1894 1173 1901 1176
rect 1842 1036 1845 1113
rect 1874 1086 1877 1163
rect 1894 1116 1897 1173
rect 1906 1143 1925 1146
rect 1906 1133 1909 1143
rect 1894 1113 1901 1116
rect 1898 1096 1901 1113
rect 1906 1103 1909 1126
rect 1914 1123 1917 1136
rect 1922 1123 1925 1143
rect 1930 1113 1933 1203
rect 1962 1193 1965 1206
rect 1938 1143 1965 1146
rect 1938 1133 1941 1143
rect 1898 1093 1917 1096
rect 1938 1093 1941 1126
rect 1874 1083 1885 1086
rect 1842 1033 1849 1036
rect 1802 1023 1813 1026
rect 1778 996 1781 1006
rect 1762 993 1781 996
rect 1754 973 1765 976
rect 1762 836 1765 973
rect 1802 886 1805 1023
rect 1826 976 1829 1016
rect 1834 1013 1837 1026
rect 1826 973 1837 976
rect 1834 923 1837 973
rect 1846 966 1849 1033
rect 1846 963 1853 966
rect 1850 916 1853 963
rect 1842 913 1853 916
rect 1802 883 1813 886
rect 1754 833 1765 836
rect 1746 796 1749 806
rect 1730 793 1749 796
rect 1690 733 1693 746
rect 1690 723 1701 726
rect 1706 723 1709 736
rect 1730 733 1733 746
rect 1738 736 1741 756
rect 1738 733 1749 736
rect 1690 613 1693 723
rect 1666 583 1669 606
rect 1602 573 1613 576
rect 1594 553 1601 556
rect 1586 516 1589 536
rect 1578 513 1589 516
rect 1482 483 1501 486
rect 1450 433 1461 436
rect 1498 436 1501 483
rect 1578 456 1581 513
rect 1598 486 1601 553
rect 1610 523 1613 573
rect 1682 543 1685 606
rect 1690 603 1701 606
rect 1706 596 1709 716
rect 1698 593 1709 596
rect 1634 513 1637 536
rect 1674 513 1677 536
rect 1682 503 1685 526
rect 1690 523 1693 536
rect 1698 506 1701 593
rect 1694 503 1701 506
rect 1594 483 1601 486
rect 1594 463 1597 483
rect 1578 453 1589 456
rect 1498 433 1509 436
rect 1418 323 1429 326
rect 1418 276 1421 323
rect 1418 273 1429 276
rect 1426 253 1429 273
rect 1266 153 1277 156
rect 1250 143 1269 146
rect 1250 123 1253 143
rect 1258 103 1261 136
rect 1266 133 1269 143
rect 1266 113 1269 126
rect 1274 103 1277 153
rect 1378 133 1381 176
rect 1290 113 1293 126
rect 1298 103 1301 126
rect 1330 113 1333 126
rect 1410 123 1413 206
rect 1418 196 1421 216
rect 1426 203 1429 216
rect 1434 213 1437 316
rect 1450 313 1453 433
rect 1474 396 1477 416
rect 1482 403 1485 416
rect 1490 413 1493 426
rect 1490 396 1493 406
rect 1474 393 1493 396
rect 1506 386 1509 433
rect 1530 413 1533 426
rect 1538 413 1549 416
rect 1570 413 1573 426
rect 1498 383 1509 386
rect 1474 313 1477 326
rect 1498 276 1501 383
rect 1514 333 1525 336
rect 1514 313 1517 326
rect 1522 296 1525 333
rect 1490 273 1501 276
rect 1506 293 1525 296
rect 1434 196 1437 206
rect 1418 193 1437 196
rect 1458 123 1461 216
rect 1466 213 1469 226
rect 1490 206 1493 273
rect 1506 213 1509 293
rect 1466 193 1469 206
rect 1490 203 1501 206
rect 1498 186 1501 203
rect 1514 186 1517 226
rect 1522 213 1525 236
rect 1570 213 1573 316
rect 1490 183 1501 186
rect 1510 183 1517 186
rect 1490 133 1493 183
rect 1510 116 1513 183
rect 1522 123 1525 206
rect 1562 193 1565 206
rect 1578 203 1581 286
rect 1586 213 1589 453
rect 1694 436 1697 503
rect 1694 433 1701 436
rect 1618 363 1621 406
rect 1610 296 1613 336
rect 1642 323 1645 416
rect 1682 403 1685 426
rect 1698 413 1701 433
rect 1690 323 1693 406
rect 1706 403 1709 476
rect 1714 413 1717 626
rect 1722 563 1725 646
rect 1730 593 1733 606
rect 1746 603 1749 733
rect 1754 713 1757 833
rect 1786 813 1789 826
rect 1794 813 1805 816
rect 1810 736 1813 883
rect 1842 843 1845 913
rect 1882 836 1885 1083
rect 1890 1013 1893 1026
rect 1914 993 1917 1093
rect 1946 1023 1949 1126
rect 1954 1123 1957 1136
rect 1962 1133 1965 1143
rect 1930 1003 1933 1016
rect 1962 963 1965 1126
rect 1970 1093 1973 1136
rect 1978 1123 1981 1146
rect 1986 1133 1989 1176
rect 1994 1036 1997 1326
rect 2002 1323 2005 1336
rect 2010 1323 2013 1343
rect 2018 1306 2021 1406
rect 2030 1346 2033 1433
rect 2042 1366 2045 1516
rect 2082 1476 2085 1526
rect 2074 1473 2085 1476
rect 2074 1376 2077 1473
rect 2094 1456 2097 1533
rect 2122 1486 2125 1546
rect 2138 1523 2141 1536
rect 2146 1496 2149 1596
rect 2162 1593 2169 1596
rect 2154 1533 2157 1586
rect 2166 1526 2169 1593
rect 2090 1453 2097 1456
rect 2114 1483 2125 1486
rect 2138 1493 2149 1496
rect 2090 1423 2093 1453
rect 2074 1373 2085 1376
rect 2042 1363 2053 1366
rect 2030 1343 2037 1346
rect 2010 1303 2021 1306
rect 2010 1206 2013 1303
rect 2026 1213 2029 1326
rect 2034 1323 2037 1343
rect 2050 1206 2053 1363
rect 2082 1336 2085 1373
rect 2090 1346 2093 1416
rect 2114 1376 2117 1483
rect 2138 1396 2141 1493
rect 2154 1476 2157 1526
rect 2150 1473 2157 1476
rect 2162 1523 2169 1526
rect 2150 1416 2153 1473
rect 2162 1423 2165 1523
rect 2150 1413 2157 1416
rect 2138 1393 2149 1396
rect 2114 1373 2133 1376
rect 2090 1343 2101 1346
rect 2082 1333 2093 1336
rect 2010 1203 2021 1206
rect 1986 1033 1997 1036
rect 1898 896 1901 926
rect 1962 906 1965 926
rect 1954 903 1965 906
rect 1898 893 1909 896
rect 1906 836 1909 893
rect 1874 833 1885 836
rect 1898 833 1909 836
rect 1826 813 1829 826
rect 1802 733 1813 736
rect 1842 733 1845 756
rect 1874 753 1877 833
rect 1898 803 1901 833
rect 1906 786 1909 816
rect 1922 796 1925 816
rect 1930 803 1933 816
rect 1938 813 1941 846
rect 1954 836 1957 903
rect 1970 896 1973 1016
rect 1986 1013 1989 1033
rect 2002 1013 2005 1126
rect 2018 1096 2021 1203
rect 2042 1203 2053 1206
rect 2042 1133 2045 1203
rect 2050 1133 2053 1146
rect 2010 1093 2021 1096
rect 1994 933 1997 996
rect 2010 976 2013 1093
rect 2018 996 2021 1056
rect 2026 1043 2029 1126
rect 2058 1113 2061 1126
rect 2066 1123 2069 1176
rect 2082 1166 2085 1326
rect 2078 1163 2085 1166
rect 2090 1163 2093 1333
rect 2098 1326 2101 1343
rect 2098 1323 2105 1326
rect 2102 1236 2105 1323
rect 2098 1233 2105 1236
rect 2078 1086 2081 1163
rect 2098 1133 2101 1233
rect 2106 1186 2109 1216
rect 2106 1183 2113 1186
rect 2098 1113 2101 1126
rect 2110 1106 2113 1183
rect 2130 1146 2133 1373
rect 2146 1313 2149 1393
rect 2154 1306 2157 1413
rect 2146 1303 2157 1306
rect 2146 1236 2149 1303
rect 2146 1233 2153 1236
rect 2150 1166 2153 1233
rect 2106 1103 2113 1106
rect 2122 1143 2133 1146
rect 2146 1163 2153 1166
rect 2034 1013 2037 1086
rect 2078 1083 2085 1086
rect 2058 1036 2061 1056
rect 2050 1033 2061 1036
rect 2018 993 2029 996
rect 2010 973 2021 976
rect 2010 923 2013 966
rect 1970 893 1981 896
rect 1954 833 1965 836
rect 1938 796 1941 806
rect 1922 793 1941 796
rect 1906 783 1917 786
rect 1754 613 1757 626
rect 1762 593 1765 726
rect 1770 616 1773 716
rect 1802 656 1805 733
rect 1818 656 1821 726
rect 1802 653 1813 656
rect 1818 653 1829 656
rect 1770 613 1781 616
rect 1770 483 1773 606
rect 1778 416 1781 613
rect 1786 613 1797 616
rect 1786 533 1789 613
rect 1802 586 1805 616
rect 1798 583 1805 586
rect 1798 496 1801 583
rect 1810 523 1813 653
rect 1818 603 1821 626
rect 1826 613 1829 653
rect 1858 613 1861 746
rect 1882 713 1885 736
rect 1890 656 1893 756
rect 1898 733 1901 746
rect 1890 653 1897 656
rect 1894 576 1897 653
rect 1906 613 1909 726
rect 1914 683 1917 783
rect 1938 713 1941 726
rect 1946 636 1949 816
rect 1954 736 1957 816
rect 1962 813 1965 833
rect 1970 786 1973 876
rect 1978 803 1981 893
rect 2010 813 2013 826
rect 2018 803 2021 973
rect 2026 883 2029 993
rect 2050 986 2053 1033
rect 2050 983 2061 986
rect 2050 946 2053 966
rect 2046 943 2053 946
rect 2046 836 2049 943
rect 2026 813 2029 836
rect 2046 833 2053 836
rect 2034 803 2037 826
rect 1970 783 1989 786
rect 1954 733 1965 736
rect 1954 693 1957 726
rect 1962 713 1965 733
rect 1946 633 1957 636
rect 1890 573 1897 576
rect 1794 493 1801 496
rect 1722 383 1725 406
rect 1730 393 1733 406
rect 1594 293 1613 296
rect 1594 176 1597 293
rect 1730 276 1733 336
rect 1746 333 1749 356
rect 1738 313 1741 326
rect 1754 323 1757 336
rect 1762 306 1765 416
rect 1770 413 1781 416
rect 1786 413 1789 426
rect 1794 403 1797 493
rect 1802 413 1805 466
rect 1810 413 1813 486
rect 1842 413 1845 526
rect 1850 513 1853 526
rect 1802 346 1805 406
rect 1802 343 1813 346
rect 1754 303 1765 306
rect 1730 273 1741 276
rect 1602 213 1605 226
rect 1602 183 1605 206
rect 1610 203 1613 216
rect 1594 173 1605 176
rect 1602 133 1605 173
rect 1618 133 1621 216
rect 1626 193 1629 206
rect 1666 203 1669 216
rect 1674 203 1677 226
rect 1690 203 1693 216
rect 1674 133 1677 146
rect 1510 113 1517 116
rect 1578 113 1581 126
rect 1618 113 1621 126
rect 1698 123 1701 216
rect 1706 193 1709 216
rect 1730 213 1733 226
rect 1738 203 1741 273
rect 1754 236 1757 303
rect 1754 233 1765 236
rect 1746 203 1749 216
rect 1762 213 1765 233
rect 1770 223 1773 336
rect 1754 123 1757 206
rect 1778 123 1781 336
rect 1786 313 1789 326
rect 1794 303 1797 336
rect 1802 323 1805 336
rect 1786 196 1789 216
rect 1794 203 1797 216
rect 1802 213 1805 256
rect 1810 213 1813 343
rect 1842 333 1845 346
rect 1826 306 1829 326
rect 1826 303 1837 306
rect 1834 236 1837 303
rect 1826 233 1837 236
rect 1802 196 1805 206
rect 1786 193 1805 196
rect 1826 183 1829 233
rect 1842 123 1845 216
rect 1858 203 1861 216
rect 1874 213 1877 256
rect 1890 226 1893 573
rect 1938 556 1941 606
rect 1954 573 1957 633
rect 1930 553 1949 556
rect 1906 513 1909 526
rect 1906 403 1909 506
rect 1906 313 1909 326
rect 1882 223 1893 226
rect 1882 166 1885 223
rect 1874 163 1885 166
rect 1874 133 1877 163
rect 1898 123 1901 226
rect 1906 163 1909 236
rect 1930 233 1933 553
rect 1946 513 1949 526
rect 1938 413 1941 436
rect 1954 413 1957 536
rect 1962 526 1965 686
rect 1986 666 1989 783
rect 2042 746 2045 816
rect 1970 663 1989 666
rect 2026 743 2045 746
rect 1970 613 1973 663
rect 2026 613 2029 743
rect 2050 613 2053 833
rect 2058 713 2061 983
rect 2082 963 2085 1083
rect 2106 1043 2109 1103
rect 2098 953 2101 1016
rect 2122 1003 2125 1143
rect 2146 1053 2149 1163
rect 2162 1063 2165 1416
rect 2170 1103 2173 1506
rect 2178 1473 2181 1833
rect 2186 1813 2205 1816
rect 2234 1806 2237 1983
rect 2242 1933 2245 2066
rect 2250 2013 2253 2136
rect 2266 2076 2269 2153
rect 2282 2133 2285 2186
rect 2290 2163 2293 2206
rect 2306 2123 2309 2216
rect 2314 2196 2317 2233
rect 2322 2213 2325 2416
rect 2330 2403 2333 2426
rect 2338 2393 2341 2536
rect 2346 2493 2349 2553
rect 2354 2523 2357 2686
rect 2362 2533 2365 2726
rect 2370 2686 2373 2736
rect 2378 2706 2381 2766
rect 2394 2746 2397 2863
rect 2414 2846 2417 2933
rect 2410 2843 2417 2846
rect 2402 2803 2405 2816
rect 2386 2743 2397 2746
rect 2386 2733 2389 2743
rect 2394 2723 2397 2736
rect 2402 2723 2405 2746
rect 2378 2703 2389 2706
rect 2370 2683 2377 2686
rect 2374 2566 2377 2683
rect 2370 2563 2377 2566
rect 2370 2476 2373 2563
rect 2386 2546 2389 2703
rect 2362 2473 2373 2476
rect 2378 2543 2389 2546
rect 2362 2356 2365 2473
rect 2378 2456 2381 2543
rect 2386 2506 2389 2526
rect 2386 2503 2397 2506
rect 2394 2456 2397 2503
rect 2410 2473 2413 2843
rect 2418 2803 2421 2826
rect 2426 2763 2429 2943
rect 2450 2936 2453 3303
rect 2458 3153 2461 3286
rect 2474 3266 2477 3503
rect 2490 3376 2493 3626
rect 2514 3603 2517 3616
rect 2530 3613 2533 3626
rect 2530 3603 2541 3606
rect 2486 3373 2493 3376
rect 2486 3286 2489 3373
rect 2498 3296 2501 3586
rect 2506 3503 2509 3556
rect 2522 3523 2525 3536
rect 2514 3496 2517 3516
rect 2546 3513 2549 3643
rect 2558 3626 2561 3713
rect 2578 3703 2581 3736
rect 2558 3623 2565 3626
rect 2570 3623 2573 3686
rect 2586 3623 2589 3823
rect 2610 3813 2613 3826
rect 2626 3793 2629 3883
rect 2650 3813 2653 3826
rect 2698 3813 2709 3816
rect 2594 3713 2597 3736
rect 2602 3723 2605 3736
rect 2642 3713 2645 3726
rect 2514 3493 2525 3496
rect 2522 3436 2525 3493
rect 2514 3433 2525 3436
rect 2506 3413 2509 3426
rect 2514 3413 2517 3433
rect 2554 3423 2557 3606
rect 2562 3533 2565 3623
rect 2586 3603 2589 3616
rect 2570 3523 2573 3546
rect 2586 3426 2589 3586
rect 2602 3533 2605 3546
rect 2562 3423 2573 3426
rect 2582 3423 2589 3426
rect 2610 3423 2613 3616
rect 2618 3583 2621 3626
rect 2658 3613 2661 3796
rect 2706 3793 2709 3813
rect 2714 3803 2717 3916
rect 2730 3843 2733 3986
rect 2754 3983 2757 4113
rect 2826 4036 2829 4163
rect 2846 4116 2849 4163
rect 2866 4156 2869 4206
rect 2874 4203 2877 4216
rect 2858 4153 2869 4156
rect 2858 4123 2861 4153
rect 2846 4113 2853 4116
rect 2826 4033 2837 4036
rect 2762 3923 2765 4016
rect 2778 3906 2781 3966
rect 2810 3923 2813 4016
rect 2818 3996 2821 4016
rect 2818 3993 2825 3996
rect 2822 3916 2825 3993
rect 2770 3903 2781 3906
rect 2818 3913 2825 3916
rect 2770 3836 2773 3903
rect 2770 3833 2781 3836
rect 2754 3783 2757 3816
rect 2778 3793 2781 3833
rect 2786 3813 2789 3826
rect 2794 3803 2797 3896
rect 2802 3803 2805 3836
rect 2810 3793 2813 3806
rect 2746 3743 2749 3766
rect 2682 3713 2685 3726
rect 2738 3703 2741 3726
rect 2786 3716 2789 3786
rect 2802 3723 2813 3726
rect 2786 3713 2793 3716
rect 2666 3533 2669 3616
rect 2682 3613 2701 3616
rect 2618 3486 2621 3526
rect 2634 3513 2637 3526
rect 2642 3503 2645 3526
rect 2674 3503 2677 3546
rect 2690 3523 2693 3546
rect 2618 3483 2629 3486
rect 2506 3393 2509 3406
rect 2498 3293 2505 3296
rect 2486 3283 2493 3286
rect 2474 3263 2485 3266
rect 2474 3213 2477 3246
rect 2482 3223 2485 3263
rect 2466 3203 2477 3206
rect 2482 3203 2485 3216
rect 2490 3213 2493 3283
rect 2502 3216 2505 3293
rect 2498 3213 2505 3216
rect 2498 3193 2501 3213
rect 2458 3113 2461 3136
rect 2474 3093 2477 3136
rect 2498 3093 2501 3126
rect 2514 3066 2517 3406
rect 2530 3333 2533 3416
rect 2562 3413 2565 3423
rect 2546 3313 2549 3326
rect 2530 3203 2533 3246
rect 2554 3243 2557 3406
rect 2570 3353 2573 3406
rect 2582 3376 2585 3423
rect 2626 3416 2629 3483
rect 2582 3373 2589 3376
rect 2562 3286 2565 3306
rect 2562 3283 2569 3286
rect 2566 3216 2569 3283
rect 2562 3213 2569 3216
rect 2554 3186 2557 3196
rect 2562 3193 2565 3213
rect 2578 3193 2581 3226
rect 2554 3183 2561 3186
rect 2538 3133 2549 3136
rect 2522 3113 2525 3126
rect 2538 3106 2541 3126
rect 2506 3063 2517 3066
rect 2534 3103 2541 3106
rect 2450 2933 2461 2936
rect 2418 2733 2421 2756
rect 2434 2746 2437 2826
rect 2442 2813 2445 2926
rect 2458 2836 2461 2933
rect 2450 2833 2461 2836
rect 2430 2743 2437 2746
rect 2418 2713 2421 2726
rect 2430 2636 2433 2743
rect 2442 2733 2445 2746
rect 2430 2633 2437 2636
rect 2418 2593 2421 2616
rect 2426 2583 2429 2606
rect 2434 2576 2437 2633
rect 2442 2603 2445 2726
rect 2426 2573 2437 2576
rect 2374 2453 2381 2456
rect 2386 2453 2397 2456
rect 2374 2376 2377 2453
rect 2374 2373 2381 2376
rect 2362 2353 2369 2356
rect 2330 2283 2333 2346
rect 2346 2316 2349 2336
rect 2342 2313 2349 2316
rect 2342 2256 2345 2313
rect 2342 2253 2349 2256
rect 2346 2236 2349 2253
rect 2354 2243 2357 2326
rect 2346 2233 2357 2236
rect 2346 2213 2349 2226
rect 2354 2196 2357 2233
rect 2366 2226 2369 2353
rect 2366 2223 2373 2226
rect 2314 2193 2325 2196
rect 2322 2116 2325 2193
rect 2350 2193 2357 2196
rect 2362 2193 2365 2206
rect 2350 2136 2353 2193
rect 2350 2133 2357 2136
rect 2314 2113 2325 2116
rect 2354 2116 2357 2133
rect 2362 2123 2365 2166
rect 2354 2113 2365 2116
rect 2266 2073 2277 2076
rect 2274 2006 2277 2073
rect 2258 2003 2277 2006
rect 2258 1856 2261 2003
rect 2266 1923 2269 1956
rect 2258 1853 2269 1856
rect 2194 1733 2197 1806
rect 2226 1803 2237 1806
rect 2202 1726 2205 1746
rect 2186 1723 2205 1726
rect 2186 1706 2189 1723
rect 2186 1703 2197 1706
rect 2194 1646 2197 1703
rect 2226 1666 2229 1803
rect 2242 1743 2245 1806
rect 2258 1803 2261 1846
rect 2242 1726 2245 1736
rect 2250 1733 2253 1746
rect 2258 1733 2261 1776
rect 2266 1756 2269 1853
rect 2274 1803 2277 1816
rect 2282 1783 2285 1806
rect 2290 1803 2293 1866
rect 2298 1793 2301 1806
rect 2266 1753 2277 1756
rect 2266 1733 2269 1746
rect 2242 1723 2261 1726
rect 2226 1663 2237 1666
rect 2190 1643 2197 1646
rect 2190 1536 2193 1643
rect 2210 1543 2213 1606
rect 2186 1533 2193 1536
rect 2178 1333 2181 1406
rect 2186 1343 2189 1533
rect 2194 1376 2197 1516
rect 2202 1403 2205 1526
rect 2234 1513 2237 1663
rect 2242 1596 2245 1723
rect 2250 1613 2253 1696
rect 2274 1656 2277 1753
rect 2282 1686 2285 1746
rect 2290 1723 2293 1736
rect 2314 1726 2317 2113
rect 2362 2096 2365 2113
rect 2354 2093 2365 2096
rect 2354 2036 2357 2093
rect 2354 2033 2365 2036
rect 2330 2013 2333 2026
rect 2354 1933 2357 2016
rect 2362 1993 2365 2033
rect 2370 1963 2373 2223
rect 2378 1983 2381 2373
rect 2386 2323 2389 2453
rect 2394 2353 2397 2436
rect 2402 2413 2405 2426
rect 2418 2416 2421 2526
rect 2426 2483 2429 2573
rect 2434 2533 2437 2566
rect 2410 2413 2421 2416
rect 2426 2406 2429 2476
rect 2442 2443 2445 2596
rect 2442 2413 2445 2426
rect 2402 2333 2405 2406
rect 2410 2403 2429 2406
rect 2394 2256 2397 2326
rect 2394 2253 2401 2256
rect 2386 2203 2389 2246
rect 2398 2196 2401 2253
rect 2394 2193 2401 2196
rect 2386 2113 2389 2126
rect 2394 2106 2397 2193
rect 2410 2123 2413 2403
rect 2450 2366 2453 2833
rect 2466 2776 2469 2816
rect 2474 2803 2477 2936
rect 2490 2923 2493 3016
rect 2498 2873 2501 3016
rect 2506 2953 2509 3063
rect 2514 2996 2517 3016
rect 2522 3003 2525 3056
rect 2534 3036 2537 3103
rect 2534 3033 2541 3036
rect 2546 3033 2549 3133
rect 2558 3086 2561 3183
rect 2586 3136 2589 3373
rect 2594 3363 2597 3416
rect 2618 3413 2629 3416
rect 2618 3353 2621 3413
rect 2594 3313 2597 3326
rect 2594 3213 2613 3216
rect 2594 3203 2597 3213
rect 2634 3196 2637 3336
rect 2650 3296 2653 3336
rect 2646 3293 2653 3296
rect 2646 3236 2649 3293
rect 2646 3233 2653 3236
rect 2642 3203 2645 3216
rect 2650 3213 2653 3233
rect 2626 3193 2637 3196
rect 2586 3133 2597 3136
rect 2578 3093 2581 3126
rect 2594 3086 2597 3133
rect 2558 3083 2565 3086
rect 2530 2996 2533 3006
rect 2538 3003 2541 3033
rect 2514 2993 2533 2996
rect 2482 2813 2485 2826
rect 2538 2816 2541 2936
rect 2554 2906 2557 2956
rect 2562 2923 2565 3083
rect 2586 3083 2597 3086
rect 2554 2903 2565 2906
rect 2562 2836 2565 2903
rect 2554 2833 2565 2836
rect 2490 2803 2493 2816
rect 2498 2803 2501 2816
rect 2538 2813 2549 2816
rect 2458 2773 2469 2776
rect 2458 2696 2461 2773
rect 2466 2716 2469 2766
rect 2482 2733 2485 2786
rect 2522 2723 2533 2726
rect 2466 2713 2485 2716
rect 2458 2693 2469 2696
rect 2466 2616 2469 2693
rect 2458 2613 2469 2616
rect 2458 2593 2461 2613
rect 2482 2556 2485 2713
rect 2530 2613 2533 2723
rect 2538 2676 2541 2806
rect 2546 2783 2549 2813
rect 2554 2803 2557 2833
rect 2562 2796 2565 2816
rect 2570 2803 2573 2816
rect 2578 2796 2581 2806
rect 2562 2793 2581 2796
rect 2578 2766 2581 2786
rect 2574 2763 2581 2766
rect 2546 2743 2565 2746
rect 2546 2723 2549 2743
rect 2554 2703 2557 2736
rect 2562 2733 2565 2743
rect 2574 2706 2577 2763
rect 2586 2713 2589 3083
rect 2602 3013 2605 3026
rect 2610 2953 2613 3056
rect 2594 2943 2613 2946
rect 2594 2923 2597 2943
rect 2602 2923 2605 2936
rect 2610 2933 2613 2943
rect 2618 2866 2621 3006
rect 2610 2863 2621 2866
rect 2574 2703 2581 2706
rect 2538 2673 2549 2676
rect 2466 2553 2485 2556
rect 2466 2536 2469 2553
rect 2458 2403 2461 2536
rect 2466 2533 2477 2536
rect 2474 2466 2477 2533
rect 2466 2463 2477 2466
rect 2442 2363 2453 2366
rect 2418 2336 2421 2356
rect 2418 2333 2429 2336
rect 2426 2206 2429 2333
rect 2442 2286 2445 2363
rect 2442 2283 2453 2286
rect 2450 2206 2453 2283
rect 2466 2276 2469 2463
rect 2490 2403 2493 2536
rect 2506 2413 2509 2466
rect 2490 2346 2493 2396
rect 2486 2343 2493 2346
rect 2462 2273 2469 2276
rect 2462 2216 2465 2273
rect 2462 2213 2469 2216
rect 2474 2213 2477 2326
rect 2486 2296 2489 2343
rect 2486 2293 2493 2296
rect 2490 2213 2493 2293
rect 2418 2203 2429 2206
rect 2442 2203 2453 2206
rect 2418 2183 2421 2203
rect 2442 2156 2445 2203
rect 2466 2196 2469 2213
rect 2442 2153 2453 2156
rect 2426 2133 2445 2136
rect 2426 2106 2429 2133
rect 2394 2103 2405 2106
rect 2402 2046 2405 2103
rect 2394 2043 2405 2046
rect 2418 2103 2429 2106
rect 2394 2023 2397 2043
rect 2418 1956 2421 2103
rect 2418 1953 2425 1956
rect 2378 1933 2397 1936
rect 2386 1913 2389 1926
rect 2346 1743 2349 1806
rect 2314 1723 2325 1726
rect 2354 1723 2357 1816
rect 2378 1813 2381 1836
rect 2378 1763 2381 1806
rect 2362 1726 2365 1736
rect 2370 1733 2373 1746
rect 2362 1723 2381 1726
rect 2394 1723 2397 1933
rect 2410 1886 2413 1936
rect 2422 1896 2425 1953
rect 2434 1906 2437 2126
rect 2450 1946 2453 2153
rect 2458 2123 2461 2196
rect 2466 2193 2477 2196
rect 2474 2136 2477 2193
rect 2514 2186 2517 2356
rect 2530 2343 2533 2526
rect 2546 2403 2549 2673
rect 2578 2573 2581 2703
rect 2594 2613 2597 2816
rect 2610 2813 2613 2863
rect 2626 2796 2629 3193
rect 2658 3133 2661 3406
rect 2674 3353 2677 3416
rect 2666 3306 2669 3326
rect 2666 3303 2677 3306
rect 2674 3246 2677 3303
rect 2666 3243 2677 3246
rect 2666 3213 2669 3243
rect 2674 3203 2677 3226
rect 2682 3196 2685 3206
rect 2674 3193 2685 3196
rect 2642 3113 2645 3126
rect 2674 3123 2677 3193
rect 2642 3013 2645 3026
rect 2690 3013 2693 3426
rect 2698 3413 2701 3613
rect 2706 3533 2709 3546
rect 2706 3513 2709 3526
rect 2738 3523 2741 3616
rect 2762 3603 2765 3616
rect 2778 3603 2781 3706
rect 2790 3666 2793 3713
rect 2786 3663 2793 3666
rect 2754 3533 2757 3556
rect 2786 3523 2789 3663
rect 2802 3606 2805 3723
rect 2802 3603 2813 3606
rect 2818 3586 2821 3913
rect 2826 3813 2829 3856
rect 2826 3733 2829 3746
rect 2834 3716 2837 4033
rect 2842 4003 2845 4026
rect 2850 3936 2853 4113
rect 2866 4063 2869 4136
rect 2882 4016 2885 4216
rect 2890 4193 2893 4226
rect 2906 4213 2909 4326
rect 2938 4313 2941 4326
rect 2930 4193 2933 4306
rect 2954 4293 2957 4336
rect 2962 4323 2965 4406
rect 2994 4403 2997 4456
rect 3010 4453 3021 4456
rect 3002 4403 3005 4436
rect 3010 4386 3013 4453
rect 3002 4383 3013 4386
rect 3002 4336 3005 4383
rect 2970 4323 2973 4336
rect 3002 4333 3013 4336
rect 2946 4213 2949 4226
rect 2954 4213 2973 4216
rect 2954 4203 2957 4213
rect 2970 4153 2973 4206
rect 2978 4203 2981 4216
rect 2986 4196 2989 4226
rect 3010 4223 3013 4333
rect 3026 4323 3029 4426
rect 3058 4383 3061 4406
rect 3066 4333 3069 4416
rect 3074 4413 3077 4436
rect 3090 4413 3093 4473
rect 3082 4393 3085 4406
rect 3098 4403 3101 4503
rect 3106 4433 3109 4526
rect 2978 4193 2989 4196
rect 2890 4106 2893 4126
rect 2898 4123 2901 4136
rect 2906 4116 2909 4136
rect 2906 4113 2917 4116
rect 2890 4103 2897 4106
rect 2894 4026 2897 4103
rect 2914 4046 2917 4113
rect 2866 4013 2885 4016
rect 2890 4023 2897 4026
rect 2906 4043 2917 4046
rect 2906 4023 2909 4043
rect 2890 4003 2893 4023
rect 2850 3933 2861 3936
rect 2850 3856 2853 3926
rect 2858 3916 2861 3933
rect 2858 3913 2865 3916
rect 2842 3853 2853 3856
rect 2842 3743 2845 3853
rect 2862 3836 2865 3913
rect 2874 3853 2877 3936
rect 2882 3933 2885 3946
rect 2898 3913 2901 4006
rect 2922 3893 2925 3926
rect 2858 3833 2865 3836
rect 2858 3816 2861 3833
rect 2850 3813 2861 3816
rect 2830 3713 2837 3716
rect 2842 3713 2845 3736
rect 2830 3646 2833 3713
rect 2850 3706 2853 3813
rect 2858 3723 2861 3806
rect 2850 3703 2857 3706
rect 2830 3643 2837 3646
rect 2826 3613 2829 3626
rect 2826 3593 2829 3606
rect 2810 3583 2821 3586
rect 2706 3413 2709 3506
rect 2810 3446 2813 3583
rect 2834 3566 2837 3643
rect 2826 3563 2837 3566
rect 2826 3466 2829 3563
rect 2842 3546 2845 3696
rect 2854 3636 2857 3703
rect 2866 3693 2869 3746
rect 2874 3703 2877 3736
rect 2838 3543 2845 3546
rect 2850 3633 2857 3636
rect 2838 3486 2841 3543
rect 2850 3496 2853 3633
rect 2858 3533 2861 3616
rect 2866 3593 2869 3626
rect 2866 3513 2869 3526
rect 2874 3506 2877 3536
rect 2882 3516 2885 3826
rect 2906 3736 2909 3816
rect 2914 3803 2917 3826
rect 2922 3803 2925 3816
rect 2930 3796 2933 3906
rect 2938 3823 2941 4116
rect 2970 4103 2973 4116
rect 2978 4113 2981 4193
rect 2986 4113 2989 4136
rect 2994 4133 2997 4196
rect 3010 4126 3013 4176
rect 3034 4133 3037 4146
rect 2994 4123 3013 4126
rect 2930 3793 2941 3796
rect 2930 3766 2933 3786
rect 2890 3733 2909 3736
rect 2922 3763 2933 3766
rect 2890 3563 2893 3606
rect 2906 3603 2909 3726
rect 2922 3636 2925 3763
rect 2938 3746 2941 3793
rect 2946 3773 2949 3936
rect 2934 3743 2941 3746
rect 2934 3676 2937 3743
rect 2946 3683 2949 3736
rect 2954 3713 2957 3826
rect 2934 3673 2941 3676
rect 2922 3633 2933 3636
rect 2914 3603 2917 3616
rect 2930 3613 2933 3633
rect 2938 3596 2941 3673
rect 2930 3593 2941 3596
rect 2906 3533 2909 3556
rect 2914 3523 2917 3536
rect 2882 3513 2917 3516
rect 2874 3503 2885 3506
rect 2850 3493 2861 3496
rect 2838 3483 2845 3486
rect 2826 3463 2837 3466
rect 2810 3443 2821 3446
rect 2730 3413 2733 3426
rect 2706 3363 2709 3406
rect 2746 3383 2749 3396
rect 2786 3383 2789 3406
rect 2706 3333 2709 3356
rect 2738 3236 2741 3326
rect 2746 3303 2749 3326
rect 2754 3313 2757 3326
rect 2770 3323 2773 3336
rect 2794 3333 2797 3406
rect 2802 3403 2805 3416
rect 2810 3366 2813 3426
rect 2802 3363 2813 3366
rect 2794 3313 2797 3326
rect 2738 3233 2749 3236
rect 2730 3166 2733 3216
rect 2730 3163 2741 3166
rect 2698 3123 2701 3136
rect 2714 3046 2717 3156
rect 2738 3123 2741 3163
rect 2746 3153 2749 3233
rect 2770 3213 2773 3306
rect 2802 3256 2805 3363
rect 2786 3253 2805 3256
rect 2786 3176 2789 3253
rect 2810 3223 2813 3356
rect 2786 3173 2797 3176
rect 2794 3136 2797 3173
rect 2794 3133 2805 3136
rect 2786 3123 2797 3126
rect 2802 3106 2805 3133
rect 2810 3123 2813 3186
rect 2794 3103 2805 3106
rect 2714 3043 2725 3046
rect 2690 2986 2693 3006
rect 2706 3003 2709 3036
rect 2722 2986 2725 3043
rect 2794 3036 2797 3103
rect 2818 3036 2821 3443
rect 2826 3383 2829 3416
rect 2834 3303 2837 3463
rect 2842 3423 2845 3483
rect 2842 3383 2845 3416
rect 2858 3376 2861 3493
rect 2882 3423 2885 3503
rect 2930 3496 2933 3593
rect 2922 3493 2933 3496
rect 2946 3526 2949 3616
rect 2962 3613 2965 3966
rect 2986 3856 2989 4016
rect 2994 3996 2997 4056
rect 3002 4013 3005 4123
rect 3050 4053 3053 4216
rect 3066 4173 3069 4326
rect 3074 4313 3077 4336
rect 3090 4333 3093 4346
rect 3090 4136 3093 4326
rect 3106 4203 3109 4226
rect 3114 4196 3117 4406
rect 3138 4343 3141 4606
rect 3162 4596 3165 4676
rect 3154 4593 3165 4596
rect 3154 4513 3157 4593
rect 3162 4523 3165 4536
rect 3170 4533 3173 4616
rect 3178 4523 3181 4546
rect 3242 4543 3245 4616
rect 3186 4523 3189 4536
rect 3162 4393 3165 4416
rect 3122 4213 3125 4316
rect 3130 4306 3133 4326
rect 3186 4313 3189 4326
rect 3194 4306 3197 4326
rect 3210 4323 3213 4536
rect 3250 4516 3253 4536
rect 3266 4533 3269 4606
rect 3282 4593 3285 4606
rect 3306 4603 3309 4616
rect 3282 4536 3285 4576
rect 3362 4543 3365 4616
rect 3242 4513 3253 4516
rect 3242 4436 3245 4513
rect 3258 4453 3261 4526
rect 3274 4523 3277 4536
rect 3282 4533 3293 4536
rect 3282 4513 3285 4526
rect 3354 4456 3357 4536
rect 3370 4533 3373 4616
rect 3434 4603 3437 4616
rect 3458 4593 3461 4606
rect 3482 4593 3485 4636
rect 3354 4453 3365 4456
rect 3242 4433 3253 4436
rect 3130 4303 3137 4306
rect 3134 4226 3137 4303
rect 3130 4223 3137 4226
rect 3186 4303 3197 4306
rect 3130 4203 3133 4223
rect 3058 4103 3061 4126
rect 3066 4013 3069 4136
rect 3082 4133 3093 4136
rect 3106 4193 3117 4196
rect 3074 4113 3077 4126
rect 2994 3993 3001 3996
rect 2998 3926 3001 3993
rect 3026 3983 3029 4006
rect 3042 3963 3045 4006
rect 3082 3986 3085 4133
rect 3090 4113 3093 4126
rect 3078 3983 3085 3986
rect 2994 3923 3001 3926
rect 3010 3923 3013 3946
rect 2994 3903 2997 3923
rect 3066 3896 3069 3926
rect 3058 3893 3069 3896
rect 2982 3853 2989 3856
rect 2970 3783 2973 3816
rect 2982 3746 2985 3853
rect 2982 3743 2989 3746
rect 2986 3726 2989 3743
rect 2994 3733 2997 3846
rect 3002 3803 3005 3816
rect 3010 3786 3013 3856
rect 3058 3846 3061 3893
rect 3058 3843 3069 3846
rect 3006 3783 3013 3786
rect 2970 3723 2989 3726
rect 3006 3716 3009 3783
rect 3018 3723 3021 3826
rect 3042 3813 3045 3826
rect 3066 3813 3069 3843
rect 3026 3793 3029 3806
rect 3034 3803 3045 3806
rect 3050 3733 3053 3806
rect 3078 3766 3081 3983
rect 3090 3766 3093 3976
rect 3106 3853 3109 4193
rect 3114 3996 3117 4186
rect 3146 4183 3149 4206
rect 3122 4116 3125 4136
rect 3154 4133 3157 4206
rect 3170 4123 3173 4146
rect 3122 4113 3133 4116
rect 3178 4113 3181 4136
rect 3130 4036 3133 4113
rect 3122 4033 3133 4036
rect 3122 4013 3125 4033
rect 3114 3993 3121 3996
rect 3106 3793 3109 3816
rect 3118 3786 3121 3993
rect 3130 3973 3133 4006
rect 3138 3933 3141 3946
rect 3162 3926 3165 3996
rect 3130 3913 3133 3926
rect 3154 3923 3165 3926
rect 3130 3796 3133 3826
rect 3130 3793 3141 3796
rect 3114 3783 3121 3786
rect 3078 3763 3085 3766
rect 3090 3763 3101 3766
rect 3082 3746 3085 3763
rect 3082 3743 3089 3746
rect 3006 3713 3013 3716
rect 3010 3646 3013 3713
rect 3010 3643 3029 3646
rect 2978 3603 2981 3626
rect 2994 3576 2997 3616
rect 2994 3573 3013 3576
rect 2946 3523 2965 3526
rect 2850 3373 2861 3376
rect 2842 3313 2845 3366
rect 2850 3296 2853 3373
rect 2858 3333 2861 3356
rect 2858 3313 2861 3326
rect 2846 3293 2853 3296
rect 2826 3213 2829 3226
rect 2834 3193 2837 3206
rect 2846 3186 2849 3293
rect 2866 3276 2869 3326
rect 2858 3273 2869 3276
rect 2846 3183 2853 3186
rect 2858 3183 2861 3273
rect 2826 3163 2845 3166
rect 2826 3143 2829 3163
rect 2834 3113 2837 3156
rect 2842 3143 2845 3163
rect 2842 3113 2845 3136
rect 2794 3033 2805 3036
rect 2794 3003 2797 3016
rect 2690 2983 2725 2986
rect 2690 2966 2693 2983
rect 2682 2963 2693 2966
rect 2666 2913 2669 2926
rect 2682 2906 2685 2963
rect 2770 2933 2773 2946
rect 2706 2913 2709 2926
rect 2754 2923 2765 2926
rect 2618 2793 2629 2796
rect 2618 2746 2621 2793
rect 2618 2743 2629 2746
rect 2626 2723 2629 2743
rect 2594 2593 2597 2606
rect 2602 2596 2605 2646
rect 2602 2593 2613 2596
rect 2610 2576 2613 2593
rect 2602 2573 2613 2576
rect 2554 2543 2573 2546
rect 2554 2523 2557 2543
rect 2562 2493 2565 2536
rect 2570 2533 2573 2543
rect 2570 2413 2573 2426
rect 2586 2416 2589 2526
rect 2602 2516 2605 2573
rect 2618 2523 2621 2616
rect 2626 2613 2629 2716
rect 2634 2666 2637 2906
rect 2658 2903 2685 2906
rect 2642 2813 2645 2826
rect 2658 2733 2661 2903
rect 2682 2813 2685 2826
rect 2730 2813 2741 2816
rect 2778 2803 2781 2876
rect 2786 2803 2789 2816
rect 2746 2783 2749 2796
rect 2802 2763 2805 3033
rect 2814 3033 2821 3036
rect 2814 2986 2817 3033
rect 2826 3013 2829 3026
rect 2834 3003 2837 3026
rect 2850 3003 2853 3183
rect 2866 3143 2869 3266
rect 2874 3226 2877 3416
rect 2882 3383 2885 3406
rect 2890 3403 2893 3476
rect 2898 3436 2901 3456
rect 2898 3433 2909 3436
rect 2882 3246 2885 3336
rect 2890 3333 2893 3366
rect 2906 3346 2909 3433
rect 2922 3356 2925 3493
rect 2946 3453 2949 3523
rect 2970 3513 2973 3536
rect 2970 3443 2973 3486
rect 2978 3473 2981 3536
rect 2946 3366 2949 3426
rect 2986 3403 2989 3526
rect 2994 3523 3005 3526
rect 3010 3516 3013 3573
rect 3026 3566 3029 3643
rect 3066 3623 3069 3726
rect 3042 3593 3045 3616
rect 3074 3613 3077 3736
rect 3086 3656 3089 3743
rect 3082 3653 3089 3656
rect 3082 3613 3085 3653
rect 3098 3636 3101 3763
rect 3090 3633 3101 3636
rect 3082 3586 3085 3606
rect 3018 3563 3029 3566
rect 3074 3583 3085 3586
rect 3018 3523 3021 3563
rect 3026 3533 3029 3546
rect 3034 3543 3053 3546
rect 3034 3526 3037 3543
rect 3050 3536 3053 3543
rect 3050 3533 3061 3536
rect 3034 3523 3045 3526
rect 3010 3513 3021 3516
rect 2994 3413 2997 3476
rect 3002 3373 3005 3486
rect 3018 3366 3021 3513
rect 3042 3413 3045 3523
rect 3050 3503 3053 3526
rect 3066 3513 3069 3526
rect 3074 3523 3077 3583
rect 3082 3573 3085 3583
rect 3082 3513 3085 3526
rect 3066 3366 3069 3386
rect 2946 3363 2957 3366
rect 3018 3363 3029 3366
rect 2922 3353 2941 3356
rect 2898 3343 2909 3346
rect 2890 3313 2893 3326
rect 2898 3256 2901 3343
rect 2938 3336 2941 3353
rect 2906 3303 2909 3326
rect 2930 3323 2933 3336
rect 2938 3333 2945 3336
rect 2922 3303 2925 3316
rect 2898 3253 2905 3256
rect 2882 3243 2893 3246
rect 2874 3223 2881 3226
rect 2878 3166 2881 3223
rect 2874 3163 2881 3166
rect 2858 3123 2861 3136
rect 2866 3113 2869 3126
rect 2858 3013 2861 3026
rect 2874 3016 2877 3163
rect 2882 3133 2885 3146
rect 2890 3123 2893 3243
rect 2902 3156 2905 3253
rect 2914 3203 2917 3256
rect 2930 3213 2933 3316
rect 2942 3206 2945 3333
rect 2922 3193 2925 3206
rect 2938 3203 2945 3206
rect 2898 3153 2905 3156
rect 2874 3013 2881 3016
rect 2814 2983 2821 2986
rect 2818 2966 2821 2983
rect 2826 2973 2829 2996
rect 2818 2963 2829 2966
rect 2826 2946 2829 2963
rect 2850 2956 2853 2996
rect 2858 2983 2861 2996
rect 2818 2943 2829 2946
rect 2818 2846 2821 2943
rect 2834 2853 2837 2936
rect 2842 2933 2845 2956
rect 2850 2953 2861 2956
rect 2818 2843 2829 2846
rect 2810 2803 2813 2816
rect 2754 2733 2757 2746
rect 2642 2713 2645 2726
rect 2658 2686 2661 2726
rect 2682 2713 2685 2726
rect 2738 2703 2741 2726
rect 2786 2706 2789 2726
rect 2786 2703 2793 2706
rect 2658 2683 2677 2686
rect 2634 2663 2645 2666
rect 2642 2546 2645 2663
rect 2666 2593 2669 2606
rect 2634 2543 2645 2546
rect 2602 2513 2613 2516
rect 2586 2413 2597 2416
rect 2562 2403 2573 2406
rect 2570 2336 2573 2403
rect 2554 2333 2573 2336
rect 2554 2226 2557 2333
rect 2554 2223 2573 2226
rect 2514 2183 2533 2186
rect 2466 2133 2477 2136
rect 2466 2113 2469 2133
rect 2490 2046 2493 2176
rect 2514 2136 2517 2176
rect 2506 2133 2517 2136
rect 2490 2043 2497 2046
rect 2466 2003 2469 2026
rect 2482 2013 2485 2036
rect 2442 1943 2453 1946
rect 2442 1923 2445 1943
rect 2434 1903 2445 1906
rect 2422 1893 2429 1896
rect 2406 1883 2413 1886
rect 2406 1786 2409 1883
rect 2418 1803 2421 1836
rect 2426 1813 2429 1893
rect 2442 1806 2445 1903
rect 2434 1803 2445 1806
rect 2458 1803 2461 1926
rect 2474 1916 2477 1926
rect 2482 1923 2485 1986
rect 2466 1896 2469 1916
rect 2474 1913 2485 1916
rect 2494 1906 2497 2043
rect 2490 1903 2497 1906
rect 2466 1893 2477 1896
rect 2474 1836 2477 1893
rect 2466 1833 2477 1836
rect 2402 1783 2409 1786
rect 2402 1723 2405 1783
rect 2434 1733 2437 1803
rect 2466 1766 2469 1833
rect 2466 1763 2477 1766
rect 2298 1696 2301 1716
rect 2298 1693 2309 1696
rect 2282 1683 2293 1686
rect 2274 1653 2281 1656
rect 2242 1593 2249 1596
rect 2246 1526 2249 1593
rect 2278 1576 2281 1653
rect 2290 1613 2293 1683
rect 2306 1636 2309 1693
rect 2298 1633 2309 1636
rect 2298 1603 2301 1633
rect 2322 1616 2325 1723
rect 2362 1676 2365 1723
rect 2426 1716 2429 1726
rect 2426 1713 2437 1716
rect 2442 1713 2445 1736
rect 2474 1733 2477 1763
rect 2314 1613 2325 1616
rect 2354 1673 2365 1676
rect 2354 1616 2357 1673
rect 2354 1613 2365 1616
rect 2274 1573 2281 1576
rect 2242 1523 2249 1526
rect 2242 1506 2245 1523
rect 2210 1483 2213 1506
rect 2218 1503 2245 1506
rect 2218 1413 2221 1503
rect 2258 1446 2261 1566
rect 2258 1443 2265 1446
rect 2250 1413 2253 1436
rect 2194 1373 2205 1376
rect 2202 1336 2205 1373
rect 2202 1333 2221 1336
rect 2178 1323 2197 1326
rect 2202 1323 2205 1333
rect 2178 1296 2181 1323
rect 2186 1313 2197 1316
rect 2210 1313 2213 1326
rect 2178 1293 2185 1296
rect 2182 1146 2185 1293
rect 2194 1183 2197 1313
rect 2218 1213 2221 1333
rect 2250 1306 2253 1406
rect 2262 1366 2265 1443
rect 2246 1303 2253 1306
rect 2258 1363 2265 1366
rect 2246 1236 2249 1303
rect 2246 1233 2253 1236
rect 2218 1193 2221 1206
rect 2242 1196 2245 1216
rect 2238 1193 2245 1196
rect 2178 1143 2185 1146
rect 2138 1023 2141 1036
rect 2146 1006 2149 1046
rect 2162 1026 2165 1046
rect 2142 1003 2149 1006
rect 2154 1023 2165 1026
rect 2034 576 2037 596
rect 2050 586 2053 606
rect 2050 583 2061 586
rect 1970 533 1973 546
rect 1962 523 1973 526
rect 1970 436 1973 523
rect 1962 433 1973 436
rect 1946 313 1949 326
rect 1954 253 1957 336
rect 1962 326 1965 433
rect 1970 333 1973 346
rect 1978 333 1981 526
rect 1994 413 1997 446
rect 1962 323 1973 326
rect 1962 306 1965 323
rect 1962 303 1969 306
rect 1966 236 1969 303
rect 1962 233 1969 236
rect 1914 203 1917 216
rect 1930 203 1933 226
rect 1946 193 1949 206
rect 1954 123 1957 216
rect 1962 203 1965 233
rect 1978 206 1981 236
rect 1986 213 1989 226
rect 1978 203 1989 206
rect 1994 203 1997 406
rect 2002 403 2005 576
rect 2010 533 2013 546
rect 2026 533 2029 576
rect 2034 573 2053 576
rect 2018 523 2029 526
rect 2010 413 2013 426
rect 2018 396 2021 446
rect 2034 443 2037 566
rect 2042 523 2045 536
rect 2026 413 2029 436
rect 2014 393 2021 396
rect 2014 336 2017 393
rect 2026 383 2029 406
rect 2034 403 2037 426
rect 2026 343 2045 346
rect 2002 316 2005 336
rect 2014 333 2021 336
rect 2002 313 2009 316
rect 2006 226 2009 313
rect 2006 223 2013 226
rect 1986 133 1989 203
rect 2002 183 2005 216
rect 2010 213 2013 223
rect 1514 93 1517 113
rect 1986 76 1989 126
rect 2018 123 2021 333
rect 2026 323 2029 343
rect 2034 323 2037 336
rect 2042 333 2045 343
rect 2050 316 2053 573
rect 2058 553 2061 583
rect 2066 536 2069 926
rect 2090 866 2093 936
rect 2106 903 2109 916
rect 2090 863 2101 866
rect 2074 816 2077 836
rect 2074 813 2081 816
rect 2078 746 2081 813
rect 2074 743 2081 746
rect 2074 723 2077 743
rect 2074 593 2077 716
rect 2098 656 2101 863
rect 2130 826 2133 956
rect 2142 906 2145 1003
rect 2154 913 2157 1023
rect 2170 1006 2173 1086
rect 2178 1023 2181 1143
rect 2194 1113 2197 1126
rect 2186 1093 2189 1106
rect 2194 1016 2197 1106
rect 2178 1013 2197 1016
rect 2170 1003 2181 1006
rect 2142 903 2149 906
rect 2162 903 2165 916
rect 2130 823 2137 826
rect 2090 653 2101 656
rect 2062 533 2069 536
rect 2062 346 2065 533
rect 2062 343 2069 346
rect 2034 313 2053 316
rect 2034 166 2037 313
rect 2058 263 2061 326
rect 2066 256 2069 343
rect 2050 253 2069 256
rect 2050 176 2053 253
rect 2050 173 2061 176
rect 2030 163 2037 166
rect 1978 73 1989 76
rect 1978 16 1981 73
rect 1978 13 1989 16
rect 1986 0 1989 13
rect 2002 0 2005 116
rect 2030 86 2033 163
rect 2050 113 2053 126
rect 2058 123 2061 173
rect 2066 96 2069 176
rect 2074 103 2077 566
rect 2090 556 2093 653
rect 2090 553 2109 556
rect 2082 396 2085 536
rect 2090 513 2093 526
rect 2098 523 2101 546
rect 2106 506 2109 553
rect 2102 503 2109 506
rect 2102 436 2105 503
rect 2102 433 2109 436
rect 2090 413 2093 426
rect 2082 393 2089 396
rect 2086 196 2089 393
rect 2098 383 2101 416
rect 2106 343 2109 433
rect 2114 366 2117 616
rect 2122 563 2125 816
rect 2134 746 2137 823
rect 2130 743 2137 746
rect 2130 533 2133 743
rect 2138 566 2141 726
rect 2146 723 2149 903
rect 2178 896 2181 1003
rect 2186 903 2189 1013
rect 2194 993 2197 1006
rect 2178 893 2189 896
rect 2178 813 2181 886
rect 2186 813 2189 893
rect 2170 733 2173 746
rect 2194 723 2197 986
rect 2202 786 2205 1136
rect 2210 1083 2213 1186
rect 2218 1103 2221 1116
rect 2210 803 2213 1056
rect 2218 993 2221 1096
rect 2226 973 2229 1166
rect 2238 1066 2241 1193
rect 2234 1063 2241 1066
rect 2218 903 2221 916
rect 2202 783 2209 786
rect 2206 716 2209 783
rect 2170 613 2173 716
rect 2202 713 2209 716
rect 2202 696 2205 713
rect 2194 693 2205 696
rect 2194 576 2197 693
rect 2226 686 2229 966
rect 2234 913 2237 1063
rect 2250 983 2253 1233
rect 2258 1166 2261 1363
rect 2274 1346 2277 1573
rect 2298 1356 2301 1546
rect 2314 1523 2317 1613
rect 2338 1523 2341 1596
rect 2362 1593 2365 1613
rect 2370 1586 2373 1666
rect 2354 1583 2373 1586
rect 2354 1486 2357 1583
rect 2394 1543 2397 1606
rect 2434 1556 2437 1713
rect 2442 1613 2445 1626
rect 2482 1613 2485 1726
rect 2490 1713 2493 1903
rect 2506 1753 2509 2126
rect 2530 2006 2533 2183
rect 2562 2113 2565 2136
rect 2522 2003 2533 2006
rect 2522 1923 2525 2003
rect 2522 1813 2525 1866
rect 2546 1853 2549 1986
rect 2554 1933 2557 2006
rect 2570 2003 2573 2223
rect 2578 2213 2581 2326
rect 2578 2123 2581 2136
rect 2594 2053 2597 2413
rect 2586 2013 2597 2016
rect 2602 2013 2605 2026
rect 2610 1996 2613 2513
rect 2626 2403 2629 2436
rect 2626 2203 2629 2216
rect 2634 2146 2637 2543
rect 2658 2513 2661 2526
rect 2674 2486 2677 2683
rect 2682 2593 2685 2616
rect 2698 2603 2701 2616
rect 2706 2583 2709 2596
rect 2746 2583 2749 2606
rect 2762 2603 2765 2656
rect 2762 2533 2765 2596
rect 2770 2526 2773 2606
rect 2698 2513 2701 2526
rect 2754 2523 2773 2526
rect 2754 2493 2757 2523
rect 2674 2483 2701 2486
rect 2642 2403 2645 2426
rect 2682 2413 2685 2426
rect 2626 2143 2637 2146
rect 2618 2123 2621 2136
rect 2602 1993 2613 1996
rect 2530 1803 2533 1816
rect 2554 1746 2557 1836
rect 2562 1813 2565 1926
rect 2570 1916 2573 1936
rect 2570 1913 2581 1916
rect 2570 1803 2573 1816
rect 2578 1813 2581 1913
rect 2602 1876 2605 1993
rect 2618 1923 2621 2056
rect 2602 1873 2613 1876
rect 2586 1806 2589 1856
rect 2610 1853 2613 1873
rect 2578 1803 2589 1806
rect 2610 1803 2613 1816
rect 2550 1743 2557 1746
rect 2434 1553 2445 1556
rect 2426 1533 2429 1546
rect 2354 1483 2365 1486
rect 2378 1483 2381 1526
rect 2442 1523 2445 1553
rect 2530 1493 2533 1726
rect 2538 1613 2541 1726
rect 2550 1696 2553 1743
rect 2550 1693 2557 1696
rect 2562 1693 2565 1736
rect 2570 1706 2573 1726
rect 2578 1713 2581 1803
rect 2626 1773 2629 2143
rect 2650 2136 2653 2326
rect 2682 2303 2685 2326
rect 2698 2323 2701 2483
rect 2778 2446 2781 2686
rect 2790 2606 2793 2703
rect 2786 2603 2793 2606
rect 2786 2523 2789 2603
rect 2802 2596 2805 2746
rect 2818 2603 2821 2616
rect 2802 2593 2809 2596
rect 2794 2533 2797 2586
rect 2806 2526 2809 2593
rect 2826 2526 2829 2843
rect 2842 2803 2845 2926
rect 2850 2793 2853 2946
rect 2858 2863 2861 2953
rect 2866 2913 2869 3006
rect 2878 2936 2881 3013
rect 2878 2933 2885 2936
rect 2882 2916 2885 2933
rect 2874 2913 2885 2916
rect 2890 2913 2893 3026
rect 2858 2813 2861 2826
rect 2874 2796 2877 2913
rect 2898 2903 2901 3153
rect 2906 3116 2909 3136
rect 2906 3113 2917 3116
rect 2914 3046 2917 3113
rect 2906 3043 2917 3046
rect 2906 3023 2909 3043
rect 2866 2793 2877 2796
rect 2842 2583 2845 2726
rect 2850 2706 2853 2766
rect 2866 2726 2869 2793
rect 2882 2746 2885 2806
rect 2890 2803 2893 2816
rect 2906 2753 2909 3006
rect 2914 2933 2917 3016
rect 2922 3003 2925 3016
rect 2914 2913 2917 2926
rect 2922 2923 2925 2936
rect 2922 2813 2925 2826
rect 2882 2743 2893 2746
rect 2866 2723 2877 2726
rect 2850 2703 2861 2706
rect 2858 2626 2861 2703
rect 2874 2636 2877 2723
rect 2882 2703 2885 2736
rect 2890 2656 2893 2743
rect 2914 2733 2917 2806
rect 2890 2653 2901 2656
rect 2850 2623 2861 2626
rect 2870 2633 2877 2636
rect 2802 2523 2809 2526
rect 2818 2523 2829 2526
rect 2770 2443 2781 2446
rect 2802 2443 2805 2523
rect 2850 2476 2853 2623
rect 2858 2533 2861 2606
rect 2870 2586 2873 2633
rect 2870 2583 2877 2586
rect 2866 2543 2869 2566
rect 2842 2473 2853 2476
rect 2722 2413 2725 2426
rect 2722 2303 2725 2326
rect 2770 2296 2773 2443
rect 2786 2413 2789 2436
rect 2818 2403 2821 2436
rect 2826 2403 2829 2426
rect 2786 2363 2789 2396
rect 2786 2306 2789 2326
rect 2842 2323 2845 2473
rect 2874 2426 2877 2583
rect 2882 2543 2885 2626
rect 2890 2613 2893 2646
rect 2898 2636 2901 2653
rect 2898 2633 2905 2636
rect 2890 2583 2893 2606
rect 2890 2513 2893 2566
rect 2902 2556 2905 2633
rect 2930 2623 2933 3116
rect 2938 2833 2941 3203
rect 2954 3176 2957 3363
rect 2946 3173 2957 3176
rect 2946 3046 2949 3173
rect 2954 3093 2957 3136
rect 2962 3133 2965 3156
rect 2970 3063 2973 3316
rect 2986 3286 2989 3326
rect 2994 3323 2997 3336
rect 3002 3303 3005 3336
rect 3010 3293 3013 3316
rect 3026 3296 3029 3363
rect 3018 3293 3029 3296
rect 3058 3363 3069 3366
rect 2986 3283 2997 3286
rect 2994 3216 2997 3283
rect 3018 3273 3021 3293
rect 3058 3286 3061 3363
rect 3074 3313 3077 3326
rect 3058 3283 3069 3286
rect 3066 3266 3069 3283
rect 2994 3213 3005 3216
rect 2994 3146 2997 3166
rect 2986 3143 2997 3146
rect 2986 3046 2989 3143
rect 3002 3126 3005 3213
rect 3034 3133 3037 3216
rect 3042 3203 3053 3206
rect 3058 3186 3061 3266
rect 3066 3263 3073 3266
rect 3070 3206 3073 3263
rect 3054 3183 3061 3186
rect 3066 3203 3073 3206
rect 3002 3123 3021 3126
rect 2946 3043 2957 3046
rect 2986 3043 2997 3046
rect 2954 2956 2957 3043
rect 2994 3023 2997 3043
rect 2946 2953 2957 2956
rect 2946 2826 2949 2953
rect 2938 2823 2949 2826
rect 2954 2823 2957 2936
rect 2970 2903 2973 2916
rect 3002 2846 3005 3123
rect 3010 3003 3013 3016
rect 2994 2843 3005 2846
rect 2938 2786 2941 2823
rect 2946 2803 2949 2816
rect 2938 2783 2949 2786
rect 2946 2646 2949 2783
rect 2938 2643 2949 2646
rect 2898 2553 2905 2556
rect 2898 2463 2901 2553
rect 2906 2523 2909 2536
rect 2914 2523 2917 2586
rect 2922 2563 2925 2606
rect 2922 2533 2925 2546
rect 2938 2506 2941 2643
rect 2930 2503 2941 2506
rect 2930 2426 2933 2503
rect 2874 2423 2885 2426
rect 2930 2423 2941 2426
rect 2866 2393 2869 2416
rect 2866 2343 2869 2376
rect 2882 2346 2885 2423
rect 2874 2343 2885 2346
rect 2786 2303 2797 2306
rect 2770 2293 2781 2296
rect 2778 2276 2781 2293
rect 2770 2273 2781 2276
rect 2658 2143 2669 2146
rect 2634 2066 2637 2136
rect 2650 2133 2669 2136
rect 2674 2133 2677 2216
rect 2642 2113 2645 2126
rect 2634 2063 2641 2066
rect 2638 2006 2641 2063
rect 2658 2053 2661 2126
rect 2634 2003 2641 2006
rect 2650 2003 2653 2026
rect 2634 1923 2637 2003
rect 2666 1906 2669 2133
rect 2714 2056 2717 2136
rect 2730 2133 2733 2216
rect 2770 2206 2773 2273
rect 2794 2236 2797 2303
rect 2786 2233 2797 2236
rect 2786 2213 2789 2233
rect 2802 2206 2805 2216
rect 2866 2213 2869 2226
rect 2770 2203 2781 2206
rect 2802 2203 2813 2206
rect 2778 2156 2781 2203
rect 2778 2153 2789 2156
rect 2770 2103 2773 2146
rect 2786 2096 2789 2153
rect 2810 2116 2813 2203
rect 2826 2123 2829 2206
rect 2842 2133 2845 2166
rect 2810 2113 2821 2116
rect 2706 2053 2717 2056
rect 2778 2093 2789 2096
rect 2690 2013 2693 2036
rect 2706 1976 2709 2053
rect 2746 2013 2749 2026
rect 2706 1973 2725 1976
rect 2658 1903 2669 1906
rect 2658 1803 2661 1903
rect 2722 1873 2725 1973
rect 2730 1913 2733 2006
rect 2778 1976 2781 2093
rect 2770 1973 2781 1976
rect 2738 1923 2741 1936
rect 2770 1916 2773 1973
rect 2794 1923 2797 1966
rect 2818 1963 2821 2113
rect 2858 2106 2861 2126
rect 2850 2103 2861 2106
rect 2850 2026 2853 2103
rect 2850 2023 2861 2026
rect 2858 2003 2861 2023
rect 2770 1913 2781 1916
rect 2818 1913 2821 1936
rect 2730 1823 2741 1826
rect 2722 1803 2741 1806
rect 2594 1713 2597 1726
rect 2602 1706 2605 1736
rect 2610 1723 2613 1736
rect 2570 1703 2589 1706
rect 2594 1703 2605 1706
rect 2626 1703 2629 1726
rect 2642 1703 2645 1716
rect 2650 1713 2653 1726
rect 2666 1713 2669 1776
rect 2674 1713 2677 1726
rect 2722 1713 2725 1726
rect 2738 1713 2741 1803
rect 2546 1506 2549 1606
rect 2554 1563 2557 1693
rect 2570 1533 2573 1546
rect 2542 1503 2549 1506
rect 2266 1343 2277 1346
rect 2290 1353 2301 1356
rect 2266 1286 2269 1343
rect 2290 1333 2293 1353
rect 2338 1336 2341 1476
rect 2362 1446 2365 1483
rect 2362 1443 2373 1446
rect 2370 1396 2373 1443
rect 2542 1436 2545 1503
rect 2542 1433 2549 1436
rect 2362 1393 2373 1396
rect 2266 1283 2293 1286
rect 2266 1213 2269 1276
rect 2290 1216 2293 1283
rect 2306 1273 2309 1336
rect 2330 1333 2341 1336
rect 2282 1213 2293 1216
rect 2306 1213 2309 1256
rect 2314 1213 2317 1316
rect 2258 1163 2269 1166
rect 2266 1056 2269 1163
rect 2282 1113 2285 1213
rect 2258 1053 2269 1056
rect 2234 853 2237 906
rect 2250 846 2253 976
rect 2258 923 2261 1053
rect 2266 923 2269 1036
rect 2274 1013 2277 1026
rect 2298 963 2301 1196
rect 2322 1096 2325 1246
rect 2330 1193 2333 1333
rect 2338 1136 2341 1326
rect 2346 1243 2349 1316
rect 2354 1303 2357 1336
rect 2346 1203 2357 1206
rect 2338 1133 2349 1136
rect 2314 1093 2325 1096
rect 2314 1046 2317 1093
rect 2314 1043 2325 1046
rect 2314 1003 2317 1026
rect 2274 906 2277 926
rect 2270 903 2277 906
rect 2250 843 2261 846
rect 2258 796 2261 843
rect 2270 836 2273 903
rect 2282 883 2285 936
rect 2290 913 2293 936
rect 2306 923 2309 936
rect 2270 833 2277 836
rect 2274 813 2277 833
rect 2306 813 2309 916
rect 2322 903 2325 1043
rect 2330 1023 2333 1126
rect 2346 1066 2349 1133
rect 2362 1086 2365 1393
rect 2370 1223 2373 1326
rect 2378 1146 2381 1366
rect 2386 1316 2389 1416
rect 2394 1333 2397 1356
rect 2418 1353 2421 1416
rect 2450 1356 2453 1396
rect 2450 1353 2469 1356
rect 2402 1333 2405 1346
rect 2410 1326 2413 1346
rect 2402 1323 2413 1326
rect 2466 1323 2469 1353
rect 2386 1313 2393 1316
rect 2390 1226 2393 1313
rect 2402 1296 2405 1323
rect 2402 1293 2413 1296
rect 2410 1236 2413 1293
rect 2386 1223 2393 1226
rect 2402 1233 2413 1236
rect 2386 1203 2389 1223
rect 2402 1213 2405 1233
rect 2434 1213 2437 1306
rect 2418 1203 2437 1206
rect 2378 1143 2385 1146
rect 2370 1093 2373 1136
rect 2362 1083 2373 1086
rect 2338 1063 2349 1066
rect 2338 1046 2341 1063
rect 2338 1043 2349 1046
rect 2346 976 2349 1043
rect 2354 1013 2357 1046
rect 2370 1013 2373 1083
rect 2382 1076 2385 1143
rect 2394 1123 2397 1166
rect 2378 1073 2385 1076
rect 2378 1053 2381 1073
rect 2354 1003 2365 1006
rect 2330 973 2349 976
rect 2314 813 2317 886
rect 2330 833 2333 973
rect 2346 916 2349 936
rect 2354 933 2357 996
rect 2402 993 2405 1126
rect 2434 1123 2437 1203
rect 2450 1193 2453 1226
rect 2458 1213 2461 1306
rect 2482 1203 2485 1216
rect 2490 1213 2493 1226
rect 2498 1216 2501 1326
rect 2522 1323 2525 1416
rect 2530 1253 2533 1356
rect 2538 1343 2541 1416
rect 2546 1363 2549 1433
rect 2554 1393 2557 1496
rect 2586 1413 2589 1526
rect 2594 1513 2597 1703
rect 2618 1656 2621 1696
rect 2650 1693 2653 1706
rect 2674 1693 2677 1706
rect 2614 1653 2621 1656
rect 2602 1456 2605 1616
rect 2614 1586 2617 1653
rect 2614 1583 2621 1586
rect 2650 1583 2653 1656
rect 2698 1633 2717 1636
rect 2658 1613 2661 1626
rect 2698 1613 2701 1633
rect 2618 1566 2621 1583
rect 2618 1563 2629 1566
rect 2626 1456 2629 1563
rect 2602 1453 2613 1456
rect 2498 1213 2509 1216
rect 2498 1193 2501 1206
rect 2490 1126 2493 1146
rect 2506 1133 2509 1213
rect 2514 1203 2517 1226
rect 2522 1203 2525 1216
rect 2546 1203 2549 1236
rect 2490 1123 2501 1126
rect 2450 1103 2469 1106
rect 2466 1086 2469 1103
rect 2462 1083 2469 1086
rect 2462 1026 2465 1083
rect 2462 1023 2469 1026
rect 2434 1003 2437 1016
rect 2450 993 2453 1006
rect 2466 1003 2469 1023
rect 2474 1013 2477 1106
rect 2498 1103 2501 1123
rect 2514 1106 2517 1146
rect 2538 1123 2549 1126
rect 2554 1123 2557 1216
rect 2562 1213 2565 1326
rect 2578 1213 2581 1226
rect 2586 1213 2589 1336
rect 2602 1316 2605 1336
rect 2598 1313 2605 1316
rect 2598 1216 2601 1313
rect 2598 1213 2605 1216
rect 2570 1133 2573 1206
rect 2506 1103 2517 1106
rect 2362 926 2365 946
rect 2342 913 2349 916
rect 2354 923 2365 926
rect 2314 796 2317 806
rect 2250 793 2261 796
rect 2298 793 2317 796
rect 2250 736 2253 793
rect 2298 783 2301 793
rect 2322 786 2325 816
rect 2330 813 2333 826
rect 2342 816 2345 913
rect 2354 826 2357 923
rect 2418 846 2421 876
rect 2410 843 2421 846
rect 2354 823 2361 826
rect 2342 813 2349 816
rect 2306 783 2325 786
rect 2218 683 2229 686
rect 2242 733 2253 736
rect 2274 733 2277 746
rect 2218 583 2221 683
rect 2242 646 2245 733
rect 2250 713 2253 726
rect 2274 656 2277 726
rect 2290 713 2293 736
rect 2306 713 2309 783
rect 2346 733 2349 813
rect 2358 736 2361 823
rect 2354 733 2361 736
rect 2354 713 2357 733
rect 2370 696 2373 836
rect 2378 736 2381 816
rect 2410 766 2413 843
rect 2450 836 2453 926
rect 2466 913 2469 936
rect 2474 873 2477 1006
rect 2482 1003 2485 1016
rect 2498 1003 2501 1086
rect 2506 1003 2509 1103
rect 2530 1013 2533 1116
rect 2546 1046 2549 1123
rect 2562 1113 2565 1126
rect 2546 1043 2557 1046
rect 2602 1043 2605 1213
rect 2610 1173 2613 1453
rect 2622 1453 2629 1456
rect 2622 1376 2625 1453
rect 2634 1413 2637 1426
rect 2658 1403 2661 1416
rect 2618 1373 2625 1376
rect 2618 1353 2621 1373
rect 2618 1313 2621 1326
rect 2618 1133 2621 1246
rect 2634 1233 2637 1326
rect 2642 1243 2645 1336
rect 2650 1323 2653 1376
rect 2674 1373 2677 1416
rect 2682 1413 2685 1606
rect 2706 1603 2709 1626
rect 2714 1613 2717 1633
rect 2714 1576 2717 1606
rect 2722 1583 2725 1596
rect 2706 1573 2717 1576
rect 2706 1466 2709 1573
rect 2706 1463 2717 1466
rect 2714 1446 2717 1463
rect 2714 1443 2721 1446
rect 2718 1386 2721 1443
rect 2714 1383 2721 1386
rect 2658 1333 2661 1356
rect 2666 1293 2669 1326
rect 2674 1256 2677 1366
rect 2714 1363 2717 1383
rect 2730 1373 2733 1546
rect 2738 1413 2741 1536
rect 2746 1523 2749 1596
rect 2754 1583 2757 1806
rect 2778 1543 2781 1913
rect 2874 1863 2877 2343
rect 2890 2313 2893 2326
rect 2882 2193 2885 2206
rect 2890 2203 2893 2216
rect 2898 2206 2901 2406
rect 2914 2393 2917 2406
rect 2938 2403 2941 2423
rect 2906 2326 2909 2336
rect 2906 2323 2925 2326
rect 2930 2323 2933 2336
rect 2922 2313 2933 2316
rect 2954 2313 2957 2626
rect 2962 2623 2965 2836
rect 2994 2676 2997 2843
rect 3026 2826 3029 3126
rect 3042 3073 3045 3136
rect 3054 3126 3057 3183
rect 3066 3133 3069 3203
rect 3054 3123 3061 3126
rect 3074 3123 3077 3186
rect 3082 3163 3085 3456
rect 3090 3366 3093 3633
rect 3098 3383 3101 3616
rect 3106 3413 3109 3536
rect 3114 3486 3117 3783
rect 3138 3736 3141 3793
rect 3154 3776 3157 3923
rect 3170 3906 3173 4106
rect 3186 4103 3189 4303
rect 3218 4286 3221 4336
rect 3210 4283 3221 4286
rect 3210 4226 3213 4283
rect 3210 4223 3221 4226
rect 3194 4173 3197 4206
rect 3218 4143 3221 4223
rect 3226 4183 3229 4416
rect 3234 4333 3237 4366
rect 3242 4323 3245 4386
rect 3250 4333 3253 4433
rect 3258 4413 3261 4426
rect 3282 4353 3285 4406
rect 3306 4363 3309 4416
rect 3362 4376 3365 4453
rect 3386 4436 3389 4516
rect 3402 4513 3405 4526
rect 3426 4523 3429 4566
rect 3434 4533 3445 4536
rect 3418 4493 3421 4506
rect 3354 4373 3365 4376
rect 3378 4433 3389 4436
rect 3354 4356 3357 4373
rect 3242 4296 3245 4316
rect 3242 4293 3253 4296
rect 3250 4246 3253 4293
rect 3242 4243 3253 4246
rect 3234 4213 3237 4226
rect 3242 4203 3245 4243
rect 3250 4193 3253 4216
rect 3258 4213 3261 4226
rect 3274 4193 3277 4276
rect 3178 4003 3181 4026
rect 3186 3983 3189 4016
rect 3194 4003 3197 4016
rect 3186 3933 3189 3946
rect 3202 3906 3205 4106
rect 3226 4103 3229 4136
rect 3218 3933 3221 3996
rect 3242 3993 3245 4186
rect 3306 4183 3309 4356
rect 3346 4353 3357 4356
rect 3330 4313 3333 4326
rect 3346 4286 3349 4353
rect 3378 4316 3381 4433
rect 3394 4423 3405 4426
rect 3394 4346 3397 4423
rect 3402 4383 3405 4416
rect 3394 4343 3401 4346
rect 3374 4313 3381 4316
rect 3346 4283 3357 4286
rect 3346 4193 3349 4216
rect 3354 4176 3357 4283
rect 3374 4236 3377 4313
rect 3374 4233 3381 4236
rect 3362 4203 3365 4226
rect 3346 4173 3357 4176
rect 3266 4113 3269 4126
rect 3290 4056 3293 4146
rect 3346 4116 3349 4173
rect 3370 4163 3373 4216
rect 3362 4123 3365 4136
rect 3346 4113 3357 4116
rect 3282 4053 3293 4056
rect 3266 4013 3269 4026
rect 3282 3976 3285 4053
rect 3346 3983 3349 4016
rect 3282 3973 3289 3976
rect 3242 3906 3245 3926
rect 3170 3903 3181 3906
rect 3202 3903 3213 3906
rect 3242 3903 3253 3906
rect 3178 3846 3181 3903
rect 3170 3843 3181 3846
rect 3170 3813 3173 3843
rect 3202 3793 3205 3806
rect 3154 3773 3173 3776
rect 3130 3733 3141 3736
rect 3170 3733 3173 3773
rect 3130 3686 3133 3733
rect 3146 3696 3149 3726
rect 3146 3693 3157 3696
rect 3130 3683 3141 3686
rect 3122 3613 3125 3626
rect 3130 3593 3133 3606
rect 3122 3503 3125 3526
rect 3138 3523 3141 3683
rect 3154 3636 3157 3693
rect 3194 3636 3197 3726
rect 3210 3676 3213 3903
rect 3226 3813 3229 3846
rect 3218 3803 3229 3806
rect 3234 3803 3237 3856
rect 3250 3816 3253 3903
rect 3286 3896 3289 3973
rect 3354 3966 3357 4113
rect 3378 4106 3381 4233
rect 3386 4223 3389 4326
rect 3398 4296 3401 4343
rect 3398 4293 3405 4296
rect 3350 3963 3357 3966
rect 3370 4103 3381 4106
rect 3298 3906 3301 3926
rect 3338 3906 3341 3926
rect 3298 3903 3309 3906
rect 3286 3893 3293 3896
rect 3242 3813 3253 3816
rect 3282 3813 3285 3846
rect 3226 3796 3229 3803
rect 3242 3796 3245 3813
rect 3226 3793 3245 3796
rect 3250 3676 3253 3726
rect 3210 3673 3221 3676
rect 3146 3633 3157 3636
rect 3186 3633 3197 3636
rect 3146 3603 3149 3633
rect 3186 3616 3189 3633
rect 3154 3523 3157 3616
rect 3182 3613 3189 3616
rect 3114 3483 3121 3486
rect 3162 3483 3165 3536
rect 3118 3406 3121 3483
rect 3170 3426 3173 3606
rect 3182 3556 3185 3613
rect 3194 3593 3197 3606
rect 3182 3553 3189 3556
rect 3186 3536 3189 3553
rect 3178 3533 3189 3536
rect 3194 3533 3197 3576
rect 3218 3536 3221 3673
rect 3242 3673 3253 3676
rect 3242 3626 3245 3673
rect 3266 3636 3269 3796
rect 3290 3786 3293 3893
rect 3306 3826 3309 3903
rect 3298 3823 3309 3826
rect 3330 3903 3341 3906
rect 3330 3826 3333 3903
rect 3350 3886 3353 3963
rect 3350 3883 3357 3886
rect 3330 3823 3341 3826
rect 3298 3803 3301 3823
rect 3338 3803 3341 3823
rect 3354 3786 3357 3883
rect 3370 3876 3373 4103
rect 3378 4003 3381 4036
rect 3386 4013 3389 4216
rect 3402 4156 3405 4293
rect 3418 4203 3421 4466
rect 3426 4433 3429 4446
rect 3434 4413 3437 4486
rect 3482 4466 3485 4556
rect 3506 4523 3509 4576
rect 3514 4533 3517 4606
rect 3530 4593 3533 4616
rect 3586 4583 3589 4616
rect 3618 4613 3621 4626
rect 3626 4573 3629 4616
rect 3634 4593 3637 4606
rect 3530 4533 3533 4546
rect 3490 4473 3493 4516
rect 3522 4513 3525 4526
rect 3538 4513 3541 4536
rect 3602 4533 3605 4556
rect 3642 4533 3645 4626
rect 3650 4543 3653 4606
rect 3682 4603 3685 4636
rect 3714 4586 3717 4636
rect 3730 4603 3733 4616
rect 3706 4583 3717 4586
rect 3482 4463 3493 4466
rect 3474 4423 3477 4436
rect 3490 4433 3493 4463
rect 3482 4366 3485 4426
rect 3498 4413 3501 4446
rect 3506 4423 3509 4456
rect 3482 4363 3489 4366
rect 3450 4213 3453 4246
rect 3394 4153 3405 4156
rect 3366 3873 3373 3876
rect 3366 3806 3369 3873
rect 3366 3803 3373 3806
rect 3370 3786 3373 3803
rect 3378 3793 3381 3966
rect 3386 3923 3389 3946
rect 3394 3876 3397 4153
rect 3402 4053 3405 4136
rect 3418 4033 3421 4126
rect 3402 4003 3405 4016
rect 3410 3963 3413 4026
rect 3426 4013 3429 4026
rect 3418 3906 3421 3936
rect 3434 3906 3437 4206
rect 3442 4163 3445 4206
rect 3458 4203 3461 4326
rect 3486 4286 3489 4363
rect 3514 4333 3517 4416
rect 3498 4306 3501 4326
rect 3498 4303 3509 4306
rect 3482 4283 3489 4286
rect 3482 4223 3485 4283
rect 3506 4246 3509 4303
rect 3554 4256 3557 4526
rect 3570 4503 3573 4526
rect 3586 4453 3589 4526
rect 3642 4513 3645 4526
rect 3650 4503 3653 4526
rect 3666 4433 3669 4526
rect 3682 4496 3685 4526
rect 3706 4516 3709 4583
rect 3722 4523 3725 4586
rect 3730 4533 3733 4546
rect 3738 4523 3741 4536
rect 3754 4533 3757 4606
rect 3770 4533 3773 4576
rect 3778 4526 3781 4616
rect 3818 4603 3821 4636
rect 3762 4523 3781 4526
rect 3706 4513 3717 4516
rect 3682 4493 3693 4496
rect 3690 4436 3693 4493
rect 3682 4433 3693 4436
rect 3570 4343 3573 4416
rect 3682 4413 3685 4433
rect 3594 4346 3597 4406
rect 3698 4356 3701 4406
rect 3586 4343 3597 4346
rect 3586 4296 3589 4343
rect 3586 4293 3597 4296
rect 3554 4253 3565 4256
rect 3498 4243 3509 4246
rect 3466 4213 3485 4216
rect 3474 4136 3477 4206
rect 3442 4023 3445 4046
rect 3450 4013 3453 4136
rect 3458 4123 3461 4136
rect 3466 4133 3477 4136
rect 3482 4133 3485 4213
rect 3498 4203 3501 4243
rect 3466 4106 3469 4133
rect 3514 4126 3517 4226
rect 3530 4183 3533 4206
rect 3538 4166 3541 4246
rect 3462 4103 3469 4106
rect 3462 4026 3465 4103
rect 3462 4023 3469 4026
rect 3474 4023 3477 4126
rect 3490 4076 3493 4126
rect 3510 4123 3517 4126
rect 3534 4163 3541 4166
rect 3486 4073 3493 4076
rect 3466 4006 3469 4023
rect 3486 4016 3489 4073
rect 3498 4023 3501 4106
rect 3486 4013 3493 4016
rect 3466 4003 3477 4006
rect 3418 3903 3437 3906
rect 3434 3876 3437 3903
rect 3394 3873 3405 3876
rect 3402 3816 3405 3873
rect 3394 3813 3405 3816
rect 3426 3873 3437 3876
rect 3290 3783 3309 3786
rect 3262 3633 3269 3636
rect 3282 3633 3285 3716
rect 3306 3656 3309 3783
rect 3346 3783 3357 3786
rect 3346 3716 3349 3783
rect 3362 3723 3365 3786
rect 3370 3783 3381 3786
rect 3290 3653 3309 3656
rect 3290 3636 3293 3653
rect 3290 3633 3301 3636
rect 3242 3623 3253 3626
rect 3250 3603 3253 3623
rect 3262 3586 3265 3633
rect 3274 3596 3277 3626
rect 3290 3613 3293 3626
rect 3274 3593 3285 3596
rect 3262 3583 3269 3586
rect 3210 3533 3221 3536
rect 3186 3523 3197 3526
rect 3170 3423 3177 3426
rect 3114 3403 3121 3406
rect 3090 3363 3101 3366
rect 3098 3266 3101 3363
rect 3114 3346 3117 3403
rect 3138 3383 3141 3406
rect 3162 3376 3165 3416
rect 3146 3373 3165 3376
rect 3110 3343 3117 3346
rect 3110 3286 3113 3343
rect 3122 3313 3125 3336
rect 3130 3333 3133 3346
rect 3146 3333 3149 3373
rect 3174 3366 3177 3423
rect 3186 3366 3189 3516
rect 3202 3456 3205 3516
rect 3210 3513 3213 3533
rect 3250 3503 3253 3566
rect 3266 3536 3269 3583
rect 3266 3533 3273 3536
rect 3258 3513 3261 3526
rect 3270 3486 3273 3533
rect 3266 3483 3273 3486
rect 3202 3453 3209 3456
rect 3206 3376 3209 3453
rect 3202 3373 3209 3376
rect 3174 3363 3181 3366
rect 3186 3363 3193 3366
rect 3170 3333 3173 3356
rect 3110 3283 3117 3286
rect 3090 3263 3101 3266
rect 3114 3263 3117 3283
rect 3090 3243 3093 3263
rect 3090 3233 3109 3236
rect 3090 3213 3093 3233
rect 3098 3203 3101 3226
rect 3106 3216 3109 3233
rect 3106 3213 3117 3216
rect 3106 3136 3109 3206
rect 3122 3193 3125 3206
rect 3130 3183 3133 3326
rect 3154 3313 3157 3326
rect 3170 3313 3173 3326
rect 3138 3213 3141 3226
rect 3138 3166 3141 3206
rect 3178 3166 3181 3363
rect 3190 3246 3193 3363
rect 3058 3026 3061 3123
rect 3082 3113 3085 3136
rect 3098 3133 3109 3136
rect 3122 3163 3141 3166
rect 3174 3163 3181 3166
rect 3186 3243 3193 3246
rect 3122 3133 3125 3163
rect 3138 3133 3141 3156
rect 3090 3093 3093 3126
rect 3098 3026 3101 3133
rect 3162 3113 3165 3126
rect 3174 3096 3177 3163
rect 3186 3103 3189 3243
rect 3202 3226 3205 3373
rect 3218 3333 3221 3416
rect 3194 3223 3205 3226
rect 3194 3166 3197 3223
rect 3202 3193 3205 3216
rect 3194 3163 3205 3166
rect 3174 3093 3181 3096
rect 3178 3036 3181 3093
rect 3178 3033 3197 3036
rect 3058 3023 3069 3026
rect 3034 2993 3037 3006
rect 3042 2923 3045 3016
rect 3066 2916 3069 3023
rect 3090 3023 3101 3026
rect 3090 3003 3093 3023
rect 3098 2933 3101 3016
rect 3130 2993 3133 3016
rect 3178 2993 3181 3006
rect 3194 2986 3197 3033
rect 3186 2983 3197 2986
rect 3058 2913 3069 2916
rect 3058 2883 3061 2913
rect 3090 2896 3093 2916
rect 3186 2906 3189 2983
rect 3202 2913 3205 3163
rect 3226 3113 3229 3386
rect 3242 3383 3245 3406
rect 3266 3396 3269 3483
rect 3282 3436 3285 3593
rect 3298 3453 3301 3633
rect 3330 3626 3333 3716
rect 3346 3713 3357 3716
rect 3330 3623 3337 3626
rect 3346 3623 3349 3636
rect 3322 3526 3325 3616
rect 3334 3556 3337 3623
rect 3314 3523 3325 3526
rect 3330 3553 3337 3556
rect 3258 3393 3269 3396
rect 3274 3433 3285 3436
rect 3242 3336 3245 3356
rect 3238 3333 3245 3336
rect 3238 3246 3241 3333
rect 3238 3243 3245 3246
rect 3210 3003 3213 3106
rect 3218 3013 3221 3026
rect 3226 3013 3237 3016
rect 3226 3003 3237 3006
rect 3186 2903 3193 2906
rect 3090 2893 3101 2896
rect 3018 2823 3029 2826
rect 3018 2806 3021 2823
rect 3026 2813 3045 2816
rect 3002 2706 3005 2796
rect 3010 2723 3013 2806
rect 3018 2803 3025 2806
rect 3022 2726 3025 2803
rect 3034 2733 3037 2766
rect 3050 2743 3053 2806
rect 3022 2723 3029 2726
rect 3002 2703 3009 2706
rect 2986 2673 2997 2676
rect 2986 2616 2989 2673
rect 2962 2613 2973 2616
rect 2978 2613 2989 2616
rect 2970 2606 2973 2613
rect 2962 2596 2965 2606
rect 2970 2603 2989 2606
rect 2962 2593 2973 2596
rect 2970 2523 2973 2593
rect 2994 2533 2997 2666
rect 3006 2636 3009 2703
rect 3002 2633 3009 2636
rect 2970 2356 2973 2516
rect 2970 2353 2981 2356
rect 2898 2203 2909 2206
rect 2890 2123 2893 2136
rect 2898 2106 2901 2176
rect 2906 2123 2909 2203
rect 2914 2186 2917 2226
rect 2922 2223 2925 2313
rect 2922 2203 2925 2216
rect 2914 2183 2925 2186
rect 2922 2116 2925 2183
rect 2890 2103 2901 2106
rect 2906 2113 2925 2116
rect 2890 2046 2893 2103
rect 2890 2043 2901 2046
rect 2898 2023 2901 2043
rect 2906 1976 2909 2113
rect 2946 2096 2949 2306
rect 2962 2236 2965 2346
rect 2958 2233 2965 2236
rect 2958 2146 2961 2233
rect 2978 2226 2981 2353
rect 2994 2303 2997 2526
rect 3002 2513 3005 2633
rect 3010 2603 3013 2616
rect 3018 2603 3021 2626
rect 3026 2556 3029 2723
rect 3034 2613 3037 2646
rect 3058 2603 3061 2816
rect 3066 2813 3069 2826
rect 3074 2803 3077 2886
rect 3098 2846 3101 2893
rect 3090 2843 3101 2846
rect 3074 2723 3077 2746
rect 3090 2656 3093 2843
rect 3114 2766 3117 2806
rect 3162 2793 3165 2816
rect 3114 2763 3125 2766
rect 3082 2653 3093 2656
rect 3026 2553 3033 2556
rect 3018 2533 3021 2546
rect 3030 2506 3033 2553
rect 3042 2513 3045 2526
rect 3030 2503 3045 2506
rect 3026 2426 3029 2486
rect 3010 2403 3013 2426
rect 3022 2423 3029 2426
rect 3022 2356 3025 2423
rect 3042 2416 3045 2503
rect 3034 2413 3045 2416
rect 3022 2353 3029 2356
rect 3018 2273 3021 2336
rect 3026 2256 3029 2353
rect 2970 2223 2981 2226
rect 3022 2253 3029 2256
rect 2958 2143 2965 2146
rect 2938 2093 2949 2096
rect 2938 2036 2941 2093
rect 2954 2083 2957 2126
rect 2962 2053 2965 2143
rect 2970 2113 2973 2223
rect 2938 2033 2949 2036
rect 2922 1996 2925 2016
rect 2938 2003 2941 2016
rect 2946 2013 2949 2033
rect 2954 2003 2957 2026
rect 2898 1973 2909 1976
rect 2914 1993 2925 1996
rect 2802 1806 2805 1816
rect 2858 1813 2861 1826
rect 2898 1823 2901 1973
rect 2914 1906 2917 1993
rect 2970 1983 2973 2026
rect 2978 2013 2981 2206
rect 2986 2133 2997 2136
rect 2986 2013 2989 2116
rect 3002 2113 3005 2126
rect 3010 2123 3013 2196
rect 3022 2166 3025 2253
rect 3022 2163 3029 2166
rect 3018 2133 3021 2146
rect 2922 1943 2933 1946
rect 2970 1933 2973 1966
rect 2994 1913 2997 1926
rect 2914 1903 2925 1906
rect 2922 1846 2925 1903
rect 2914 1843 2925 1846
rect 2914 1826 2917 1843
rect 3002 1833 3005 2106
rect 3026 2103 3029 2163
rect 3018 1963 3021 2016
rect 3034 2013 3037 2413
rect 3050 2403 3053 2456
rect 3058 2323 3061 2596
rect 3082 2576 3085 2653
rect 3114 2613 3117 2626
rect 3082 2573 3093 2576
rect 3090 2556 3093 2573
rect 3090 2553 3101 2556
rect 3082 2486 3085 2526
rect 3066 2483 3085 2486
rect 3066 2403 3069 2483
rect 3098 2476 3101 2553
rect 3122 2543 3125 2763
rect 3170 2716 3173 2746
rect 3162 2713 3173 2716
rect 3162 2666 3165 2713
rect 3162 2663 3173 2666
rect 3154 2543 3157 2606
rect 3170 2576 3173 2663
rect 3166 2573 3173 2576
rect 3090 2473 3101 2476
rect 3074 2413 3077 2426
rect 3090 2396 3093 2473
rect 3106 2413 3109 2426
rect 3082 2393 3093 2396
rect 3042 2203 3045 2226
rect 3050 2193 3053 2266
rect 3066 2203 3069 2286
rect 3074 2213 3077 2276
rect 3082 2216 3085 2393
rect 3122 2366 3125 2426
rect 3138 2403 3141 2526
rect 3146 2513 3149 2526
rect 3166 2496 3169 2573
rect 3162 2493 3169 2496
rect 3162 2446 3165 2493
rect 3162 2443 3173 2446
rect 3170 2423 3173 2443
rect 3178 2416 3181 2896
rect 3190 2766 3193 2903
rect 3170 2413 3181 2416
rect 3186 2763 3193 2766
rect 3122 2363 3133 2366
rect 3090 2283 3093 2326
rect 3106 2226 3109 2326
rect 3130 2306 3133 2363
rect 3170 2353 3173 2413
rect 3186 2366 3189 2763
rect 3194 2733 3197 2746
rect 3194 2703 3197 2726
rect 3202 2696 3205 2836
rect 3210 2763 3213 2826
rect 3226 2816 3229 2996
rect 3226 2813 3233 2816
rect 3198 2693 3205 2696
rect 3198 2646 3201 2693
rect 3194 2643 3201 2646
rect 3194 2586 3197 2643
rect 3210 2593 3213 2746
rect 3218 2733 3221 2806
rect 3230 2766 3233 2813
rect 3242 2803 3245 3243
rect 3250 3076 3253 3376
rect 3258 3193 3261 3393
rect 3274 3363 3277 3433
rect 3282 3333 3285 3416
rect 3314 3373 3317 3523
rect 3322 3503 3325 3516
rect 3298 3333 3301 3356
rect 3266 3263 3269 3326
rect 3274 3306 3277 3326
rect 3282 3323 3309 3326
rect 3314 3306 3317 3366
rect 3322 3333 3325 3416
rect 3274 3303 3285 3306
rect 3258 3093 3261 3126
rect 3250 3073 3257 3076
rect 3254 2966 3257 3073
rect 3266 2986 3269 3246
rect 3282 3236 3285 3303
rect 3274 3233 3285 3236
rect 3306 3303 3317 3306
rect 3306 3236 3309 3303
rect 3330 3276 3333 3553
rect 3354 3536 3357 3713
rect 3370 3703 3373 3776
rect 3370 3613 3373 3626
rect 3362 3603 3373 3606
rect 3378 3586 3381 3783
rect 3374 3583 3381 3586
rect 3338 3523 3341 3536
rect 3354 3533 3365 3536
rect 3346 3513 3349 3526
rect 3338 3383 3341 3416
rect 3346 3413 3349 3496
rect 3362 3446 3365 3533
rect 3354 3443 3365 3446
rect 3330 3273 3341 3276
rect 3306 3233 3317 3236
rect 3274 3183 3277 3233
rect 3290 3213 3309 3216
rect 3282 3153 3285 3206
rect 3290 3203 3293 3213
rect 3298 3163 3301 3206
rect 3314 3166 3317 3233
rect 3322 3203 3325 3266
rect 3338 3196 3341 3273
rect 3354 3263 3357 3443
rect 3362 3413 3365 3426
rect 3374 3396 3377 3583
rect 3374 3393 3381 3396
rect 3378 3373 3381 3393
rect 3354 3206 3357 3226
rect 3330 3193 3341 3196
rect 3350 3203 3357 3206
rect 3314 3163 3321 3166
rect 3282 2993 3285 3136
rect 3306 3123 3309 3156
rect 3318 3116 3321 3163
rect 3314 3113 3321 3116
rect 3314 3026 3317 3113
rect 3314 3023 3321 3026
rect 3306 3003 3309 3016
rect 3266 2983 3277 2986
rect 3254 2963 3261 2966
rect 3258 2856 3261 2963
rect 3250 2853 3261 2856
rect 3250 2833 3253 2853
rect 3250 2813 3253 2826
rect 3258 2793 3261 2806
rect 3226 2763 3233 2766
rect 3226 2743 3229 2763
rect 3266 2746 3269 2816
rect 3274 2803 3277 2983
rect 3306 2903 3309 2976
rect 3318 2966 3321 3023
rect 3330 2973 3333 3193
rect 3350 3116 3353 3203
rect 3362 3123 3365 3206
rect 3378 3196 3381 3316
rect 3386 3293 3389 3736
rect 3394 3306 3397 3813
rect 3402 3463 3405 3796
rect 3426 3766 3429 3873
rect 3426 3763 3437 3766
rect 3410 3713 3413 3726
rect 3410 3596 3413 3626
rect 3418 3603 3421 3716
rect 3434 3623 3437 3763
rect 3450 3743 3453 3966
rect 3474 3843 3477 4003
rect 3490 3963 3493 4013
rect 3510 3956 3513 4123
rect 3522 3966 3525 4116
rect 3534 4066 3537 4163
rect 3534 4063 3541 4066
rect 3522 3963 3529 3966
rect 3510 3953 3517 3956
rect 3490 3933 3493 3946
rect 3498 3933 3509 3936
rect 3514 3926 3517 3953
rect 3458 3803 3461 3826
rect 3482 3823 3485 3926
rect 3498 3906 3501 3926
rect 3494 3903 3501 3906
rect 3506 3923 3517 3926
rect 3466 3783 3469 3816
rect 3494 3806 3497 3903
rect 3482 3803 3497 3806
rect 3458 3676 3461 3726
rect 3442 3673 3461 3676
rect 3426 3603 3429 3616
rect 3434 3603 3437 3616
rect 3442 3603 3445 3673
rect 3466 3666 3469 3766
rect 3458 3663 3469 3666
rect 3410 3593 3429 3596
rect 3458 3593 3461 3663
rect 3474 3646 3477 3746
rect 3470 3643 3477 3646
rect 3410 3533 3413 3556
rect 3426 3476 3429 3593
rect 3470 3556 3473 3643
rect 3482 3593 3485 3803
rect 3506 3786 3509 3923
rect 3526 3916 3529 3963
rect 3538 3923 3541 4063
rect 3522 3913 3529 3916
rect 3522 3826 3525 3913
rect 3522 3823 3529 3826
rect 3502 3783 3509 3786
rect 3502 3636 3505 3783
rect 3514 3733 3517 3816
rect 3526 3746 3529 3823
rect 3522 3743 3529 3746
rect 3502 3633 3509 3636
rect 3498 3603 3501 3616
rect 3470 3553 3477 3556
rect 3466 3523 3469 3536
rect 3410 3473 3429 3476
rect 3410 3403 3413 3473
rect 3434 3446 3437 3466
rect 3474 3446 3477 3553
rect 3506 3536 3509 3633
rect 3514 3603 3517 3726
rect 3498 3533 3509 3536
rect 3498 3446 3501 3533
rect 3514 3513 3517 3526
rect 3522 3506 3525 3743
rect 3530 3713 3533 3726
rect 3538 3706 3541 3846
rect 3546 3776 3549 4186
rect 3562 4176 3565 4253
rect 3554 4173 3565 4176
rect 3554 3976 3557 4173
rect 3562 4103 3565 4156
rect 3570 4113 3573 4126
rect 3586 4103 3589 4276
rect 3594 4213 3597 4293
rect 3602 4206 3605 4336
rect 3594 4203 3605 4206
rect 3610 4203 3613 4346
rect 3642 4333 3645 4356
rect 3694 4353 3701 4356
rect 3618 4213 3621 4326
rect 3626 4243 3629 4326
rect 3634 4196 3637 4216
rect 3618 4193 3637 4196
rect 3594 4093 3597 4126
rect 3602 4113 3605 4156
rect 3618 4133 3621 4193
rect 3626 4113 3629 4126
rect 3562 3993 3565 4016
rect 3586 3983 3589 4056
rect 3554 3973 3565 3976
rect 3562 3796 3565 3973
rect 3578 3933 3581 3966
rect 3602 3963 3605 4006
rect 3634 4003 3637 4186
rect 3642 4133 3645 4226
rect 3650 4203 3653 4286
rect 3658 4223 3661 4336
rect 3666 4213 3669 4326
rect 3674 4306 3677 4336
rect 3694 4306 3697 4353
rect 3674 4303 3685 4306
rect 3694 4303 3701 4306
rect 3682 4216 3685 4303
rect 3674 4213 3685 4216
rect 3674 4193 3677 4213
rect 3650 4123 3653 4136
rect 3642 4013 3645 4036
rect 3650 3993 3653 4006
rect 3658 3986 3661 4106
rect 3666 4073 3669 4136
rect 3674 4003 3677 4016
rect 3690 4003 3693 4166
rect 3698 4133 3701 4303
rect 3714 4203 3717 4513
rect 3762 4506 3765 4523
rect 3722 4413 3725 4426
rect 3738 4413 3741 4476
rect 3754 4413 3757 4506
rect 3762 4503 3773 4506
rect 3770 4426 3773 4503
rect 3762 4423 3773 4426
rect 3730 4393 3733 4406
rect 3762 4403 3765 4423
rect 3762 4323 3765 4346
rect 3730 4213 3733 4226
rect 3714 4123 3717 4136
rect 3738 4086 3741 4266
rect 3786 4236 3789 4586
rect 3794 4516 3797 4536
rect 3810 4533 3813 4586
rect 3842 4583 3845 4616
rect 3826 4533 3829 4576
rect 3818 4523 3837 4526
rect 3850 4516 3853 4536
rect 3898 4533 3901 4616
rect 3794 4513 3805 4516
rect 3802 4446 3805 4513
rect 3846 4513 3853 4516
rect 3794 4443 3805 4446
rect 3794 4413 3797 4443
rect 3802 4406 3805 4426
rect 3802 4403 3813 4406
rect 3810 4286 3813 4403
rect 3802 4283 3813 4286
rect 3802 4246 3805 4283
rect 3834 4266 3837 4466
rect 3846 4426 3849 4513
rect 3858 4506 3861 4526
rect 3922 4523 3925 4536
rect 3930 4523 3933 4616
rect 3938 4533 3941 4606
rect 3954 4533 3957 4616
rect 4002 4603 4005 4616
rect 4050 4593 4053 4606
rect 3858 4503 3869 4506
rect 3866 4456 3869 4503
rect 3962 4493 3965 4536
rect 3858 4453 3869 4456
rect 3846 4423 3853 4426
rect 3850 4316 3853 4423
rect 3858 4403 3861 4453
rect 3866 4413 3869 4436
rect 3882 4413 3885 4426
rect 3906 4366 3909 4426
rect 3922 4403 3925 4426
rect 3938 4373 3941 4436
rect 3946 4423 3949 4436
rect 3986 4426 3989 4526
rect 3946 4383 3949 4416
rect 3962 4413 3965 4426
rect 3978 4423 3989 4426
rect 3978 4376 3981 4423
rect 3978 4373 3989 4376
rect 3882 4333 3885 4346
rect 3826 4263 3837 4266
rect 3846 4313 3853 4316
rect 3858 4323 3877 4326
rect 3890 4323 3893 4366
rect 3906 4363 3913 4366
rect 3802 4243 3813 4246
rect 3786 4233 3797 4236
rect 3770 4133 3773 4166
rect 3778 4103 3781 4206
rect 3786 4113 3789 4126
rect 3794 4123 3797 4233
rect 3810 4156 3813 4243
rect 3826 4193 3829 4263
rect 3846 4236 3849 4313
rect 3846 4233 3853 4236
rect 3834 4203 3837 4226
rect 3802 4153 3813 4156
rect 3842 4153 3845 4216
rect 3730 4083 3741 4086
rect 3658 3983 3669 3986
rect 3618 3946 3621 3966
rect 3594 3933 3597 3946
rect 3618 3943 3629 3946
rect 3602 3933 3613 3936
rect 3586 3813 3589 3926
rect 3602 3883 3605 3926
rect 3610 3803 3613 3926
rect 3626 3836 3629 3943
rect 3650 3923 3653 3946
rect 3666 3916 3669 3983
rect 3658 3913 3669 3916
rect 3618 3833 3629 3836
rect 3562 3793 3573 3796
rect 3546 3773 3557 3776
rect 3530 3703 3541 3706
rect 3530 3533 3533 3703
rect 3554 3696 3557 3773
rect 3546 3693 3557 3696
rect 3546 3636 3549 3693
rect 3542 3633 3549 3636
rect 3542 3586 3545 3633
rect 3570 3626 3573 3793
rect 3618 3786 3621 3833
rect 3610 3783 3621 3786
rect 3610 3706 3613 3783
rect 3626 3713 3629 3816
rect 3634 3733 3637 3806
rect 3642 3713 3645 3886
rect 3658 3883 3661 3913
rect 3650 3763 3653 3806
rect 3610 3703 3629 3706
rect 3626 3636 3629 3703
rect 3554 3623 3573 3626
rect 3618 3633 3629 3636
rect 3554 3603 3557 3623
rect 3542 3583 3549 3586
rect 3546 3563 3549 3583
rect 3538 3533 3549 3536
rect 3530 3523 3541 3526
rect 3554 3506 3557 3596
rect 3570 3546 3573 3566
rect 3562 3533 3565 3546
rect 3570 3543 3581 3546
rect 3434 3443 3445 3446
rect 3474 3443 3485 3446
rect 3498 3443 3509 3446
rect 3442 3396 3445 3443
rect 3458 3403 3461 3416
rect 3434 3393 3445 3396
rect 3418 3356 3421 3376
rect 3418 3353 3425 3356
rect 3402 3313 3405 3326
rect 3394 3303 3405 3306
rect 3410 3303 3413 3336
rect 3402 3296 3405 3303
rect 3402 3293 3413 3296
rect 3386 3233 3397 3236
rect 3402 3213 3405 3246
rect 3410 3223 3413 3293
rect 3422 3216 3425 3353
rect 3418 3213 3425 3216
rect 3378 3193 3389 3196
rect 3350 3113 3357 3116
rect 3314 2963 3321 2966
rect 3242 2743 3261 2746
rect 3266 2743 3277 2746
rect 3242 2736 3245 2743
rect 3234 2733 3245 2736
rect 3226 2663 3229 2726
rect 3234 2686 3237 2716
rect 3242 2703 3245 2726
rect 3234 2683 3241 2686
rect 3238 2596 3241 2683
rect 3250 2613 3253 2736
rect 3258 2613 3261 2743
rect 3266 2723 3269 2736
rect 3274 2723 3277 2743
rect 3282 2636 3285 2786
rect 3290 2706 3293 2806
rect 3298 2733 3301 2746
rect 3290 2703 3301 2706
rect 3278 2633 3285 2636
rect 3238 2593 3245 2596
rect 3194 2583 3205 2586
rect 3202 2566 3205 2583
rect 3202 2563 3209 2566
rect 3194 2413 3197 2536
rect 3206 2406 3209 2563
rect 3178 2363 3189 2366
rect 3202 2403 3209 2406
rect 3130 2303 3141 2306
rect 3138 2226 3141 2303
rect 3106 2223 3117 2226
rect 3138 2223 3149 2226
rect 3082 2213 3093 2216
rect 3082 2173 3085 2206
rect 3090 2146 3093 2213
rect 3114 2176 3117 2223
rect 3146 2203 3149 2223
rect 3154 2203 3157 2326
rect 3178 2323 3181 2363
rect 3186 2333 3189 2346
rect 3162 2213 3165 2226
rect 3170 2216 3173 2306
rect 3186 2273 3189 2326
rect 3202 2313 3205 2403
rect 3218 2343 3221 2566
rect 3226 2556 3229 2576
rect 3226 2553 3233 2556
rect 3230 2456 3233 2553
rect 3226 2453 3233 2456
rect 3226 2353 3229 2453
rect 3242 2436 3245 2593
rect 3278 2566 3281 2633
rect 3290 2613 3293 2626
rect 3298 2603 3301 2703
rect 3314 2596 3317 2963
rect 3322 2783 3325 2906
rect 3330 2893 3333 2936
rect 3322 2603 3325 2626
rect 3274 2563 3281 2566
rect 3290 2593 3317 2596
rect 3234 2433 3245 2436
rect 3234 2326 3237 2433
rect 3226 2323 3237 2326
rect 3242 2323 3245 2416
rect 3170 2213 3181 2216
rect 3186 2213 3189 2226
rect 3210 2216 3213 2276
rect 3194 2213 3213 2216
rect 3074 2143 3093 2146
rect 3106 2173 3117 2176
rect 3058 2123 3061 2136
rect 3074 2096 3077 2143
rect 3106 2133 3109 2173
rect 3130 2113 3133 2156
rect 3170 2123 3173 2206
rect 3178 2203 3189 2206
rect 3194 2166 3197 2213
rect 3194 2163 3201 2166
rect 3074 2093 3085 2096
rect 3082 2026 3085 2093
rect 3082 2023 3089 2026
rect 3026 1993 3029 2006
rect 3042 1973 3045 2006
rect 3066 2003 3069 2016
rect 3010 1923 3013 1936
rect 3042 1933 3045 1946
rect 3050 1923 3053 1966
rect 3074 1933 3077 2016
rect 3086 1966 3089 2023
rect 3106 1993 3109 2016
rect 3086 1963 3093 1966
rect 3090 1916 3093 1963
rect 2906 1823 2917 1826
rect 2802 1803 2821 1806
rect 2874 1786 2877 1806
rect 2882 1803 2885 1816
rect 2866 1783 2877 1786
rect 2786 1623 2789 1636
rect 2802 1613 2805 1726
rect 2810 1716 2813 1776
rect 2866 1733 2869 1783
rect 2810 1713 2821 1716
rect 2818 1606 2821 1713
rect 2842 1633 2845 1726
rect 2810 1603 2821 1606
rect 2754 1513 2757 1526
rect 2682 1333 2693 1336
rect 2738 1333 2741 1396
rect 2762 1376 2765 1416
rect 2778 1413 2781 1536
rect 2794 1513 2797 1526
rect 2802 1426 2805 1516
rect 2810 1503 2813 1603
rect 2850 1526 2853 1616
rect 2866 1603 2869 1726
rect 2922 1723 2925 1806
rect 2930 1713 2933 1826
rect 2970 1803 2973 1826
rect 2994 1773 2997 1826
rect 2938 1743 2941 1756
rect 2954 1716 2957 1736
rect 3002 1733 3005 1806
rect 3034 1773 3037 1876
rect 3074 1873 3077 1916
rect 3082 1913 3093 1916
rect 3082 1893 3085 1913
rect 3066 1823 3077 1826
rect 3066 1813 3069 1823
rect 3106 1786 3109 1986
rect 3138 1923 3141 1996
rect 3154 1986 3157 2006
rect 3170 1986 3173 2116
rect 3198 2106 3201 2163
rect 3210 2123 3213 2206
rect 3226 2156 3229 2323
rect 3242 2296 3245 2316
rect 3238 2293 3245 2296
rect 3238 2176 3241 2293
rect 3238 2173 3245 2176
rect 3226 2153 3237 2156
rect 3234 2133 3237 2153
rect 3154 1983 3173 1986
rect 3194 2103 3201 2106
rect 3194 1976 3197 2103
rect 3218 2056 3221 2126
rect 3242 2116 3245 2173
rect 3238 2113 3245 2116
rect 3146 1913 3149 1976
rect 3186 1973 3197 1976
rect 3210 2053 3221 2056
rect 3122 1903 3133 1906
rect 3130 1833 3133 1886
rect 3138 1813 3141 1906
rect 3186 1896 3189 1973
rect 3210 1946 3213 2053
rect 3210 1943 3221 1946
rect 3194 1903 3197 1926
rect 3202 1913 3205 1926
rect 3218 1923 3221 1943
rect 3210 1903 3213 1916
rect 3146 1823 3149 1896
rect 3186 1893 3205 1896
rect 3106 1783 3113 1786
rect 2946 1713 2957 1716
rect 2962 1713 2965 1726
rect 2946 1656 2949 1713
rect 2970 1696 2973 1726
rect 3018 1716 3021 1736
rect 2962 1693 2973 1696
rect 3010 1713 3021 1716
rect 2946 1653 2957 1656
rect 2906 1623 2925 1626
rect 2866 1533 2869 1546
rect 2842 1523 2869 1526
rect 2882 1503 2885 1606
rect 2906 1603 2909 1623
rect 2938 1613 2941 1636
rect 2954 1633 2957 1653
rect 2962 1626 2965 1693
rect 3010 1636 3013 1713
rect 3010 1633 3021 1636
rect 2954 1623 2965 1626
rect 2954 1613 2957 1623
rect 3010 1593 3013 1616
rect 3018 1583 3021 1633
rect 3034 1613 3037 1756
rect 3058 1633 3061 1726
rect 3066 1723 3069 1736
rect 3074 1716 3077 1736
rect 3066 1713 3077 1716
rect 3074 1693 3077 1713
rect 2914 1523 2917 1536
rect 2922 1533 2933 1536
rect 2914 1503 2917 1516
rect 2922 1513 2925 1526
rect 2786 1413 2789 1426
rect 2794 1423 2805 1426
rect 2786 1393 2789 1406
rect 2746 1333 2749 1356
rect 2682 1323 2685 1333
rect 2690 1313 2693 1326
rect 2674 1253 2685 1256
rect 2634 1213 2637 1226
rect 2642 1163 2645 1216
rect 2666 1156 2669 1176
rect 2658 1153 2669 1156
rect 2610 1083 2613 1126
rect 2626 1106 2629 1126
rect 2634 1116 2637 1136
rect 2634 1113 2645 1116
rect 2622 1103 2629 1106
rect 2554 1013 2557 1043
rect 2622 1036 2625 1103
rect 2642 1066 2645 1113
rect 2634 1063 2645 1066
rect 2658 1066 2661 1153
rect 2682 1146 2685 1253
rect 2674 1143 2685 1146
rect 2658 1063 2665 1066
rect 2622 1033 2629 1036
rect 2482 903 2485 926
rect 2410 763 2421 766
rect 2378 733 2389 736
rect 2274 653 2285 656
rect 2242 643 2253 646
rect 2250 596 2253 643
rect 2266 613 2269 626
rect 2242 593 2253 596
rect 2194 573 2205 576
rect 2138 563 2149 566
rect 2130 513 2133 526
rect 2146 506 2149 563
rect 2202 556 2205 573
rect 2138 503 2149 506
rect 2130 413 2133 426
rect 2138 393 2141 503
rect 2178 403 2181 556
rect 2202 553 2213 556
rect 2210 506 2213 553
rect 2202 503 2213 506
rect 2202 436 2205 503
rect 2198 433 2205 436
rect 2114 363 2121 366
rect 2098 213 2101 326
rect 2118 306 2121 363
rect 2138 333 2141 346
rect 2178 336 2181 396
rect 2198 386 2201 433
rect 2242 426 2245 593
rect 2282 566 2285 653
rect 2274 563 2285 566
rect 2274 466 2277 563
rect 2274 463 2285 466
rect 2282 446 2285 463
rect 2282 443 2289 446
rect 2242 423 2253 426
rect 2198 383 2205 386
rect 2202 366 2205 383
rect 2202 363 2209 366
rect 2178 333 2185 336
rect 2118 303 2133 306
rect 2130 246 2133 303
rect 2170 286 2173 326
rect 2162 283 2173 286
rect 2130 243 2141 246
rect 2082 193 2089 196
rect 2122 193 2125 206
rect 2082 173 2085 193
rect 2138 186 2141 243
rect 2146 213 2149 266
rect 2122 183 2141 186
rect 2122 166 2125 183
rect 2118 163 2125 166
rect 2098 133 2101 146
rect 2118 106 2121 163
rect 2162 156 2165 283
rect 2182 276 2185 333
rect 2206 286 2209 363
rect 2218 343 2221 406
rect 2242 356 2245 416
rect 2250 373 2253 423
rect 2286 376 2289 443
rect 2298 413 2301 696
rect 2362 693 2373 696
rect 2362 636 2365 693
rect 2386 686 2389 733
rect 2402 713 2405 736
rect 2418 733 2421 763
rect 2434 743 2437 836
rect 2442 833 2453 836
rect 2490 833 2493 926
rect 2506 913 2509 936
rect 2522 883 2525 986
rect 2538 906 2541 926
rect 2546 906 2549 926
rect 2554 923 2557 1006
rect 2562 923 2565 1026
rect 2602 1013 2605 1026
rect 2626 1013 2629 1033
rect 2570 993 2573 1006
rect 2618 1003 2629 1006
rect 2634 996 2637 1063
rect 2618 993 2637 996
rect 2578 916 2581 976
rect 2538 903 2549 906
rect 2546 846 2549 903
rect 2570 913 2581 916
rect 2610 913 2613 926
rect 2546 843 2557 846
rect 2442 803 2445 833
rect 2434 723 2437 736
rect 2450 733 2453 796
rect 2382 683 2389 686
rect 2362 633 2373 636
rect 2306 603 2309 626
rect 2314 533 2317 616
rect 2338 523 2341 626
rect 2362 536 2365 546
rect 2346 533 2365 536
rect 2370 516 2373 633
rect 2382 576 2385 683
rect 2362 513 2373 516
rect 2378 573 2385 576
rect 2306 383 2309 396
rect 2314 393 2317 406
rect 2282 373 2289 376
rect 2226 353 2245 356
rect 2218 323 2221 336
rect 2178 273 2185 276
rect 2202 283 2209 286
rect 2178 256 2181 273
rect 2174 253 2181 256
rect 2174 176 2177 253
rect 2202 226 2205 283
rect 2226 246 2229 353
rect 2198 223 2205 226
rect 2218 243 2229 246
rect 2198 176 2201 223
rect 2174 173 2181 176
rect 2198 173 2205 176
rect 2162 153 2173 156
rect 2138 133 2141 146
rect 2066 93 2077 96
rect 2030 83 2037 86
rect 2018 0 2021 36
rect 2034 0 2037 83
rect 2058 0 2061 16
rect 2074 0 2077 93
rect 2090 0 2093 86
rect 2106 0 2109 106
rect 2118 103 2125 106
rect 2122 0 2125 103
rect 2138 0 2141 116
rect 2162 113 2165 126
rect 2154 0 2157 96
rect 2170 76 2173 153
rect 2178 93 2181 173
rect 2202 83 2205 173
rect 2170 73 2181 76
rect 2178 16 2181 73
rect 2170 13 2181 16
rect 2170 0 2173 13
rect 2210 0 2213 216
rect 2218 176 2221 243
rect 2250 236 2253 346
rect 2282 283 2285 373
rect 2314 356 2317 376
rect 2314 353 2321 356
rect 2242 233 2253 236
rect 2218 173 2237 176
rect 2218 123 2221 166
rect 2234 0 2237 173
rect 2242 143 2245 233
rect 2258 133 2261 146
rect 2274 143 2277 206
rect 2298 186 2301 326
rect 2294 183 2301 186
rect 2250 0 2253 106
rect 2282 103 2285 126
rect 2294 116 2297 183
rect 2294 113 2301 116
rect 2274 0 2277 96
rect 2298 93 2301 113
rect 2306 33 2309 286
rect 2318 246 2321 353
rect 2330 323 2333 446
rect 2362 426 2365 513
rect 2378 496 2381 573
rect 2394 556 2397 616
rect 2410 613 2437 616
rect 2410 603 2413 613
rect 2418 593 2421 606
rect 2466 593 2469 746
rect 2482 713 2485 726
rect 2506 636 2509 806
rect 2538 776 2541 816
rect 2554 783 2557 843
rect 2570 803 2573 913
rect 2618 896 2621 993
rect 2642 973 2645 1046
rect 2662 976 2665 1063
rect 2662 973 2669 976
rect 2650 946 2653 966
rect 2646 943 2653 946
rect 2666 946 2669 973
rect 2674 963 2677 1143
rect 2698 1123 2701 1306
rect 2754 1303 2757 1376
rect 2762 1373 2773 1376
rect 2770 1296 2773 1373
rect 2794 1303 2797 1423
rect 2810 1363 2813 1416
rect 2890 1343 2893 1356
rect 2898 1343 2901 1396
rect 2906 1336 2909 1366
rect 2898 1333 2909 1336
rect 2914 1326 2917 1446
rect 2930 1413 2933 1533
rect 3026 1526 3029 1546
rect 3034 1533 3045 1536
rect 3050 1533 3053 1626
rect 3074 1606 3077 1636
rect 3082 1613 3085 1726
rect 3090 1703 3093 1726
rect 3098 1643 3101 1756
rect 3110 1656 3113 1783
rect 3122 1713 3125 1726
rect 3138 1703 3141 1716
rect 3146 1703 3149 1716
rect 3154 1686 3157 1816
rect 3106 1653 3113 1656
rect 3146 1683 3157 1686
rect 3090 1623 3093 1636
rect 3058 1603 3077 1606
rect 2938 1496 2941 1526
rect 3026 1523 3037 1526
rect 2938 1493 2949 1496
rect 2946 1406 2949 1493
rect 2938 1403 2949 1406
rect 2938 1383 2941 1403
rect 2762 1293 2773 1296
rect 2722 1136 2725 1216
rect 2738 1213 2741 1226
rect 2762 1213 2765 1293
rect 2802 1223 2805 1326
rect 2906 1323 2917 1326
rect 2930 1323 2933 1346
rect 2962 1333 2965 1466
rect 3018 1436 3021 1506
rect 3018 1433 3025 1436
rect 2802 1193 2805 1216
rect 2826 1203 2829 1216
rect 2842 1213 2845 1306
rect 2842 1193 2845 1206
rect 2850 1196 2853 1226
rect 2850 1193 2861 1196
rect 2706 1133 2725 1136
rect 2738 1133 2741 1146
rect 2850 1143 2853 1166
rect 2858 1133 2861 1193
rect 2866 1156 2869 1236
rect 2906 1233 2909 1323
rect 2874 1203 2877 1216
rect 2970 1203 2973 1386
rect 2978 1333 2981 1346
rect 2994 1343 2997 1396
rect 3002 1323 3005 1356
rect 3010 1333 3013 1426
rect 3022 1366 3025 1433
rect 3018 1363 3025 1366
rect 3010 1223 3013 1236
rect 3018 1206 3021 1363
rect 3034 1333 3037 1523
rect 3042 1503 3045 1526
rect 3042 1403 3045 1426
rect 3050 1423 3053 1436
rect 3058 1433 3061 1576
rect 3042 1343 3053 1346
rect 3050 1233 3053 1326
rect 3058 1323 3061 1416
rect 2978 1196 2981 1206
rect 2962 1193 2981 1196
rect 2866 1153 2877 1156
rect 2682 1013 2685 1046
rect 2706 986 2709 1133
rect 2754 1113 2757 1126
rect 2762 1033 2765 1126
rect 2722 993 2725 1006
rect 2666 943 2677 946
rect 2578 813 2581 826
rect 2586 813 2589 896
rect 2614 893 2621 896
rect 2614 826 2617 893
rect 2626 833 2629 926
rect 2634 903 2637 926
rect 2646 826 2649 943
rect 2674 886 2677 943
rect 2690 923 2693 986
rect 2706 983 2717 986
rect 2730 983 2733 1016
rect 2746 1013 2749 1026
rect 2714 906 2717 983
rect 2730 923 2733 936
rect 2754 933 2757 1016
rect 2850 1003 2853 1036
rect 2842 973 2845 996
rect 2858 956 2861 1056
rect 2866 1043 2869 1146
rect 2874 1053 2877 1153
rect 2986 1143 2989 1156
rect 2882 1113 2885 1136
rect 2994 1133 2997 1206
rect 3010 1203 3021 1206
rect 3002 1133 3005 1166
rect 3010 1126 3013 1203
rect 3018 1133 3021 1156
rect 3026 1136 3029 1226
rect 3034 1213 3061 1216
rect 3066 1146 3069 1596
rect 3098 1583 3101 1596
rect 3106 1573 3109 1653
rect 3114 1613 3117 1636
rect 3122 1603 3125 1636
rect 3130 1623 3133 1646
rect 3146 1606 3149 1683
rect 3162 1613 3165 1716
rect 3170 1703 3173 1726
rect 3178 1713 3181 1816
rect 3202 1753 3205 1893
rect 3226 1826 3229 2106
rect 3238 1966 3241 2113
rect 3238 1963 3245 1966
rect 3242 1943 3245 1963
rect 3234 1926 3237 1936
rect 3234 1923 3245 1926
rect 3250 1906 3253 2396
rect 3258 2346 3261 2526
rect 3274 2466 3277 2563
rect 3274 2463 3285 2466
rect 3266 2363 3269 2446
rect 3274 2403 3277 2416
rect 3282 2396 3285 2463
rect 3290 2423 3293 2593
rect 3330 2586 3333 2826
rect 3338 2803 3341 2816
rect 3354 2766 3357 3113
rect 3370 3046 3373 3116
rect 3366 3043 3373 3046
rect 3366 2976 3369 3043
rect 3386 3036 3389 3193
rect 3410 3123 3413 3156
rect 3418 3113 3421 3213
rect 3434 3106 3437 3393
rect 3458 3333 3469 3336
rect 3442 3303 3445 3316
rect 3450 3236 3453 3326
rect 3466 3313 3469 3326
rect 3474 3306 3477 3436
rect 3482 3363 3485 3443
rect 3482 3333 3485 3356
rect 3446 3233 3453 3236
rect 3466 3303 3477 3306
rect 3466 3233 3469 3303
rect 3482 3276 3485 3326
rect 3490 3323 3493 3426
rect 3498 3333 3501 3416
rect 3506 3316 3509 3443
rect 3514 3403 3517 3506
rect 3522 3503 3529 3506
rect 3526 3386 3529 3503
rect 3550 3503 3557 3506
rect 3550 3436 3553 3503
rect 3578 3496 3581 3543
rect 3570 3493 3581 3496
rect 3550 3433 3557 3436
rect 3538 3413 3541 3426
rect 3554 3413 3557 3433
rect 3538 3403 3549 3406
rect 3562 3403 3565 3486
rect 3526 3383 3533 3386
rect 3502 3313 3509 3316
rect 3482 3273 3493 3276
rect 3446 3126 3449 3233
rect 3446 3123 3453 3126
rect 3402 3083 3405 3106
rect 3418 3103 3437 3106
rect 3378 3033 3389 3036
rect 3418 3036 3421 3103
rect 3418 3033 3425 3036
rect 3366 2973 3373 2976
rect 3346 2763 3357 2766
rect 3346 2686 3349 2763
rect 3362 2723 3365 2956
rect 3370 2876 3373 2973
rect 3378 2953 3381 3033
rect 3386 3013 3397 3016
rect 3410 2996 3413 3026
rect 3402 2993 3413 2996
rect 3378 2923 3381 2946
rect 3370 2873 3381 2876
rect 3378 2816 3381 2873
rect 3402 2836 3405 2993
rect 3422 2986 3425 3033
rect 3418 2983 3425 2986
rect 3402 2833 3413 2836
rect 3370 2813 3381 2816
rect 3370 2706 3373 2813
rect 3366 2703 3373 2706
rect 3346 2683 3357 2686
rect 3326 2583 3333 2586
rect 3314 2533 3317 2546
rect 3290 2403 3293 2416
rect 3282 2393 3293 2396
rect 3298 2393 3301 2426
rect 3258 2343 3269 2346
rect 3266 2276 3269 2343
rect 3290 2336 3293 2393
rect 3290 2333 3297 2336
rect 3258 2273 3269 2276
rect 3258 2133 3261 2273
rect 3258 2103 3261 2116
rect 3274 2103 3277 2256
rect 3282 2203 3285 2326
rect 3294 2196 3297 2333
rect 3306 2273 3309 2516
rect 3326 2496 3329 2583
rect 3338 2543 3341 2616
rect 3346 2613 3349 2666
rect 3354 2596 3357 2683
rect 3366 2626 3369 2703
rect 3362 2623 3369 2626
rect 3362 2603 3365 2623
rect 3378 2613 3381 2796
rect 3350 2593 3357 2596
rect 3350 2526 3353 2593
rect 3346 2523 3353 2526
rect 3338 2503 3341 2516
rect 3346 2506 3349 2523
rect 3362 2516 3365 2596
rect 3354 2513 3365 2516
rect 3378 2506 3381 2606
rect 3386 2603 3389 2616
rect 3394 2533 3397 2616
rect 3402 2603 3405 2816
rect 3410 2683 3413 2833
rect 3418 2776 3421 2983
rect 3434 2963 3437 3036
rect 3442 3013 3445 3106
rect 3450 3076 3453 3123
rect 3458 3093 3461 3226
rect 3466 3206 3469 3226
rect 3482 3223 3485 3266
rect 3466 3203 3477 3206
rect 3474 3086 3477 3203
rect 3466 3083 3477 3086
rect 3450 3073 3457 3076
rect 3454 3006 3457 3073
rect 3466 3023 3469 3083
rect 3490 3053 3493 3273
rect 3502 3246 3505 3313
rect 3502 3243 3509 3246
rect 3506 3223 3509 3243
rect 3514 3216 3517 3376
rect 3530 3256 3533 3383
rect 3570 3373 3573 3493
rect 3594 3486 3597 3606
rect 3618 3556 3621 3633
rect 3618 3553 3629 3556
rect 3602 3513 3605 3536
rect 3618 3513 3621 3526
rect 3594 3483 3605 3486
rect 3578 3403 3581 3476
rect 3602 3396 3605 3483
rect 3626 3473 3629 3553
rect 3642 3446 3645 3576
rect 3650 3566 3653 3756
rect 3698 3753 3701 3986
rect 3714 3933 3717 3956
rect 3666 3723 3669 3736
rect 3714 3733 3717 3756
rect 3698 3576 3701 3616
rect 3698 3573 3709 3576
rect 3650 3563 3669 3566
rect 3594 3393 3605 3396
rect 3634 3443 3645 3446
rect 3506 3213 3517 3216
rect 3522 3253 3533 3256
rect 3506 3046 3509 3213
rect 3522 3163 3525 3253
rect 3538 3213 3541 3236
rect 3546 3223 3549 3296
rect 3546 3146 3549 3216
rect 3538 3143 3549 3146
rect 3514 3113 3517 3136
rect 3538 3126 3541 3143
rect 3522 3123 3541 3126
rect 3506 3043 3513 3046
rect 3450 3003 3457 3006
rect 3442 2916 3445 2936
rect 3434 2913 3445 2916
rect 3434 2836 3437 2913
rect 3434 2833 3445 2836
rect 3426 2793 3429 2816
rect 3442 2813 3445 2833
rect 3450 2826 3453 3003
rect 3466 2933 3469 2956
rect 3482 2946 3485 3006
rect 3510 2976 3513 3043
rect 3506 2973 3513 2976
rect 3506 2953 3509 2973
rect 3474 2943 3485 2946
rect 3450 2823 3461 2826
rect 3418 2773 3425 2776
rect 3422 2676 3425 2773
rect 3418 2673 3425 2676
rect 3418 2593 3421 2673
rect 3346 2503 3357 2506
rect 3326 2493 3333 2496
rect 3314 2433 3325 2436
rect 3290 2193 3297 2196
rect 3290 2113 3293 2193
rect 3282 2033 3285 2046
rect 3242 1903 3253 1906
rect 3242 1846 3245 1903
rect 3242 1843 3253 1846
rect 3226 1823 3237 1826
rect 3170 1623 3173 1636
rect 3146 1603 3157 1606
rect 3098 1533 3101 1546
rect 3146 1533 3149 1546
rect 3074 1386 3077 1526
rect 3082 1403 3085 1446
rect 3090 1423 3093 1436
rect 3130 1413 3133 1426
rect 3138 1406 3141 1516
rect 3114 1393 3117 1406
rect 3074 1383 3085 1386
rect 3082 1176 3085 1383
rect 3098 1193 3101 1336
rect 3122 1333 3125 1346
rect 3122 1313 3125 1326
rect 3130 1226 3133 1406
rect 3138 1403 3145 1406
rect 3142 1336 3145 1403
rect 3138 1333 3145 1336
rect 3138 1313 3141 1333
rect 3130 1223 3141 1226
rect 3026 1133 3037 1136
rect 3042 1133 3045 1146
rect 3058 1143 3069 1146
rect 3074 1173 3085 1176
rect 2866 1003 2869 1036
rect 2898 1033 2901 1126
rect 3010 1123 3021 1126
rect 2874 983 2877 996
rect 2858 953 2877 956
rect 2850 943 2869 946
rect 2850 933 2861 936
rect 2866 933 2869 943
rect 2874 926 2877 953
rect 2714 903 2725 906
rect 2658 883 2677 886
rect 2614 823 2621 826
rect 2530 773 2541 776
rect 2530 666 2533 773
rect 2546 733 2549 746
rect 2530 663 2541 666
rect 2498 633 2509 636
rect 2386 553 2397 556
rect 2386 523 2389 553
rect 2498 546 2501 633
rect 2530 626 2533 646
rect 2538 636 2541 663
rect 2554 643 2557 736
rect 2562 706 2565 726
rect 2578 723 2581 736
rect 2586 733 2589 806
rect 2602 743 2605 816
rect 2610 786 2613 806
rect 2618 786 2621 823
rect 2626 813 2629 826
rect 2646 823 2653 826
rect 2634 803 2645 806
rect 2610 783 2621 786
rect 2618 736 2621 783
rect 2562 703 2573 706
rect 2570 646 2573 703
rect 2562 643 2573 646
rect 2538 633 2557 636
rect 2514 603 2517 616
rect 2522 593 2525 626
rect 2530 623 2541 626
rect 2538 613 2541 623
rect 2546 613 2549 626
rect 2554 616 2557 633
rect 2562 623 2565 643
rect 2554 613 2565 616
rect 2530 593 2533 606
rect 2538 603 2557 606
rect 2498 543 2509 546
rect 2442 513 2445 536
rect 2378 493 2389 496
rect 2386 426 2389 493
rect 2354 423 2365 426
rect 2378 423 2389 426
rect 2354 413 2357 423
rect 2338 383 2341 406
rect 2354 323 2357 396
rect 2370 376 2373 416
rect 2378 403 2381 423
rect 2366 373 2373 376
rect 2366 286 2369 373
rect 2434 333 2437 346
rect 2458 343 2461 536
rect 2498 506 2501 526
rect 2490 503 2501 506
rect 2490 436 2493 503
rect 2490 433 2501 436
rect 2498 416 2501 433
rect 2410 313 2413 326
rect 2466 316 2469 336
rect 2474 323 2477 416
rect 2482 413 2501 416
rect 2482 403 2485 413
rect 2506 346 2509 543
rect 2538 523 2541 603
rect 2562 596 2565 613
rect 2554 593 2565 596
rect 2554 526 2557 593
rect 2570 533 2573 546
rect 2586 543 2589 726
rect 2610 693 2613 736
rect 2618 733 2629 736
rect 2618 613 2621 726
rect 2626 613 2629 696
rect 2634 636 2637 726
rect 2642 723 2645 803
rect 2634 633 2645 636
rect 2642 613 2645 633
rect 2546 523 2557 526
rect 2562 513 2565 526
rect 2506 343 2517 346
rect 2458 313 2469 316
rect 2366 283 2373 286
rect 2314 243 2321 246
rect 2314 206 2317 243
rect 2322 213 2325 226
rect 2370 213 2373 283
rect 2458 246 2461 313
rect 2458 243 2469 246
rect 2314 203 2325 206
rect 2322 166 2325 203
rect 2322 163 2329 166
rect 2326 106 2329 163
rect 2338 123 2341 186
rect 2326 103 2333 106
rect 2330 36 2333 103
rect 2322 33 2333 36
rect 2322 13 2325 33
rect 2362 13 2365 146
rect 2386 143 2389 206
rect 2386 3 2389 126
rect 2410 123 2413 226
rect 2458 133 2461 226
rect 2466 213 2469 243
rect 2474 203 2477 316
rect 2482 123 2485 216
rect 2490 213 2493 336
rect 2514 256 2517 343
rect 2538 333 2541 416
rect 2578 393 2581 406
rect 2594 386 2597 526
rect 2650 523 2653 823
rect 2658 766 2661 883
rect 2698 813 2701 826
rect 2722 786 2725 903
rect 2738 813 2741 836
rect 2746 823 2749 926
rect 2722 783 2733 786
rect 2658 763 2665 766
rect 2662 666 2665 763
rect 2706 723 2709 736
rect 2658 663 2665 666
rect 2658 603 2661 663
rect 2674 533 2677 546
rect 2730 543 2733 783
rect 2762 723 2765 926
rect 2866 923 2877 926
rect 2810 813 2813 826
rect 2850 813 2853 886
rect 2866 846 2869 923
rect 2858 843 2869 846
rect 2962 846 2965 1016
rect 2970 1013 2973 1026
rect 3018 1016 3021 1123
rect 3026 1103 3029 1126
rect 3010 1013 3021 1016
rect 3026 1013 3029 1036
rect 2978 946 2981 1006
rect 2986 973 2989 1006
rect 2978 943 2989 946
rect 2986 846 2989 943
rect 2962 843 2973 846
rect 2858 813 2861 843
rect 2834 783 2837 806
rect 2850 733 2853 806
rect 2874 746 2877 816
rect 2898 776 2901 816
rect 2970 803 2973 843
rect 2978 843 2989 846
rect 2978 823 2981 843
rect 2978 796 2981 806
rect 2898 773 2909 776
rect 2874 743 2885 746
rect 2858 733 2877 736
rect 2738 613 2741 636
rect 2762 566 2765 606
rect 2802 603 2805 726
rect 2850 706 2853 726
rect 2842 703 2853 706
rect 2842 646 2845 703
rect 2842 643 2853 646
rect 2850 613 2853 643
rect 2866 633 2869 726
rect 2690 513 2693 526
rect 2746 523 2749 566
rect 2762 563 2773 566
rect 2874 563 2877 733
rect 2882 723 2885 743
rect 2890 723 2893 736
rect 2906 716 2909 773
rect 2898 713 2909 716
rect 2898 613 2901 713
rect 2770 533 2773 563
rect 2618 403 2621 416
rect 2570 313 2573 326
rect 2506 253 2517 256
rect 2506 183 2509 253
rect 2514 213 2517 226
rect 2514 126 2517 206
rect 2522 193 2525 236
rect 2530 203 2549 206
rect 2530 166 2533 186
rect 2530 163 2541 166
rect 2498 123 2517 126
rect 2538 86 2541 163
rect 2554 123 2557 216
rect 2562 213 2565 236
rect 2562 193 2565 206
rect 2578 203 2581 386
rect 2586 383 2597 386
rect 2642 383 2645 416
rect 2586 313 2589 383
rect 2594 303 2597 336
rect 2586 176 2589 236
rect 2602 223 2605 346
rect 2642 316 2645 326
rect 2618 223 2621 236
rect 2626 216 2629 316
rect 2642 313 2653 316
rect 2658 313 2661 326
rect 2666 316 2669 356
rect 2698 346 2701 416
rect 2706 353 2709 416
rect 2762 403 2765 416
rect 2786 403 2789 546
rect 2882 533 2885 546
rect 2906 543 2909 556
rect 2802 443 2805 526
rect 2858 513 2861 526
rect 2898 513 2901 536
rect 2834 413 2837 436
rect 2850 426 2853 446
rect 2922 433 2925 606
rect 2946 446 2949 796
rect 2962 793 2981 796
rect 2994 733 2997 746
rect 2970 713 2973 726
rect 2978 703 2981 726
rect 2970 543 2973 626
rect 2994 623 2997 726
rect 3002 713 3005 736
rect 3010 723 3013 1013
rect 3018 983 3021 1006
rect 3026 926 3029 946
rect 3022 923 3029 926
rect 3022 816 3025 923
rect 3022 813 3029 816
rect 3026 793 3029 813
rect 3034 743 3037 1133
rect 3042 976 3045 1116
rect 3058 1113 3061 1143
rect 3066 1113 3069 1126
rect 3050 1023 3053 1036
rect 3074 1016 3077 1173
rect 3082 1133 3085 1156
rect 3082 1123 3101 1126
rect 3106 1123 3109 1136
rect 3082 1103 3085 1116
rect 3058 993 3061 1016
rect 3074 1013 3081 1016
rect 3090 1013 3093 1026
rect 3098 1013 3109 1016
rect 3066 983 3069 1006
rect 3042 973 3053 976
rect 3050 846 3053 973
rect 3078 966 3081 1013
rect 3098 1003 3109 1006
rect 3114 1003 3117 1026
rect 3098 983 3101 996
rect 3074 963 3081 966
rect 3074 943 3077 963
rect 3042 843 3053 846
rect 3042 763 3045 843
rect 3050 783 3053 816
rect 3058 813 3061 826
rect 3066 813 3069 936
rect 3082 926 3085 936
rect 3122 933 3125 1216
rect 3138 1176 3141 1223
rect 3130 1173 3141 1176
rect 3130 1126 3133 1173
rect 3146 1143 3149 1156
rect 3130 1123 3141 1126
rect 3138 1106 3141 1123
rect 3138 1103 3145 1106
rect 3142 966 3145 1103
rect 3138 963 3145 966
rect 3138 946 3141 963
rect 3130 943 3141 946
rect 3154 943 3157 1603
rect 3170 1513 3173 1536
rect 3178 1426 3181 1626
rect 3186 1533 3189 1706
rect 3194 1516 3197 1616
rect 3202 1603 3205 1716
rect 3210 1713 3213 1726
rect 3210 1693 3213 1706
rect 3218 1663 3221 1816
rect 3234 1746 3237 1823
rect 3226 1743 3237 1746
rect 3218 1623 3221 1636
rect 3226 1623 3229 1743
rect 3242 1636 3245 1726
rect 3234 1633 3245 1636
rect 3234 1613 3237 1633
rect 3210 1533 3213 1566
rect 3190 1513 3197 1516
rect 3190 1446 3193 1513
rect 3190 1443 3197 1446
rect 3162 1413 3165 1426
rect 3178 1423 3185 1426
rect 3170 1403 3173 1416
rect 3182 1376 3185 1423
rect 3178 1373 3185 1376
rect 3178 1353 3181 1373
rect 3170 1333 3173 1346
rect 3162 1313 3165 1326
rect 3170 1213 3173 1326
rect 3178 1313 3181 1336
rect 3194 1333 3197 1443
rect 3202 1366 3205 1526
rect 3210 1403 3213 1526
rect 3218 1453 3221 1586
rect 3250 1583 3253 1843
rect 3258 1813 3261 2026
rect 3266 1933 3269 2016
rect 3290 2013 3293 2036
rect 3298 2023 3301 2136
rect 3306 1993 3309 2226
rect 3314 1973 3317 2426
rect 3322 2406 3325 2433
rect 3330 2423 3333 2493
rect 3354 2486 3357 2503
rect 3346 2483 3357 2486
rect 3362 2503 3381 2506
rect 3386 2503 3389 2526
rect 3402 2513 3405 2586
rect 3346 2416 3349 2483
rect 3362 2416 3365 2503
rect 3418 2483 3421 2526
rect 3434 2523 3437 2776
rect 3450 2726 3453 2746
rect 3446 2723 3453 2726
rect 3446 2626 3449 2723
rect 3446 2623 3453 2626
rect 3450 2533 3453 2623
rect 3458 2526 3461 2823
rect 3466 2606 3469 2706
rect 3474 2673 3477 2943
rect 3482 2916 3485 2926
rect 3490 2923 3493 2936
rect 3498 2933 3501 2946
rect 3506 2916 3509 2926
rect 3482 2913 3509 2916
rect 3498 2896 3501 2913
rect 3490 2893 3501 2896
rect 3490 2826 3493 2893
rect 3506 2836 3509 2906
rect 3506 2833 3513 2836
rect 3490 2823 3501 2826
rect 3498 2803 3501 2823
rect 3482 2633 3485 2656
rect 3474 2613 3477 2626
rect 3490 2613 3493 2686
rect 3498 2653 3501 2756
rect 3510 2746 3513 2833
rect 3506 2743 3513 2746
rect 3466 2603 3477 2606
rect 3474 2546 3477 2603
rect 3474 2543 3481 2546
rect 3446 2523 3461 2526
rect 3370 2433 3381 2436
rect 3346 2413 3357 2416
rect 3362 2413 3373 2416
rect 3386 2413 3389 2426
rect 3426 2423 3429 2476
rect 3322 2403 3333 2406
rect 3330 2356 3333 2403
rect 3354 2396 3357 2413
rect 3322 2353 3333 2356
rect 3322 2333 3325 2353
rect 3346 2336 3349 2396
rect 3354 2393 3361 2396
rect 3338 2333 3349 2336
rect 3338 2236 3341 2333
rect 3358 2326 3361 2393
rect 3354 2323 3361 2326
rect 3354 2246 3357 2323
rect 3354 2243 3361 2246
rect 3322 2163 3325 2236
rect 3338 2233 3349 2236
rect 3346 2213 3349 2233
rect 3322 2116 3325 2136
rect 3322 2113 3329 2116
rect 3326 2026 3329 2113
rect 3338 2103 3341 2126
rect 3346 2123 3349 2206
rect 3358 2186 3361 2243
rect 3354 2183 3361 2186
rect 3354 2126 3357 2183
rect 3370 2166 3373 2413
rect 3386 2283 3389 2336
rect 3362 2163 3373 2166
rect 3362 2133 3365 2163
rect 3354 2123 3365 2126
rect 3362 2106 3365 2123
rect 3370 2113 3373 2126
rect 3354 2103 3365 2106
rect 3322 2023 3329 2026
rect 3322 1983 3325 2023
rect 3346 2013 3349 2026
rect 3330 1993 3333 2006
rect 3274 1923 3277 1946
rect 3306 1923 3309 1936
rect 3314 1913 3317 1926
rect 3266 1803 3269 1846
rect 3330 1813 3333 1926
rect 3354 1813 3357 2103
rect 3370 2003 3373 2086
rect 3386 1946 3389 2216
rect 3394 2213 3397 2326
rect 3402 2316 3405 2336
rect 3426 2323 3429 2336
rect 3402 2313 3413 2316
rect 3410 2266 3413 2313
rect 3402 2263 3413 2266
rect 3402 2206 3405 2263
rect 3418 2233 3421 2246
rect 3418 2213 3421 2226
rect 3402 2203 3413 2206
rect 3410 2123 3413 2203
rect 3434 2166 3437 2486
rect 3446 2456 3449 2523
rect 3458 2483 3461 2516
rect 3442 2453 3449 2456
rect 3442 2353 3445 2453
rect 3450 2403 3453 2436
rect 3458 2413 3461 2426
rect 3442 2313 3445 2336
rect 3458 2206 3461 2406
rect 3466 2346 3469 2536
rect 3478 2486 3481 2543
rect 3490 2503 3493 2556
rect 3498 2523 3501 2616
rect 3506 2513 3509 2743
rect 3514 2713 3517 2726
rect 3522 2703 3525 3056
rect 3546 3033 3549 3136
rect 3530 2993 3533 3016
rect 3538 2686 3541 2936
rect 3546 2916 3549 2936
rect 3554 2923 3557 3366
rect 3570 3333 3573 3366
rect 3594 3346 3597 3393
rect 3634 3376 3637 3443
rect 3666 3436 3669 3563
rect 3698 3523 3701 3556
rect 3706 3533 3709 3573
rect 3714 3506 3717 3716
rect 3722 3533 3725 3546
rect 3650 3433 3669 3436
rect 3706 3503 3717 3506
rect 3706 3436 3709 3503
rect 3730 3456 3733 4083
rect 3738 3923 3741 4006
rect 3746 3933 3749 3946
rect 3762 3863 3765 4076
rect 3786 3963 3789 4016
rect 3762 3773 3765 3816
rect 3738 3716 3741 3736
rect 3786 3733 3789 3776
rect 3802 3736 3805 4153
rect 3818 4133 3829 4136
rect 3850 4133 3853 4233
rect 3858 4223 3861 4323
rect 3898 4306 3901 4356
rect 3890 4303 3901 4306
rect 3866 4203 3869 4246
rect 3890 4236 3893 4303
rect 3910 4286 3913 4363
rect 3906 4283 3913 4286
rect 3906 4263 3909 4283
rect 3890 4233 3901 4236
rect 3882 4203 3885 4216
rect 3898 4203 3901 4233
rect 3818 4056 3821 4126
rect 3834 4113 3837 4126
rect 3866 4123 3869 4196
rect 3906 4153 3909 4216
rect 3914 4203 3917 4226
rect 3922 4213 3925 4326
rect 3954 4316 3957 4336
rect 3946 4313 3957 4316
rect 3946 4236 3949 4313
rect 3946 4233 3957 4236
rect 3954 4213 3957 4233
rect 3962 4206 3965 4336
rect 3986 4333 3989 4373
rect 3994 4323 3997 4416
rect 4002 4356 4005 4526
rect 4018 4423 4021 4536
rect 4026 4506 4029 4526
rect 4034 4523 4037 4536
rect 4074 4523 4077 4556
rect 4082 4533 4085 4606
rect 4098 4593 4101 4606
rect 4122 4603 4125 4616
rect 4114 4576 4117 4596
rect 4114 4573 4125 4576
rect 4090 4533 4101 4536
rect 4090 4513 4093 4526
rect 4098 4523 4101 4533
rect 4106 4523 4109 4556
rect 4122 4516 4125 4573
rect 4178 4533 4181 4616
rect 4218 4593 4221 4606
rect 4242 4596 4245 4616
rect 4234 4593 4245 4596
rect 4114 4513 4125 4516
rect 4026 4503 4037 4506
rect 4034 4436 4037 4503
rect 4026 4433 4037 4436
rect 4010 4393 4013 4416
rect 4002 4353 4013 4356
rect 4002 4333 4005 4346
rect 3994 4213 3997 4226
rect 3818 4053 3837 4056
rect 3834 3976 3837 4053
rect 3882 4026 3885 4136
rect 3890 4113 3893 4136
rect 3906 4043 3909 4126
rect 3922 4106 3925 4206
rect 3954 4203 3965 4206
rect 3938 4156 3941 4166
rect 3954 4163 3957 4203
rect 3938 4153 3973 4156
rect 3962 4113 3965 4136
rect 3970 4133 3973 4153
rect 3978 4106 3981 4156
rect 3882 4023 3893 4026
rect 3826 3973 3837 3976
rect 3826 3923 3829 3973
rect 3842 3883 3845 3936
rect 3858 3933 3861 3966
rect 3850 3923 3861 3926
rect 3818 3783 3821 3816
rect 3842 3793 3845 3866
rect 3802 3733 3813 3736
rect 3738 3713 3749 3716
rect 3746 3636 3749 3713
rect 3778 3706 3781 3726
rect 3770 3703 3781 3706
rect 3786 3706 3789 3726
rect 3786 3703 3797 3706
rect 3770 3656 3773 3703
rect 3770 3653 3781 3656
rect 3738 3633 3749 3636
rect 3738 3613 3741 3633
rect 3770 3613 3773 3636
rect 3730 3453 3741 3456
rect 3706 3433 3717 3436
rect 3634 3373 3645 3376
rect 3594 3343 3605 3346
rect 3602 3296 3605 3343
rect 3618 3323 3621 3336
rect 3594 3293 3605 3296
rect 3594 3276 3597 3293
rect 3562 3223 3565 3246
rect 3562 2986 3565 3166
rect 3570 3003 3573 3276
rect 3590 3273 3597 3276
rect 3590 3226 3593 3273
rect 3602 3233 3605 3256
rect 3590 3223 3597 3226
rect 3578 3116 3581 3136
rect 3594 3133 3597 3223
rect 3610 3203 3621 3206
rect 3578 3113 3589 3116
rect 3586 3036 3589 3113
rect 3578 3033 3589 3036
rect 3578 3013 3581 3033
rect 3562 2983 3573 2986
rect 3570 2926 3573 2983
rect 3586 2933 3589 3016
rect 3602 3013 3605 3116
rect 3618 3073 3621 3126
rect 3626 3113 3629 3126
rect 3634 3103 3637 3116
rect 3594 2993 3597 3006
rect 3610 2976 3613 3006
rect 3594 2973 3613 2976
rect 3594 2933 3597 2973
rect 3562 2923 3573 2926
rect 3546 2913 3557 2916
rect 3530 2683 3541 2686
rect 3514 2616 3517 2676
rect 3522 2623 3525 2646
rect 3514 2613 3525 2616
rect 3522 2546 3525 2613
rect 3530 2593 3533 2683
rect 3538 2613 3541 2626
rect 3546 2603 3549 2716
rect 3554 2546 3557 2913
rect 3562 2903 3565 2923
rect 3594 2906 3597 2926
rect 3586 2903 3597 2906
rect 3586 2836 3589 2903
rect 3562 2813 3565 2836
rect 3586 2833 3597 2836
rect 3578 2736 3581 2816
rect 3594 2743 3597 2833
rect 3602 2793 3605 2956
rect 3610 2923 3613 2966
rect 3618 2933 3621 2946
rect 3626 2906 3629 2926
rect 3618 2903 3629 2906
rect 3618 2846 3621 2903
rect 3618 2843 3629 2846
rect 3626 2823 3629 2843
rect 3562 2646 3565 2736
rect 3570 2733 3581 2736
rect 3610 2733 3613 2746
rect 3626 2733 3629 2806
rect 3634 2743 3637 3006
rect 3642 2823 3645 3373
rect 3650 3363 3653 3433
rect 3714 3416 3717 3433
rect 3658 3353 3661 3416
rect 3666 3333 3669 3406
rect 3682 3403 3685 3416
rect 3706 3413 3717 3416
rect 3690 3386 3693 3406
rect 3682 3383 3693 3386
rect 3674 3323 3677 3356
rect 3682 3333 3685 3383
rect 3682 3323 3693 3326
rect 3706 3323 3709 3356
rect 3682 3283 3685 3323
rect 3690 3156 3693 3316
rect 3706 3223 3709 3236
rect 3714 3203 3717 3326
rect 3722 3313 3725 3446
rect 3738 3376 3741 3453
rect 3730 3373 3741 3376
rect 3690 3153 3709 3156
rect 3682 3103 3685 3146
rect 3706 3036 3709 3153
rect 3730 3116 3733 3373
rect 3754 3136 3757 3606
rect 3762 3593 3765 3606
rect 3770 3533 3773 3606
rect 3778 3553 3781 3653
rect 3794 3626 3797 3703
rect 3786 3623 3797 3626
rect 3786 3603 3789 3623
rect 3778 3533 3789 3536
rect 3794 3533 3797 3606
rect 3778 3503 3781 3526
rect 3770 3403 3773 3416
rect 3778 3413 3781 3426
rect 3794 3366 3797 3526
rect 3810 3373 3813 3733
rect 3818 3713 3821 3736
rect 3850 3733 3853 3786
rect 3826 3723 3845 3726
rect 3850 3696 3853 3716
rect 3834 3693 3853 3696
rect 3834 3586 3837 3693
rect 3834 3583 3853 3586
rect 3818 3533 3821 3556
rect 3826 3413 3829 3566
rect 3834 3533 3837 3546
rect 3842 3523 3845 3536
rect 3850 3423 3853 3583
rect 3858 3563 3861 3923
rect 3866 3906 3869 4016
rect 3874 3993 3877 4016
rect 3890 3966 3893 4023
rect 3882 3963 3893 3966
rect 3882 3933 3885 3963
rect 3866 3903 3877 3906
rect 3874 3836 3877 3903
rect 3866 3833 3877 3836
rect 3866 3813 3869 3833
rect 3874 3796 3877 3816
rect 3874 3793 3881 3796
rect 3866 3683 3869 3766
rect 3878 3676 3881 3793
rect 3890 3713 3893 3936
rect 3914 3933 3917 4106
rect 3922 4103 3933 4106
rect 3930 4026 3933 4103
rect 3974 4103 3981 4106
rect 3974 4036 3977 4103
rect 3974 4033 3981 4036
rect 3986 4033 3989 4136
rect 4002 4133 4005 4166
rect 4010 4153 4013 4353
rect 4018 4333 4021 4416
rect 4026 4413 4029 4433
rect 4090 4413 4093 4426
rect 4026 4323 4029 4406
rect 4066 4323 4069 4346
rect 4042 4156 4045 4216
rect 4082 4163 4085 4306
rect 4114 4213 4117 4513
rect 4138 4393 4141 4406
rect 4154 4386 4157 4526
rect 4186 4456 4189 4526
rect 4194 4523 4197 4536
rect 4234 4533 4237 4593
rect 4226 4513 4229 4526
rect 4242 4523 4261 4526
rect 4182 4453 4189 4456
rect 4138 4383 4157 4386
rect 4130 4273 4133 4366
rect 4138 4333 4141 4383
rect 4122 4213 4125 4226
rect 4146 4213 4149 4336
rect 4154 4333 4157 4346
rect 4162 4323 4165 4406
rect 4170 4403 4173 4416
rect 4182 4406 4185 4453
rect 4194 4413 4197 4446
rect 4242 4436 4245 4523
rect 4218 4413 4221 4436
rect 4234 4433 4245 4436
rect 4182 4403 4189 4406
rect 4234 4403 4237 4433
rect 4170 4283 4173 4376
rect 4186 4313 4189 4403
rect 4250 4393 4253 4416
rect 4202 4253 4205 4336
rect 4226 4323 4229 4346
rect 4266 4323 4269 4536
rect 4298 4533 4301 4616
rect 4338 4593 4341 4606
rect 4290 4513 4293 4526
rect 4274 4393 4277 4416
rect 4282 4323 4285 4406
rect 4290 4333 4293 4406
rect 4306 4403 4309 4546
rect 4322 4523 4325 4536
rect 4330 4533 4333 4586
rect 4362 4583 4365 4616
rect 4338 4523 4341 4546
rect 4346 4523 4349 4556
rect 4362 4506 4365 4536
rect 4402 4533 4405 4546
rect 4418 4533 4421 4616
rect 4450 4593 4453 4616
rect 4498 4603 4501 4616
rect 4546 4606 4549 4616
rect 4354 4503 4365 4506
rect 4354 4446 4357 4503
rect 4354 4443 4365 4446
rect 4362 4426 4365 4443
rect 4338 4423 4365 4426
rect 4338 4413 4341 4423
rect 4346 4363 4349 4416
rect 4362 4413 4365 4423
rect 4370 4413 4373 4526
rect 4394 4483 4397 4526
rect 4298 4303 4301 4356
rect 4314 4313 4317 4326
rect 4322 4323 4325 4336
rect 4354 4333 4357 4406
rect 4370 4373 4373 4406
rect 4266 4233 4269 4296
rect 4194 4203 4197 4216
rect 4202 4203 4205 4216
rect 4034 4153 4045 4156
rect 3994 4113 3997 4126
rect 4010 4113 4013 4126
rect 4034 4056 4037 4153
rect 4130 4146 4133 4166
rect 4210 4156 4213 4216
rect 4218 4203 4221 4226
rect 4226 4203 4229 4216
rect 4202 4153 4213 4156
rect 4130 4143 4141 4146
rect 4034 4053 4045 4056
rect 4050 4053 4053 4136
rect 4066 4103 4069 4136
rect 4114 4113 4117 4126
rect 3930 4023 3949 4026
rect 3922 3993 3925 4016
rect 3946 3946 3949 4023
rect 3970 4003 3973 4016
rect 3978 3966 3981 4033
rect 4018 4013 4021 4036
rect 3994 3983 3997 4006
rect 3978 3963 3985 3966
rect 3942 3943 3949 3946
rect 3942 3896 3945 3943
rect 3938 3893 3945 3896
rect 3874 3673 3881 3676
rect 3874 3613 3877 3673
rect 3882 3593 3885 3616
rect 3898 3486 3901 3796
rect 3906 3723 3909 3816
rect 3914 3793 3917 3806
rect 3922 3803 3925 3886
rect 3914 3603 3917 3726
rect 3922 3523 3925 3546
rect 3898 3483 3909 3486
rect 3866 3423 3877 3426
rect 3858 3413 3877 3416
rect 3850 3403 3861 3406
rect 3874 3396 3877 3413
rect 3866 3393 3877 3396
rect 3794 3363 3813 3366
rect 3770 3313 3773 3326
rect 3794 3323 3797 3336
rect 3810 3323 3813 3363
rect 3778 3203 3781 3216
rect 3786 3213 3805 3216
rect 3642 2736 3645 2756
rect 3634 2733 3645 2736
rect 3570 2683 3573 2733
rect 3578 2706 3581 2726
rect 3610 2723 3621 2726
rect 3578 2703 3589 2706
rect 3562 2643 3573 2646
rect 3562 2613 3565 2626
rect 3570 2603 3573 2643
rect 3586 2626 3589 2703
rect 3578 2623 3589 2626
rect 3578 2603 3581 2623
rect 3522 2543 3533 2546
rect 3478 2483 3485 2486
rect 3482 2436 3485 2483
rect 3514 2453 3517 2536
rect 3530 2466 3533 2543
rect 3522 2463 3533 2466
rect 3546 2543 3557 2546
rect 3474 2433 3485 2436
rect 3474 2413 3477 2433
rect 3498 2376 3501 2416
rect 3506 2403 3509 2416
rect 3522 2376 3525 2463
rect 3546 2403 3549 2543
rect 3554 2506 3557 2536
rect 3570 2533 3573 2596
rect 3562 2523 3589 2526
rect 3570 2513 3581 2516
rect 3554 2503 3561 2506
rect 3558 2436 3561 2503
rect 3554 2433 3561 2436
rect 3554 2413 3557 2433
rect 3570 2376 3573 2513
rect 3586 2413 3589 2523
rect 3602 2413 3605 2536
rect 3618 2426 3621 2536
rect 3610 2423 3621 2426
rect 3610 2406 3613 2423
rect 3602 2403 3613 2406
rect 3498 2373 3517 2376
rect 3522 2373 3541 2376
rect 3570 2373 3581 2376
rect 3466 2343 3477 2346
rect 3466 2303 3469 2326
rect 3474 2213 3477 2343
rect 3482 2243 3485 2326
rect 3490 2306 3493 2356
rect 3498 2323 3501 2346
rect 3490 2303 3501 2306
rect 3498 2236 3501 2303
rect 3490 2233 3501 2236
rect 3490 2216 3493 2233
rect 3482 2213 3493 2216
rect 3426 2163 3437 2166
rect 3454 2203 3461 2206
rect 3426 2086 3429 2163
rect 3454 2136 3457 2203
rect 3454 2133 3461 2136
rect 3458 2116 3461 2133
rect 3466 2123 3469 2206
rect 3474 2133 3477 2196
rect 3482 2176 3485 2213
rect 3490 2193 3493 2206
rect 3498 2203 3501 2216
rect 3482 2173 3493 2176
rect 3474 2116 3477 2126
rect 3458 2113 3477 2116
rect 3474 2096 3477 2113
rect 3466 2093 3477 2096
rect 3426 2083 3437 2086
rect 3402 2013 3405 2026
rect 3386 1943 3397 1946
rect 3370 1813 3373 1936
rect 3394 1866 3397 1943
rect 3418 1933 3421 2016
rect 3426 1966 3429 2006
rect 3434 1986 3437 2083
rect 3466 2036 3469 2093
rect 3490 2086 3493 2173
rect 3514 2146 3517 2373
rect 3522 2333 3525 2356
rect 3538 2333 3541 2373
rect 3522 2213 3525 2226
rect 3530 2203 3533 2306
rect 3570 2303 3573 2326
rect 3538 2203 3541 2226
rect 3570 2213 3573 2226
rect 3486 2083 3493 2086
rect 3506 2143 3517 2146
rect 3546 2143 3549 2206
rect 3554 2203 3565 2206
rect 3578 2146 3581 2373
rect 3602 2366 3605 2403
rect 3618 2383 3621 2406
rect 3626 2403 3629 2456
rect 3634 2413 3637 2726
rect 3650 2723 3653 2966
rect 3658 2833 3661 3026
rect 3674 3013 3677 3036
rect 3690 3033 3709 3036
rect 3722 3113 3733 3116
rect 3750 3133 3757 3136
rect 3682 2993 3685 3006
rect 3690 2966 3693 3033
rect 3698 3003 3701 3016
rect 3686 2963 3693 2966
rect 3706 2963 3709 3016
rect 3722 3006 3725 3113
rect 3738 3013 3741 3106
rect 3750 3076 3753 3133
rect 3762 3096 3765 3126
rect 3770 3103 3773 3116
rect 3778 3113 3781 3156
rect 3802 3136 3805 3213
rect 3810 3203 3813 3316
rect 3818 3213 3821 3226
rect 3826 3193 3829 3206
rect 3802 3133 3813 3136
rect 3794 3123 3805 3126
rect 3786 3113 3797 3116
rect 3786 3096 3789 3106
rect 3762 3093 3789 3096
rect 3750 3073 3757 3076
rect 3754 3053 3757 3073
rect 3818 3056 3821 3156
rect 3786 3036 3789 3056
rect 3818 3053 3825 3056
rect 3834 3053 3837 3376
rect 3866 3336 3869 3393
rect 3858 3333 3869 3336
rect 3882 3333 3885 3426
rect 3890 3383 3893 3406
rect 3906 3403 3909 3483
rect 3938 3443 3941 3893
rect 3946 3813 3949 3826
rect 3954 3803 3957 3926
rect 3982 3886 3985 3963
rect 4018 3933 4021 3946
rect 3978 3883 3985 3886
rect 3978 3823 3981 3883
rect 3962 3813 3981 3816
rect 3962 3793 3965 3813
rect 3986 3793 3989 3806
rect 3994 3803 3997 3926
rect 3970 3696 3973 3716
rect 3994 3713 3997 3726
rect 3962 3693 3973 3696
rect 3962 3636 3965 3693
rect 3962 3633 3973 3636
rect 3946 3613 3965 3616
rect 3954 3583 3957 3606
rect 3970 3603 3973 3633
rect 3986 3603 3989 3686
rect 4010 3613 4013 3826
rect 4034 3803 4037 3856
rect 4042 3816 4045 4053
rect 4074 4013 4077 4056
rect 4050 3853 4053 3976
rect 4058 3906 4061 3926
rect 4098 3906 4101 3926
rect 4058 3903 4065 3906
rect 4062 3836 4065 3903
rect 4058 3833 4065 3836
rect 4090 3903 4101 3906
rect 4090 3836 4093 3903
rect 4090 3833 4101 3836
rect 4042 3813 4053 3816
rect 4050 3786 4053 3813
rect 4058 3803 4061 3833
rect 4066 3813 4085 3816
rect 4042 3783 4053 3786
rect 3994 3546 3997 3606
rect 3994 3543 4005 3546
rect 3994 3523 3997 3536
rect 3930 3403 3933 3416
rect 3850 3286 3853 3326
rect 3866 3303 3869 3326
rect 3850 3283 3861 3286
rect 3858 3186 3861 3283
rect 3850 3183 3861 3186
rect 3850 3163 3853 3183
rect 3882 3153 3885 3326
rect 3898 3323 3901 3336
rect 3906 3323 3909 3366
rect 3946 3333 3949 3406
rect 3970 3366 3973 3446
rect 3986 3403 3989 3416
rect 3994 3403 3997 3416
rect 3966 3363 3973 3366
rect 3898 3213 3901 3236
rect 3890 3193 3893 3206
rect 3914 3176 3917 3316
rect 3954 3306 3957 3326
rect 3946 3303 3957 3306
rect 3946 3246 3949 3303
rect 3966 3286 3969 3363
rect 4002 3336 4005 3543
rect 4026 3413 4029 3616
rect 4042 3593 4045 3783
rect 4074 3696 4077 3806
rect 4098 3803 4101 3833
rect 4066 3693 4077 3696
rect 4066 3636 4069 3693
rect 4066 3633 4077 3636
rect 4090 3633 4093 3706
rect 4106 3653 4109 4106
rect 4138 4086 4141 4143
rect 4186 4123 4189 4136
rect 4194 4123 4197 4146
rect 4202 4093 4205 4153
rect 4210 4113 4213 4136
rect 4218 4123 4221 4136
rect 4234 4106 4237 4206
rect 4250 4126 4253 4226
rect 4218 4103 4237 4106
rect 4246 4123 4253 4126
rect 4130 4083 4141 4086
rect 4130 4046 4133 4083
rect 4130 4043 4141 4046
rect 4138 3996 4141 4043
rect 4130 3993 4141 3996
rect 4154 3993 4157 4016
rect 4130 3933 4133 3993
rect 4178 3913 4181 3926
rect 4114 3813 4117 3846
rect 4138 3803 4149 3806
rect 4074 3616 4077 3633
rect 4050 3533 4053 3606
rect 4058 3603 4061 3616
rect 4066 3613 4077 3616
rect 4066 3526 4069 3613
rect 4082 3573 4085 3626
rect 4098 3613 4101 3646
rect 4050 3523 4069 3526
rect 4042 3413 4045 3426
rect 4034 3403 4045 3406
rect 3994 3333 4005 3336
rect 4034 3333 4037 3366
rect 4050 3353 4053 3523
rect 4090 3486 4093 3596
rect 4114 3583 4117 3626
rect 4122 3603 4125 3616
rect 4130 3586 4133 3736
rect 4146 3733 4149 3803
rect 4162 3786 4165 3806
rect 4158 3783 4165 3786
rect 4158 3716 4161 3783
rect 4170 3733 4173 3816
rect 4178 3783 4181 3886
rect 4194 3876 4197 4006
rect 4202 3956 4205 4016
rect 4210 3973 4213 4026
rect 4202 3953 4209 3956
rect 4190 3873 4197 3876
rect 4158 3713 4165 3716
rect 4162 3696 4165 3713
rect 4162 3693 4181 3696
rect 4138 3593 4141 3606
rect 4154 3603 4157 3656
rect 4178 3613 4181 3693
rect 4190 3676 4193 3873
rect 4206 3866 4209 3953
rect 4218 3883 4221 4103
rect 4226 4013 4229 4026
rect 4234 4013 4237 4096
rect 4246 4036 4249 4123
rect 4258 4036 4261 4116
rect 4266 4103 4269 4226
rect 4274 4213 4277 4246
rect 4290 4223 4317 4226
rect 4314 4213 4317 4223
rect 4274 4113 4277 4126
rect 4282 4103 4285 4116
rect 4246 4033 4253 4036
rect 4258 4033 4277 4036
rect 4226 3923 4229 3946
rect 4234 3933 4237 3956
rect 4202 3863 4209 3866
rect 4190 3673 4197 3676
rect 4126 3583 4133 3586
rect 4114 3523 4117 3536
rect 4090 3483 4101 3486
rect 4098 3403 4101 3483
rect 4126 3436 4129 3583
rect 4138 3446 4141 3576
rect 4162 3456 4165 3546
rect 4170 3523 4173 3596
rect 4186 3533 4189 3656
rect 4194 3573 4197 3673
rect 4202 3543 4205 3863
rect 4218 3656 4221 3856
rect 4234 3746 4237 3926
rect 4242 3923 4245 4016
rect 4250 4013 4253 4033
rect 4258 4013 4261 4026
rect 4250 3993 4253 4006
rect 4250 3913 4253 3936
rect 4230 3743 4237 3746
rect 4250 3746 4253 3816
rect 4258 3803 4261 3926
rect 4266 3883 4269 4006
rect 4274 3956 4277 4033
rect 4282 4003 4285 4026
rect 4274 3953 4285 3956
rect 4274 3933 4277 3946
rect 4282 3936 4285 3953
rect 4282 3933 4289 3936
rect 4274 3893 4277 3926
rect 4286 3886 4289 3933
rect 4298 3916 4301 4206
rect 4306 4203 4317 4206
rect 4306 4133 4317 4136
rect 4314 4103 4317 4126
rect 4314 4013 4317 4036
rect 4314 3933 4317 3976
rect 4298 3913 4309 3916
rect 4282 3883 4289 3886
rect 4282 3836 4285 3883
rect 4306 3836 4309 3913
rect 4330 3853 4333 4216
rect 4346 3876 4349 4316
rect 4378 4283 4381 4436
rect 4410 4433 4413 4526
rect 4426 4523 4429 4546
rect 4442 4523 4445 4536
rect 4410 4403 4413 4416
rect 4418 4383 4421 4416
rect 4434 4406 4437 4466
rect 4426 4403 4437 4406
rect 4442 4363 4445 4416
rect 4450 4403 4453 4426
rect 4458 4393 4461 4536
rect 4522 4523 4525 4536
rect 4530 4533 4533 4606
rect 4538 4603 4549 4606
rect 4482 4413 4485 4426
rect 4498 4413 4501 4426
rect 4394 4323 4397 4336
rect 4354 4203 4357 4226
rect 4362 4203 4365 4236
rect 4370 4146 4373 4256
rect 4386 4213 4389 4226
rect 4378 4193 4381 4206
rect 4370 4143 4381 4146
rect 4362 4113 4365 4136
rect 4370 4123 4373 4136
rect 4370 4033 4373 4066
rect 4378 4046 4381 4143
rect 4386 4133 4389 4146
rect 4394 4136 4397 4306
rect 4410 4266 4413 4286
rect 4406 4263 4413 4266
rect 4406 4186 4409 4263
rect 4418 4253 4421 4336
rect 4450 4323 4453 4336
rect 4474 4323 4477 4406
rect 4490 4373 4493 4406
rect 4522 4403 4525 4416
rect 4538 4413 4541 4603
rect 4546 4533 4549 4556
rect 4562 4533 4565 4556
rect 4554 4513 4557 4526
rect 4570 4523 4573 4566
rect 4586 4466 4589 4526
rect 4594 4523 4597 4536
rect 4586 4463 4597 4466
rect 4594 4446 4597 4463
rect 4586 4443 4597 4446
rect 4530 4323 4533 4406
rect 4538 4373 4541 4406
rect 4406 4183 4413 4186
rect 4410 4136 4413 4183
rect 4426 4156 4429 4266
rect 4538 4233 4541 4336
rect 4546 4306 4549 4326
rect 4562 4323 4565 4416
rect 4570 4373 4573 4406
rect 4586 4356 4589 4443
rect 4602 4413 4605 4536
rect 4610 4493 4613 4536
rect 4610 4393 4613 4406
rect 4618 4403 4621 4416
rect 4626 4403 4629 4496
rect 4650 4386 4653 4526
rect 4658 4523 4661 4616
rect 4682 4603 4685 4616
rect 4682 4533 4685 4596
rect 4706 4593 4709 4616
rect 4674 4513 4677 4526
rect 4690 4523 4693 4556
rect 4778 4553 4781 4616
rect 4698 4533 4701 4546
rect 4738 4533 4741 4546
rect 4642 4383 4653 4386
rect 4586 4353 4597 4356
rect 4546 4303 4553 4306
rect 4550 4236 4553 4303
rect 4546 4233 4553 4236
rect 4450 4193 4453 4216
rect 4522 4213 4525 4226
rect 4546 4216 4549 4233
rect 4562 4216 4565 4246
rect 4570 4223 4573 4336
rect 4594 4333 4597 4353
rect 4578 4323 4597 4326
rect 4578 4306 4581 4323
rect 4602 4316 4605 4376
rect 4578 4303 4585 4306
rect 4582 4226 4585 4303
rect 4578 4223 4585 4226
rect 4538 4213 4549 4216
rect 4466 4166 4469 4186
rect 4466 4163 4473 4166
rect 4426 4153 4437 4156
rect 4394 4133 4405 4136
rect 4410 4133 4421 4136
rect 4378 4043 4389 4046
rect 4354 4013 4357 4026
rect 4354 4003 4365 4006
rect 4354 3913 4357 3936
rect 4362 3923 4365 4003
rect 4346 3873 4357 3876
rect 4354 3856 4357 3873
rect 4354 3853 4361 3856
rect 4266 3833 4285 3836
rect 4298 3833 4309 3836
rect 4330 3833 4341 3836
rect 4250 3743 4257 3746
rect 4230 3676 4233 3743
rect 4230 3673 4237 3676
rect 4218 3653 4225 3656
rect 4222 3576 4225 3653
rect 4218 3573 4225 3576
rect 4218 3496 4221 3573
rect 4202 3493 4221 3496
rect 4162 3453 4169 3456
rect 4138 3443 4145 3446
rect 4126 3433 4133 3436
rect 4122 3403 4125 3416
rect 4130 3386 4133 3433
rect 4126 3383 4133 3386
rect 3966 3283 3973 3286
rect 3946 3243 3957 3246
rect 3930 3193 3933 3216
rect 3938 3203 3941 3226
rect 3954 3203 3957 3243
rect 3890 3173 3917 3176
rect 3890 3146 3893 3173
rect 3922 3166 3925 3176
rect 3866 3143 3893 3146
rect 3850 3106 3853 3126
rect 3842 3103 3853 3106
rect 3858 3103 3861 3136
rect 3866 3133 3869 3143
rect 3786 3033 3793 3036
rect 3722 3003 3733 3006
rect 3666 2906 3669 2926
rect 3666 2903 3677 2906
rect 3674 2826 3677 2903
rect 3686 2886 3689 2963
rect 3706 2923 3709 2946
rect 3714 2916 3717 2956
rect 3730 2946 3733 3003
rect 3754 2953 3757 3006
rect 3778 2993 3781 3016
rect 3790 2986 3793 3033
rect 3822 2986 3825 3053
rect 3866 3043 3869 3126
rect 3882 3103 3885 3126
rect 3858 3013 3861 3036
rect 3866 2996 3869 3016
rect 3858 2993 3869 2996
rect 3786 2983 3793 2986
rect 3818 2983 3825 2986
rect 3706 2913 3717 2916
rect 3726 2943 3733 2946
rect 3686 2883 3693 2886
rect 3690 2836 3693 2883
rect 3666 2823 3677 2826
rect 3686 2833 3693 2836
rect 3666 2803 3669 2823
rect 3686 2786 3689 2833
rect 3682 2783 3689 2786
rect 3650 2413 3653 2436
rect 3602 2363 3609 2366
rect 3606 2286 3609 2363
rect 3602 2283 3609 2286
rect 3602 2256 3605 2283
rect 3602 2253 3609 2256
rect 3586 2213 3589 2226
rect 3450 2023 3453 2036
rect 3466 2033 3477 2036
rect 3442 2003 3445 2016
rect 3474 2013 3477 2033
rect 3486 2006 3489 2083
rect 3498 2033 3501 2056
rect 3506 2026 3509 2143
rect 3514 2033 3517 2136
rect 3506 2023 3517 2026
rect 3482 2003 3489 2006
rect 3434 1983 3453 1986
rect 3426 1963 3437 1966
rect 3434 1906 3437 1963
rect 3426 1903 3437 1906
rect 3426 1886 3429 1903
rect 3386 1863 3397 1866
rect 3418 1883 3429 1886
rect 3258 1736 3261 1756
rect 3258 1733 3265 1736
rect 3262 1646 3265 1733
rect 3258 1643 3265 1646
rect 3258 1553 3261 1643
rect 3226 1523 3229 1536
rect 3266 1533 3269 1626
rect 3274 1613 3277 1806
rect 3338 1773 3341 1806
rect 3386 1793 3389 1863
rect 3418 1836 3421 1883
rect 3450 1876 3453 1983
rect 3434 1873 3453 1876
rect 3434 1853 3437 1873
rect 3482 1836 3485 2003
rect 3498 1923 3501 1936
rect 3506 1923 3509 2016
rect 3514 1926 3517 2023
rect 3522 1933 3525 2126
rect 3530 2083 3533 2136
rect 3562 2126 3565 2146
rect 3570 2143 3581 2146
rect 3594 2143 3597 2246
rect 3606 2176 3609 2253
rect 3618 2203 3621 2326
rect 3626 2323 3629 2336
rect 3634 2243 3637 2406
rect 3642 2393 3645 2406
rect 3658 2403 3661 2746
rect 3682 2606 3685 2783
rect 3698 2766 3701 2826
rect 3694 2763 3701 2766
rect 3694 2696 3697 2763
rect 3706 2706 3709 2913
rect 3726 2896 3729 2943
rect 3726 2893 3733 2896
rect 3714 2833 3717 2846
rect 3730 2823 3733 2893
rect 3754 2806 3757 2936
rect 3786 2826 3789 2983
rect 3818 2966 3821 2983
rect 3810 2963 3821 2966
rect 3810 2876 3813 2963
rect 3834 2886 3837 2986
rect 3858 2916 3861 2993
rect 3882 2923 3885 3056
rect 3898 2946 3901 3166
rect 3914 3163 3925 3166
rect 3906 3133 3909 3156
rect 3914 3133 3917 3163
rect 3930 3133 3933 3146
rect 3906 3123 3925 3126
rect 3938 3123 3941 3166
rect 3946 3053 3949 3186
rect 3970 3166 3973 3283
rect 3994 3266 3997 3333
rect 4010 3276 4013 3326
rect 4010 3273 4021 3276
rect 3994 3263 4001 3266
rect 3986 3183 3989 3216
rect 3998 3166 4001 3263
rect 4010 3193 4013 3216
rect 4018 3203 4021 3273
rect 4026 3186 4029 3236
rect 4034 3203 4037 3326
rect 4042 3193 4045 3206
rect 3970 3163 3981 3166
rect 3954 3123 3957 3156
rect 3978 3116 3981 3163
rect 3970 3113 3981 3116
rect 3994 3163 4001 3166
rect 4010 3183 4029 3186
rect 3890 2943 3901 2946
rect 3858 2913 3869 2916
rect 3834 2883 3845 2886
rect 3810 2873 3821 2876
rect 3794 2833 3797 2856
rect 3786 2823 3797 2826
rect 3746 2803 3757 2806
rect 3746 2756 3749 2803
rect 3746 2753 3757 2756
rect 3706 2703 3713 2706
rect 3694 2693 3701 2696
rect 3698 2616 3701 2693
rect 3710 2636 3713 2703
rect 3710 2633 3717 2636
rect 3698 2613 3705 2616
rect 3682 2603 3693 2606
rect 3690 2583 3693 2603
rect 3674 2513 3677 2526
rect 3690 2523 3693 2536
rect 3702 2516 3705 2613
rect 3698 2513 3705 2516
rect 3666 2403 3669 2456
rect 3698 2453 3701 2513
rect 3642 2306 3645 2386
rect 3658 2313 3661 2336
rect 3666 2323 3669 2356
rect 3642 2303 3649 2306
rect 3646 2236 3649 2303
rect 3642 2233 3649 2236
rect 3626 2183 3629 2206
rect 3602 2173 3609 2176
rect 3570 2133 3573 2143
rect 3554 2123 3565 2126
rect 3530 1976 3533 2036
rect 3554 2026 3557 2123
rect 3554 2023 3565 2026
rect 3578 2023 3581 2136
rect 3538 1993 3541 2006
rect 3530 1973 3537 1976
rect 3514 1923 3525 1926
rect 3522 1893 3525 1923
rect 3418 1833 3429 1836
rect 3426 1813 3429 1833
rect 3474 1833 3485 1836
rect 3450 1793 3453 1806
rect 3474 1786 3477 1833
rect 3522 1806 3525 1856
rect 3534 1836 3537 1973
rect 3530 1833 3537 1836
rect 3530 1813 3533 1833
rect 3498 1793 3501 1806
rect 3522 1803 3533 1806
rect 3474 1783 3485 1786
rect 3298 1726 3301 1746
rect 3282 1713 3285 1726
rect 3290 1723 3301 1726
rect 3290 1696 3293 1723
rect 3386 1696 3389 1726
rect 3394 1706 3397 1776
rect 3402 1733 3405 1746
rect 3410 1723 3413 1736
rect 3434 1733 3437 1746
rect 3426 1713 3429 1726
rect 3394 1703 3405 1706
rect 3434 1703 3437 1726
rect 3466 1706 3469 1726
rect 3458 1703 3469 1706
rect 3474 1706 3477 1736
rect 3482 1733 3485 1783
rect 3498 1733 3509 1736
rect 3514 1733 3517 1746
rect 3482 1723 3501 1726
rect 3506 1706 3509 1733
rect 3530 1726 3533 1803
rect 3474 1703 3485 1706
rect 3290 1693 3301 1696
rect 3298 1636 3301 1693
rect 3378 1693 3389 1696
rect 3378 1646 3381 1693
rect 3378 1643 3389 1646
rect 3290 1633 3301 1636
rect 3290 1613 3293 1633
rect 3274 1593 3277 1606
rect 3314 1523 3317 1546
rect 3258 1486 3261 1506
rect 3258 1483 3265 1486
rect 3250 1436 3253 1456
rect 3218 1413 3221 1436
rect 3246 1433 3253 1436
rect 3226 1373 3229 1406
rect 3234 1383 3237 1406
rect 3202 1363 3213 1366
rect 3202 1333 3205 1356
rect 3186 1223 3189 1326
rect 3210 1303 3213 1363
rect 3226 1323 3229 1366
rect 3246 1346 3249 1433
rect 3262 1426 3265 1483
rect 3258 1423 3265 1426
rect 3246 1343 3253 1346
rect 3242 1313 3245 1326
rect 3250 1296 3253 1343
rect 3258 1333 3261 1423
rect 3274 1383 3277 1416
rect 3282 1413 3285 1506
rect 3322 1496 3325 1546
rect 3330 1533 3333 1626
rect 3386 1623 3389 1643
rect 3386 1596 3389 1616
rect 3402 1596 3405 1703
rect 3458 1636 3461 1703
rect 3458 1633 3469 1636
rect 3338 1543 3341 1596
rect 3378 1593 3389 1596
rect 3394 1593 3405 1596
rect 3426 1593 3429 1606
rect 3378 1546 3381 1593
rect 3378 1543 3385 1546
rect 3314 1493 3325 1496
rect 3314 1426 3317 1493
rect 3314 1423 3325 1426
rect 3266 1326 3269 1346
rect 3266 1323 3273 1326
rect 3234 1293 3253 1296
rect 3234 1176 3237 1293
rect 3258 1276 3261 1316
rect 3250 1273 3261 1276
rect 3250 1206 3253 1273
rect 3270 1266 3273 1323
rect 3266 1263 3273 1266
rect 3266 1213 3269 1263
rect 3282 1246 3285 1376
rect 3290 1316 3293 1396
rect 3298 1333 3301 1406
rect 3322 1393 3325 1423
rect 3330 1356 3333 1526
rect 3338 1413 3341 1536
rect 3346 1413 3357 1416
rect 3322 1353 3333 1356
rect 3290 1313 3297 1316
rect 3278 1243 3285 1246
rect 3250 1203 3261 1206
rect 3234 1173 3245 1176
rect 3218 1136 3221 1156
rect 3210 1133 3221 1136
rect 3162 953 3165 1116
rect 3178 1106 3181 1126
rect 3202 1113 3205 1126
rect 3178 1103 3197 1106
rect 3074 903 3077 926
rect 3082 923 3101 926
rect 3098 906 3101 923
rect 3094 903 3101 906
rect 3094 846 3097 903
rect 3094 843 3101 846
rect 3090 806 3093 826
rect 3082 803 3093 806
rect 3042 733 3045 756
rect 3066 733 3069 776
rect 3042 723 3061 726
rect 3018 703 3021 716
rect 2986 613 3005 616
rect 3010 613 3013 636
rect 3042 603 3045 646
rect 2970 523 2973 536
rect 2978 516 2981 556
rect 3042 543 3045 556
rect 2978 513 2989 516
rect 2938 443 2949 446
rect 2850 423 2857 426
rect 2674 333 2677 346
rect 2698 343 2709 346
rect 2706 323 2709 343
rect 2730 333 2733 346
rect 2746 333 2749 396
rect 2802 393 2805 406
rect 2842 333 2845 416
rect 2854 356 2857 423
rect 2898 413 2901 426
rect 2922 376 2925 416
rect 2938 403 2941 443
rect 2922 373 2941 376
rect 2850 353 2857 356
rect 2850 333 2853 353
rect 2666 313 2677 316
rect 2602 213 2629 216
rect 2634 213 2637 226
rect 2650 213 2653 313
rect 2674 236 2677 313
rect 2666 233 2677 236
rect 2666 213 2669 233
rect 2618 193 2621 206
rect 2626 203 2629 213
rect 2714 203 2717 286
rect 2722 203 2725 226
rect 2746 223 2757 226
rect 2586 173 2597 176
rect 2578 133 2581 146
rect 2594 113 2597 173
rect 2634 123 2637 136
rect 2642 133 2645 196
rect 2658 123 2661 146
rect 2706 123 2709 146
rect 2762 123 2765 216
rect 2770 183 2773 206
rect 2778 193 2781 206
rect 2786 186 2789 216
rect 2794 203 2797 326
rect 2778 183 2789 186
rect 2770 133 2773 146
rect 2778 123 2781 183
rect 2802 113 2805 216
rect 2818 193 2821 216
rect 2826 213 2829 326
rect 2834 306 2837 326
rect 2834 303 2845 306
rect 2842 236 2845 303
rect 2834 233 2845 236
rect 2834 203 2837 233
rect 2850 203 2853 216
rect 2866 203 2869 336
rect 2874 283 2877 326
rect 2842 133 2845 146
rect 2858 133 2869 136
rect 2874 126 2877 136
rect 2890 133 2893 336
rect 2914 213 2917 226
rect 2906 153 2909 206
rect 2922 203 2925 336
rect 2938 333 2941 373
rect 2962 323 2965 406
rect 2986 403 2989 513
rect 3010 506 3013 526
rect 3002 503 3013 506
rect 3018 506 3021 526
rect 3018 503 3029 506
rect 3002 446 3005 503
rect 3026 456 3029 503
rect 3018 453 3029 456
rect 3002 443 3013 446
rect 2994 403 2997 426
rect 3010 393 3013 443
rect 3018 423 3021 453
rect 3042 416 3045 436
rect 3050 433 3053 536
rect 3066 513 3069 526
rect 3050 423 3069 426
rect 3042 413 3053 416
rect 3066 413 3069 423
rect 3026 333 3029 346
rect 3026 316 3029 326
rect 3042 323 3045 346
rect 3050 326 3053 413
rect 3082 403 3085 803
rect 3098 723 3101 843
rect 3106 833 3109 926
rect 3114 903 3117 916
rect 3114 813 3117 826
rect 3122 743 3125 756
rect 3130 726 3133 943
rect 3154 933 3165 936
rect 3146 913 3149 926
rect 3154 896 3157 926
rect 3146 893 3157 896
rect 3146 756 3149 893
rect 3146 753 3157 756
rect 3122 723 3133 726
rect 3122 666 3125 723
rect 3138 706 3141 736
rect 3146 713 3149 726
rect 3138 703 3145 706
rect 3122 663 3133 666
rect 3130 643 3133 663
rect 3142 646 3145 703
rect 3142 643 3149 646
rect 3098 403 3101 636
rect 3114 583 3117 606
rect 3106 513 3109 526
rect 3122 503 3125 616
rect 3138 613 3141 626
rect 3146 603 3149 643
rect 3154 596 3157 753
rect 3162 706 3165 916
rect 3170 903 3173 1016
rect 3178 1013 3181 1036
rect 3178 923 3181 996
rect 3186 963 3189 1006
rect 3210 993 3213 1016
rect 3218 933 3221 1116
rect 3226 1103 3229 1116
rect 3242 1046 3245 1173
rect 3258 1056 3261 1203
rect 3278 1156 3281 1243
rect 3294 1236 3297 1313
rect 3290 1233 3297 1236
rect 3278 1153 3285 1156
rect 3282 1133 3285 1153
rect 3274 1103 3277 1126
rect 3258 1053 3277 1056
rect 3242 1043 3269 1046
rect 3226 1003 3229 1016
rect 3258 1013 3261 1036
rect 3210 906 3213 926
rect 3218 913 3221 926
rect 3202 903 3213 906
rect 3202 856 3205 903
rect 3202 853 3213 856
rect 3186 823 3189 836
rect 3210 826 3213 853
rect 3194 813 3197 826
rect 3210 823 3221 826
rect 3202 793 3205 806
rect 3170 723 3173 746
rect 3210 736 3213 816
rect 3218 803 3221 823
rect 3226 803 3229 876
rect 3210 733 3221 736
rect 3194 723 3213 726
rect 3162 703 3169 706
rect 3166 636 3169 703
rect 3162 633 3169 636
rect 3178 633 3181 716
rect 3186 703 3189 716
rect 3218 713 3221 733
rect 3226 713 3229 766
rect 3234 696 3237 956
rect 3242 936 3245 1006
rect 3242 933 3253 936
rect 3258 933 3261 946
rect 3266 926 3269 1043
rect 3274 996 3277 1053
rect 3274 993 3281 996
rect 3242 773 3245 926
rect 3254 923 3269 926
rect 3254 866 3257 923
rect 3250 863 3257 866
rect 3242 713 3245 736
rect 3226 693 3237 696
rect 3162 616 3165 633
rect 3226 616 3229 693
rect 3162 613 3173 616
rect 3130 523 3133 596
rect 3150 593 3157 596
rect 3162 593 3165 606
rect 3138 513 3141 586
rect 3150 506 3153 593
rect 3170 586 3173 613
rect 3178 603 3181 616
rect 3226 613 3237 616
rect 3162 583 3173 586
rect 3162 513 3165 583
rect 3178 553 3181 596
rect 3234 593 3237 613
rect 3250 576 3253 863
rect 3258 813 3261 846
rect 3258 693 3261 806
rect 3266 803 3269 916
rect 3278 866 3281 993
rect 3290 936 3293 1233
rect 3298 1106 3301 1136
rect 3306 1113 3309 1316
rect 3322 1286 3325 1353
rect 3362 1336 3365 1456
rect 3354 1333 3365 1336
rect 3322 1283 3333 1286
rect 3330 1216 3333 1283
rect 3322 1213 3333 1216
rect 3322 1193 3325 1213
rect 3322 1123 3325 1136
rect 3330 1123 3333 1156
rect 3338 1123 3349 1126
rect 3298 1103 3317 1106
rect 3298 1003 3301 1026
rect 3290 933 3301 936
rect 3274 863 3281 866
rect 3274 843 3277 863
rect 3274 813 3277 836
rect 3282 793 3285 806
rect 3290 803 3293 926
rect 3298 906 3301 933
rect 3306 923 3309 1016
rect 3298 903 3305 906
rect 3302 806 3305 903
rect 3298 803 3305 806
rect 3298 783 3301 803
rect 3314 793 3317 1103
rect 3354 1046 3357 1333
rect 3370 1296 3373 1526
rect 3382 1466 3385 1543
rect 3394 1476 3397 1593
rect 3402 1543 3405 1556
rect 3418 1533 3421 1576
rect 3442 1573 3445 1606
rect 3450 1593 3453 1616
rect 3394 1473 3401 1476
rect 3382 1463 3389 1466
rect 3378 1403 3381 1446
rect 3386 1393 3389 1463
rect 3398 1426 3401 1473
rect 3394 1423 3401 1426
rect 3394 1403 3397 1423
rect 3410 1413 3413 1446
rect 3442 1433 3445 1526
rect 3458 1503 3461 1606
rect 3466 1523 3469 1633
rect 3482 1626 3485 1703
rect 3498 1703 3509 1706
rect 3498 1656 3501 1703
rect 3514 1663 3517 1726
rect 3530 1723 3537 1726
rect 3546 1723 3549 1896
rect 3562 1856 3565 2023
rect 3562 1853 3569 1856
rect 3566 1776 3569 1853
rect 3578 1813 3581 1936
rect 3586 1906 3589 2126
rect 3594 1933 3597 2136
rect 3602 2116 3605 2173
rect 3610 2133 3613 2156
rect 3602 2113 3609 2116
rect 3606 1946 3609 2113
rect 3618 2106 3621 2136
rect 3642 2123 3645 2233
rect 3650 2193 3653 2206
rect 3658 2203 3661 2216
rect 3674 2206 3677 2406
rect 3690 2403 3693 2416
rect 3674 2203 3685 2206
rect 3618 2103 3629 2106
rect 3626 2036 3629 2103
rect 3618 2033 3629 2036
rect 3618 1993 3621 2033
rect 3650 2003 3653 2066
rect 3658 2023 3661 2036
rect 3666 2023 3669 2136
rect 3674 2096 3677 2126
rect 3682 2113 3685 2203
rect 3690 2173 3693 2386
rect 3714 2306 3717 2633
rect 3722 2563 3725 2746
rect 3746 2686 3749 2726
rect 3738 2683 3749 2686
rect 3730 2596 3733 2616
rect 3738 2603 3741 2683
rect 3746 2613 3749 2626
rect 3754 2613 3757 2753
rect 3762 2676 3765 2796
rect 3770 2723 3773 2736
rect 3762 2673 3773 2676
rect 3762 2613 3765 2666
rect 3770 2613 3773 2673
rect 3730 2593 3741 2596
rect 3722 2523 3725 2536
rect 3722 2393 3725 2416
rect 3730 2383 3733 2586
rect 3738 2533 3741 2593
rect 3754 2553 3757 2606
rect 3754 2423 3757 2536
rect 3778 2513 3781 2616
rect 3794 2566 3797 2823
rect 3802 2813 3813 2816
rect 3794 2563 3801 2566
rect 3786 2523 3789 2556
rect 3798 2516 3801 2563
rect 3794 2513 3801 2516
rect 3818 2513 3821 2873
rect 3842 2816 3845 2883
rect 3834 2813 3845 2816
rect 3834 2743 3837 2813
rect 3842 2733 3845 2796
rect 3866 2736 3869 2913
rect 3890 2786 3893 2943
rect 3898 2933 3909 2936
rect 3906 2823 3909 2926
rect 3922 2796 3925 3046
rect 3938 2983 3941 3036
rect 3922 2793 3929 2796
rect 3890 2783 3917 2786
rect 3858 2733 3869 2736
rect 3858 2716 3861 2733
rect 3850 2713 3861 2716
rect 3850 2636 3853 2713
rect 3842 2633 3853 2636
rect 3834 2603 3837 2626
rect 3842 2576 3845 2633
rect 3850 2613 3861 2616
rect 3866 2613 3869 2646
rect 3858 2576 3861 2606
rect 3842 2573 3853 2576
rect 3858 2573 3869 2576
rect 3738 2313 3741 2326
rect 3706 2303 3717 2306
rect 3674 2093 3681 2096
rect 3658 2003 3661 2016
rect 3666 2003 3669 2016
rect 3678 1996 3681 2093
rect 3690 2013 3693 2136
rect 3706 2096 3709 2303
rect 3794 2226 3797 2513
rect 3818 2413 3821 2436
rect 3834 2406 3837 2556
rect 3850 2413 3853 2573
rect 3866 2526 3869 2573
rect 3874 2553 3877 2746
rect 3890 2733 3901 2736
rect 3882 2686 3885 2726
rect 3890 2703 3893 2726
rect 3906 2713 3909 2726
rect 3914 2696 3917 2783
rect 3926 2706 3929 2793
rect 3906 2693 3917 2696
rect 3922 2703 3929 2706
rect 3882 2683 3893 2686
rect 3890 2626 3893 2683
rect 3882 2623 3893 2626
rect 3882 2603 3885 2623
rect 3906 2606 3909 2693
rect 3922 2613 3925 2703
rect 3930 2673 3933 2686
rect 3906 2603 3917 2606
rect 3890 2533 3901 2536
rect 3866 2523 3877 2526
rect 3882 2513 3885 2526
rect 3834 2403 3845 2406
rect 3810 2323 3813 2356
rect 3818 2306 3821 2366
rect 3842 2333 3845 2403
rect 3810 2303 3821 2306
rect 3810 2236 3813 2303
rect 3810 2233 3821 2236
rect 3786 2223 3797 2226
rect 3730 2193 3733 2216
rect 3722 2123 3725 2176
rect 3706 2093 3725 2096
rect 3706 2003 3709 2016
rect 3674 1993 3681 1996
rect 3602 1943 3609 1946
rect 3586 1903 3593 1906
rect 3590 1836 3593 1903
rect 3586 1833 3593 1836
rect 3586 1813 3589 1833
rect 3562 1773 3569 1776
rect 3498 1653 3509 1656
rect 3474 1623 3485 1626
rect 3474 1603 3477 1623
rect 3506 1613 3509 1653
rect 3482 1523 3485 1596
rect 3490 1533 3493 1556
rect 3498 1523 3501 1606
rect 3506 1593 3517 1596
rect 3514 1543 3517 1593
rect 3522 1583 3525 1716
rect 3534 1656 3537 1723
rect 3562 1716 3565 1773
rect 3530 1653 3537 1656
rect 3554 1713 3565 1716
rect 3530 1573 3533 1653
rect 3538 1516 3541 1636
rect 3546 1613 3549 1626
rect 3554 1603 3557 1713
rect 3570 1673 3573 1736
rect 3586 1733 3589 1806
rect 3602 1753 3605 1943
rect 3610 1906 3613 1926
rect 3650 1923 3653 1936
rect 3674 1913 3677 1993
rect 3698 1933 3701 1946
rect 3722 1943 3725 2093
rect 3786 2066 3789 2223
rect 3818 2216 3821 2233
rect 3802 2203 3805 2216
rect 3810 2213 3821 2216
rect 3810 2196 3813 2213
rect 3810 2193 3821 2196
rect 3802 2183 3813 2186
rect 3802 2096 3805 2176
rect 3802 2093 3813 2096
rect 3786 2063 3793 2066
rect 3746 2013 3749 2026
rect 3790 1976 3793 2063
rect 3810 2023 3813 2093
rect 3818 2016 3821 2193
rect 3826 2163 3829 2306
rect 3874 2216 3877 2496
rect 3898 2473 3901 2526
rect 3906 2456 3909 2516
rect 3914 2493 3917 2603
rect 3938 2536 3941 2956
rect 3970 2953 3973 3113
rect 3994 3066 3997 3163
rect 3994 3063 4005 3066
rect 3986 3003 3989 3016
rect 4002 2966 4005 3063
rect 3994 2963 4005 2966
rect 3946 2683 3949 2766
rect 3954 2753 3957 2936
rect 3962 2883 3965 2936
rect 3994 2866 3997 2963
rect 4010 2876 4013 3183
rect 4034 3123 4037 3146
rect 4042 3106 4045 3186
rect 4034 3103 4045 3106
rect 4034 3036 4037 3103
rect 4050 3036 4053 3206
rect 4058 3143 4061 3366
rect 4090 3296 4093 3376
rect 4082 3293 4093 3296
rect 4082 3206 4085 3293
rect 4114 3276 4117 3326
rect 4098 3273 4117 3276
rect 4090 3213 4093 3226
rect 4074 3203 4085 3206
rect 4074 3086 4077 3203
rect 4074 3083 4085 3086
rect 4034 3033 4045 3036
rect 4050 3033 4069 3036
rect 4034 3006 4037 3016
rect 4018 2933 4021 3006
rect 4026 3003 4037 3006
rect 4026 2923 4029 3003
rect 4042 2996 4045 3033
rect 4034 2993 4045 2996
rect 4034 2886 4037 2993
rect 4050 2896 4053 3006
rect 4050 2893 4057 2896
rect 4026 2883 4037 2886
rect 4010 2873 4021 2876
rect 3994 2863 4005 2866
rect 3962 2733 3965 2806
rect 3978 2743 3981 2806
rect 4002 2786 4005 2863
rect 4010 2803 4013 2816
rect 4018 2796 4021 2873
rect 3998 2783 4005 2786
rect 4010 2793 4021 2796
rect 3970 2733 3981 2736
rect 3954 2646 3957 2726
rect 3970 2723 3989 2726
rect 3986 2676 3989 2723
rect 3998 2696 4001 2783
rect 3998 2693 4005 2696
rect 3986 2673 3997 2676
rect 3950 2643 3957 2646
rect 3950 2596 3953 2643
rect 3962 2603 3965 2626
rect 3950 2593 3957 2596
rect 3930 2533 3941 2536
rect 3930 2486 3933 2533
rect 3954 2526 3957 2593
rect 3970 2583 3973 2616
rect 3978 2613 3989 2616
rect 3994 2603 3997 2673
rect 3898 2453 3909 2456
rect 3922 2483 3933 2486
rect 3950 2523 3957 2526
rect 3898 2376 3901 2453
rect 3898 2373 3909 2376
rect 3906 2356 3909 2373
rect 3922 2366 3925 2483
rect 3938 2403 3941 2446
rect 3950 2436 3953 2523
rect 3946 2433 3953 2436
rect 3922 2363 3933 2366
rect 3906 2353 3913 2356
rect 3890 2313 3893 2326
rect 3910 2286 3913 2353
rect 3906 2283 3913 2286
rect 3842 2213 3861 2216
rect 3834 2146 3837 2206
rect 3850 2173 3853 2206
rect 3858 2203 3861 2213
rect 3866 2213 3877 2216
rect 3866 2203 3869 2213
rect 3874 2193 3877 2206
rect 3834 2143 3845 2146
rect 3842 2123 3845 2143
rect 3790 1973 3797 1976
rect 3714 1913 3717 1926
rect 3610 1903 3621 1906
rect 3618 1826 3621 1903
rect 3746 1843 3749 1936
rect 3778 1933 3781 1946
rect 3786 1933 3789 1956
rect 3794 1933 3797 1973
rect 3802 1943 3805 2016
rect 3810 2013 3821 2016
rect 3810 1996 3813 2013
rect 3810 1993 3821 1996
rect 3794 1903 3797 1926
rect 3610 1823 3621 1826
rect 3610 1803 3613 1823
rect 3714 1813 3717 1836
rect 3810 1833 3813 1966
rect 3818 1943 3821 1993
rect 3826 1896 3829 2016
rect 3850 2013 3853 2166
rect 3882 2123 3885 2216
rect 3890 2173 3893 2276
rect 3898 2163 3901 2246
rect 3906 2106 3909 2283
rect 3922 2243 3925 2326
rect 3922 2203 3925 2226
rect 3930 2213 3933 2363
rect 3938 2323 3941 2336
rect 3946 2303 3949 2433
rect 3962 2413 3965 2526
rect 3978 2516 3981 2536
rect 3974 2513 3981 2516
rect 3974 2436 3977 2513
rect 3974 2433 3981 2436
rect 3978 2413 3981 2433
rect 3986 2406 3989 2596
rect 4002 2466 4005 2693
rect 4010 2576 4013 2793
rect 4026 2716 4029 2883
rect 4042 2743 4045 2886
rect 4054 2836 4057 2893
rect 4050 2833 4057 2836
rect 4050 2773 4053 2833
rect 4066 2826 4069 3033
rect 4074 3003 4077 3076
rect 4082 3036 4085 3083
rect 4090 3043 4093 3206
rect 4098 3203 4101 3273
rect 4126 3266 4129 3383
rect 4142 3376 4145 3443
rect 4166 3376 4169 3453
rect 4138 3373 4145 3376
rect 4162 3373 4169 3376
rect 4138 3276 4141 3373
rect 4138 3273 4149 3276
rect 4126 3263 4133 3266
rect 4106 3156 4109 3236
rect 4114 3213 4117 3226
rect 4098 3153 4109 3156
rect 4114 3153 4117 3206
rect 4130 3173 4133 3263
rect 4146 3166 4149 3273
rect 4142 3163 4149 3166
rect 4082 3033 4089 3036
rect 4086 2946 4089 3033
rect 4086 2943 4093 2946
rect 4082 2906 4085 2926
rect 4078 2903 4085 2906
rect 4078 2846 4081 2903
rect 4078 2843 4085 2846
rect 4066 2823 4073 2826
rect 4058 2766 4061 2816
rect 4070 2766 4073 2823
rect 4082 2803 4085 2843
rect 4090 2803 4093 2943
rect 4050 2763 4061 2766
rect 4066 2763 4073 2766
rect 4018 2713 4029 2716
rect 4018 2673 4021 2713
rect 4034 2696 4037 2726
rect 4042 2713 4045 2736
rect 4050 2733 4053 2763
rect 4058 2733 4061 2746
rect 4066 2723 4069 2763
rect 4074 2733 4077 2746
rect 4082 2723 4085 2756
rect 4090 2703 4093 2736
rect 4098 2733 4101 3153
rect 4106 2973 4109 3056
rect 4114 3033 4117 3146
rect 4142 3096 4145 3163
rect 4154 3123 4157 3146
rect 4138 3093 4145 3096
rect 4138 3026 4141 3093
rect 4162 3086 4165 3373
rect 4170 3306 4173 3326
rect 4178 3323 4181 3426
rect 4186 3333 4189 3416
rect 4170 3303 4181 3306
rect 4178 3226 4181 3303
rect 4194 3273 4197 3406
rect 4202 3396 4205 3493
rect 4218 3413 4221 3446
rect 4226 3403 4229 3526
rect 4234 3443 4237 3673
rect 4242 3613 4245 3736
rect 4254 3646 4257 3743
rect 4250 3643 4257 3646
rect 4250 3566 4253 3643
rect 4250 3563 4257 3566
rect 4254 3486 4257 3563
rect 4250 3483 4257 3486
rect 4250 3426 4253 3483
rect 4250 3423 4257 3426
rect 4234 3413 4245 3416
rect 4202 3393 4213 3396
rect 4210 3376 4213 3393
rect 4242 3383 4245 3406
rect 4254 3376 4257 3423
rect 4210 3373 4221 3376
rect 4218 3266 4221 3373
rect 4250 3373 4257 3376
rect 4250 3356 4253 3373
rect 4170 3223 4181 3226
rect 4210 3263 4221 3266
rect 4242 3353 4253 3356
rect 4170 3203 4173 3223
rect 4194 3123 4197 3206
rect 4202 3106 4205 3176
rect 4210 3163 4213 3263
rect 4194 3103 4205 3106
rect 4162 3083 4173 3086
rect 4118 3023 4141 3026
rect 4106 2726 4109 2866
rect 4118 2766 4121 3023
rect 4130 2993 4133 3016
rect 4146 3013 4165 3016
rect 4130 2813 4133 2946
rect 4138 2923 4141 3006
rect 4146 2943 4149 3013
rect 4154 2983 4157 3006
rect 4162 3003 4165 3013
rect 4170 3006 4173 3083
rect 4178 3013 4181 3056
rect 4194 3036 4197 3103
rect 4194 3033 4205 3036
rect 4186 3013 4197 3016
rect 4202 3006 4205 3033
rect 4170 3003 4181 3006
rect 4162 2913 4165 2936
rect 4178 2846 4181 3003
rect 4198 3003 4205 3006
rect 4186 2933 4189 2976
rect 4198 2926 4201 3003
rect 4210 2973 4213 3156
rect 4218 3116 4221 3206
rect 4226 3193 4229 3216
rect 4234 3186 4237 3216
rect 4242 3213 4245 3353
rect 4258 3333 4261 3356
rect 4226 3183 4237 3186
rect 4226 3133 4229 3183
rect 4242 3173 4245 3206
rect 4250 3123 4253 3196
rect 4258 3153 4261 3216
rect 4266 3203 4269 3833
rect 4274 3813 4277 3826
rect 4282 3803 4285 3816
rect 4298 3736 4301 3833
rect 4306 3796 4309 3816
rect 4306 3793 4317 3796
rect 4290 3733 4301 3736
rect 4274 3706 4277 3726
rect 4274 3703 4281 3706
rect 4278 3626 4281 3703
rect 4274 3623 4281 3626
rect 4290 3623 4293 3733
rect 4314 3726 4317 3793
rect 4306 3723 4317 3726
rect 4274 3603 4277 3623
rect 4290 3583 4293 3616
rect 4274 3533 4293 3536
rect 4274 3363 4277 3533
rect 4282 3413 4285 3526
rect 4290 3513 4293 3526
rect 4306 3436 4309 3723
rect 4322 3523 4325 3616
rect 4330 3543 4333 3826
rect 4338 3823 4349 3826
rect 4346 3753 4349 3816
rect 4346 3716 4349 3736
rect 4342 3713 4349 3716
rect 4342 3636 4345 3713
rect 4358 3706 4361 3853
rect 4370 3786 4373 4026
rect 4378 4023 4381 4036
rect 4378 4003 4381 4016
rect 4386 3996 4389 4043
rect 4394 4013 4397 4126
rect 4402 4116 4405 4133
rect 4402 4113 4409 4116
rect 4406 4046 4409 4113
rect 4402 4043 4409 4046
rect 4402 4023 4405 4043
rect 4378 3993 4389 3996
rect 4378 3906 4381 3993
rect 4394 3933 4397 3966
rect 4418 3936 4421 4133
rect 4434 3963 4437 4153
rect 4458 4123 4461 4146
rect 4470 4116 4473 4163
rect 4538 4146 4541 4213
rect 4538 4143 4549 4146
rect 4466 4113 4473 4116
rect 4450 4003 4453 4026
rect 4418 3933 4437 3936
rect 4418 3913 4421 3926
rect 4378 3903 4389 3906
rect 4386 3803 4389 3903
rect 4434 3856 4437 3933
rect 4466 3923 4469 4113
rect 4514 4023 4517 4126
rect 4538 4026 4541 4126
rect 4546 4036 4549 4143
rect 4554 4093 4557 4216
rect 4562 4213 4573 4216
rect 4562 4193 4565 4206
rect 4578 4203 4581 4223
rect 4594 4213 4597 4316
rect 4602 4313 4613 4316
rect 4610 4266 4613 4313
rect 4602 4263 4613 4266
rect 4642 4266 4645 4383
rect 4642 4263 4653 4266
rect 4562 4113 4565 4136
rect 4570 4103 4573 4126
rect 4546 4033 4565 4036
rect 4538 4023 4549 4026
rect 4514 3993 4517 4016
rect 4546 4006 4549 4023
rect 4554 4013 4557 4026
rect 4546 4003 4557 4006
rect 4430 3853 4437 3856
rect 4370 3783 4381 3786
rect 4378 3736 4381 3783
rect 4418 3763 4421 3816
rect 4430 3776 4433 3853
rect 4430 3773 4437 3776
rect 4378 3733 4389 3736
rect 4354 3703 4361 3706
rect 4342 3633 4349 3636
rect 4338 3593 4341 3606
rect 4346 3603 4349 3633
rect 4354 3613 4357 3703
rect 4330 3533 4341 3536
rect 4346 3533 4349 3566
rect 4354 3526 4357 3606
rect 4362 3603 4365 3626
rect 4370 3593 4373 3726
rect 4386 3666 4389 3733
rect 4434 3716 4437 3773
rect 4466 3736 4469 3816
rect 4442 3723 4445 3736
rect 4450 3733 4469 3736
rect 4474 3733 4477 3956
rect 4490 3923 4493 3936
rect 4498 3933 4501 3976
rect 4554 3953 4557 4003
rect 4498 3776 4501 3926
rect 4514 3793 4517 3926
rect 4538 3923 4541 3946
rect 4562 3943 4565 4033
rect 4578 4013 4581 4136
rect 4586 4133 4589 4206
rect 4594 4123 4597 4136
rect 4602 4106 4605 4263
rect 4642 4213 4645 4226
rect 4618 4183 4621 4206
rect 4634 4126 4637 4156
rect 4650 4153 4653 4263
rect 4666 4256 4669 4406
rect 4690 4393 4693 4416
rect 4662 4253 4669 4256
rect 4662 4206 4665 4253
rect 4682 4216 4685 4336
rect 4698 4223 4701 4526
rect 4722 4513 4725 4526
rect 4682 4213 4701 4216
rect 4662 4203 4669 4206
rect 4666 4183 4669 4203
rect 4642 4133 4645 4146
rect 4594 4103 4605 4106
rect 4594 4036 4597 4103
rect 4594 4033 4605 4036
rect 4570 3993 4573 4006
rect 4586 3936 4589 4006
rect 4546 3813 4549 3936
rect 4578 3933 4589 3936
rect 4554 3923 4573 3926
rect 4578 3856 4581 3933
rect 4578 3853 4585 3856
rect 4490 3773 4501 3776
rect 4434 3713 4445 3716
rect 4378 3663 4389 3666
rect 4378 3563 4381 3663
rect 4442 3656 4445 3713
rect 4434 3653 4445 3656
rect 4418 3613 4421 3626
rect 4378 3533 4381 3556
rect 4394 3553 4397 3606
rect 4434 3576 4437 3653
rect 4474 3613 4477 3726
rect 4482 3713 4485 3726
rect 4482 3603 4485 3616
rect 4490 3583 4493 3773
rect 4498 3733 4501 3766
rect 4506 3713 4509 3726
rect 4514 3603 4517 3706
rect 4522 3613 4525 3626
rect 4434 3573 4445 3576
rect 4442 3556 4445 3573
rect 4442 3553 4449 3556
rect 4338 3503 4341 3526
rect 4346 3523 4357 3526
rect 4402 3523 4405 3536
rect 4298 3433 4309 3436
rect 4298 3336 4301 3433
rect 4282 3333 4293 3336
rect 4298 3333 4309 3336
rect 4314 3333 4317 3416
rect 4322 3403 4325 3416
rect 4274 3293 4277 3326
rect 4274 3193 4277 3206
rect 4258 3133 4261 3146
rect 4274 3133 4277 3186
rect 4282 3133 4285 3156
rect 4218 3113 4229 3116
rect 4226 3046 4229 3113
rect 4266 3083 4269 3126
rect 4218 3043 4229 3046
rect 4194 2923 4201 2926
rect 4178 2843 4185 2846
rect 4098 2723 4109 2726
rect 4114 2763 4121 2766
rect 4034 2693 4045 2696
rect 4026 2603 4029 2686
rect 4042 2616 4045 2693
rect 4034 2613 4045 2616
rect 4034 2593 4037 2613
rect 4058 2583 4061 2616
rect 4074 2613 4077 2626
rect 4066 2603 4077 2606
rect 4010 2573 4021 2576
rect 3954 2393 3957 2406
rect 3978 2403 3989 2406
rect 3998 2463 4005 2466
rect 3962 2313 3965 2336
rect 3938 2203 3941 2286
rect 3946 2213 3957 2216
rect 3962 2203 3965 2246
rect 3970 2213 3973 2326
rect 3978 2273 3981 2403
rect 3986 2323 3989 2336
rect 3998 2306 4001 2463
rect 4018 2376 4021 2573
rect 3994 2303 4001 2306
rect 4010 2373 4021 2376
rect 3994 2236 3997 2303
rect 3994 2233 4005 2236
rect 3986 2213 3997 2216
rect 3914 2123 3917 2196
rect 3938 2176 3941 2196
rect 3986 2183 3989 2213
rect 3938 2173 3949 2176
rect 3898 2103 3909 2106
rect 3858 2006 3861 2046
rect 3874 2013 3877 2026
rect 3898 2013 3901 2103
rect 3834 1933 3837 2006
rect 3850 2003 3861 2006
rect 3850 1993 3853 2003
rect 3898 1966 3901 2006
rect 3906 2003 3909 2016
rect 3914 2013 3917 2036
rect 3922 1993 3925 2156
rect 3930 2023 3933 2126
rect 3946 2106 3949 2173
rect 3938 2103 3949 2106
rect 3938 2016 3941 2103
rect 3930 2013 3941 2016
rect 3890 1963 3901 1966
rect 3930 1963 3933 2013
rect 3946 2003 3949 2086
rect 3970 2076 3973 2136
rect 3986 2133 3989 2176
rect 3994 2163 3997 2206
rect 4002 2143 4005 2233
rect 3978 2123 3997 2126
rect 4010 2123 4013 2373
rect 4018 2333 4021 2346
rect 4026 2283 4029 2406
rect 4034 2393 4037 2416
rect 4042 2333 4045 2536
rect 4066 2393 4069 2576
rect 4082 2533 4085 2676
rect 4090 2613 4093 2626
rect 4026 2216 4029 2226
rect 4026 2213 4045 2216
rect 4058 2206 4061 2336
rect 4082 2323 4085 2406
rect 4090 2403 4093 2416
rect 4098 2313 4101 2723
rect 4114 2593 4117 2763
rect 4130 2573 4133 2806
rect 4154 2803 4157 2826
rect 4182 2786 4185 2843
rect 4178 2783 4185 2786
rect 4178 2766 4181 2783
rect 4170 2763 4181 2766
rect 4194 2766 4197 2923
rect 4210 2903 4213 2966
rect 4218 2953 4221 3043
rect 4234 3013 4237 3026
rect 4218 2866 4221 2936
rect 4226 2923 4229 3006
rect 4234 2923 4237 2946
rect 4242 2876 4245 2936
rect 4250 2923 4253 2936
rect 4258 2896 4261 3016
rect 4202 2863 4221 2866
rect 4234 2873 4245 2876
rect 4250 2893 4261 2896
rect 4202 2813 4205 2863
rect 4234 2813 4237 2873
rect 4194 2763 4205 2766
rect 4154 2723 4157 2746
rect 4170 2686 4173 2763
rect 4202 2706 4205 2763
rect 4234 2726 4237 2756
rect 4234 2723 4245 2726
rect 4194 2703 4205 2706
rect 4114 2523 4117 2536
rect 4122 2446 4125 2536
rect 4114 2443 4125 2446
rect 4114 2413 4117 2443
rect 4130 2423 4133 2536
rect 4138 2513 4141 2586
rect 4146 2443 4149 2686
rect 4170 2683 4181 2686
rect 4194 2683 4197 2703
rect 4178 2663 4181 2683
rect 4250 2673 4253 2893
rect 4266 2876 4269 2956
rect 4262 2873 4269 2876
rect 4262 2816 4265 2873
rect 4274 2823 4277 3126
rect 4290 3003 4293 3326
rect 4306 3213 4309 3333
rect 4322 3263 4325 3316
rect 4330 3303 4333 3396
rect 4338 3333 4341 3346
rect 4306 2996 4309 3166
rect 4322 3103 4325 3136
rect 4330 3123 4341 3126
rect 4346 3123 4349 3523
rect 4426 3506 4429 3546
rect 4362 3313 4365 3416
rect 4370 3403 4373 3506
rect 4418 3503 4429 3506
rect 4378 3403 4381 3416
rect 4370 3333 4373 3366
rect 4418 3356 4421 3503
rect 4446 3486 4449 3553
rect 4458 3506 4461 3526
rect 4458 3503 4469 3506
rect 4442 3483 4449 3486
rect 4418 3353 4429 3356
rect 4370 3126 4373 3306
rect 4378 3133 4381 3156
rect 4338 3113 4341 3123
rect 4354 3083 4357 3126
rect 4370 3123 4381 3126
rect 4322 3013 4325 3026
rect 4338 3013 4341 3046
rect 4294 2993 4309 2996
rect 4282 2933 4285 2976
rect 4294 2886 4297 2993
rect 4306 2903 4309 2926
rect 4294 2883 4301 2886
rect 4282 2833 4285 2876
rect 4262 2813 4269 2816
rect 4242 2623 4245 2666
rect 4266 2646 4269 2813
rect 4282 2813 4293 2816
rect 4282 2803 4285 2813
rect 4298 2806 4301 2883
rect 4314 2833 4317 2936
rect 4322 2923 4325 3006
rect 4330 2933 4333 2946
rect 4346 2926 4349 3036
rect 4354 3013 4357 3056
rect 4362 2993 4365 3016
rect 4330 2923 4349 2926
rect 4354 2923 4357 2936
rect 4330 2836 4333 2923
rect 4378 2916 4381 3123
rect 4386 3113 4389 3146
rect 4394 3123 4397 3326
rect 4402 3323 4405 3336
rect 4410 3323 4413 3336
rect 4418 3306 4421 3336
rect 4410 3303 4421 3306
rect 4410 3236 4413 3303
rect 4426 3246 4429 3353
rect 4442 3303 4445 3483
rect 4466 3436 4469 3503
rect 4458 3433 4469 3436
rect 4458 3416 4461 3433
rect 4450 3413 4461 3416
rect 4458 3356 4461 3406
rect 4466 3393 4469 3406
rect 4450 3353 4461 3356
rect 4426 3243 4437 3246
rect 4410 3233 4421 3236
rect 4402 3133 4405 3146
rect 4418 3133 4421 3233
rect 4434 3126 4437 3243
rect 4450 3156 4453 3353
rect 4474 3343 4477 3416
rect 4482 3323 4485 3336
rect 4490 3313 4493 3576
rect 4498 3533 4501 3556
rect 4514 3533 4517 3546
rect 4506 3413 4509 3526
rect 4522 3523 4525 3586
rect 4530 3553 4533 3776
rect 4538 3713 4541 3736
rect 4546 3683 4549 3746
rect 4554 3646 4557 3806
rect 4582 3796 4585 3853
rect 4594 3803 4597 4016
rect 4602 4003 4605 4033
rect 4610 4013 4613 4126
rect 4626 4123 4637 4126
rect 4626 4026 4629 4123
rect 4650 4113 4653 4126
rect 4622 4023 4629 4026
rect 4602 3906 4605 3936
rect 4610 3923 4613 4006
rect 4622 3956 4625 4023
rect 4650 4016 4653 4096
rect 4634 4003 4637 4016
rect 4642 4013 4653 4016
rect 4622 3953 4629 3956
rect 4602 3903 4609 3906
rect 4606 3836 4609 3903
rect 4602 3833 4609 3836
rect 4602 3813 4605 3833
rect 4610 3803 4613 3816
rect 4578 3793 4585 3796
rect 4578 3773 4581 3793
rect 4562 3723 4565 3756
rect 4578 3733 4581 3766
rect 4578 3646 4581 3726
rect 4550 3643 4557 3646
rect 4570 3643 4581 3646
rect 4538 3556 4541 3616
rect 4550 3596 4553 3643
rect 4562 3606 4565 3636
rect 4570 3613 4573 3643
rect 4586 3613 4589 3646
rect 4594 3633 4597 3796
rect 4618 3736 4621 3936
rect 4626 3926 4629 3953
rect 4634 3933 4637 3976
rect 4642 3933 4645 4013
rect 4650 3956 4653 4006
rect 4658 4003 4661 4026
rect 4666 4013 4669 4036
rect 4674 4026 4677 4166
rect 4674 4023 4685 4026
rect 4674 3993 4677 4016
rect 4650 3953 4661 3956
rect 4650 3933 4653 3946
rect 4626 3923 4637 3926
rect 4658 3923 4661 3953
rect 4634 3906 4637 3923
rect 4634 3903 4645 3906
rect 4642 3836 4645 3903
rect 4634 3833 4645 3836
rect 4626 3743 4629 3806
rect 4618 3733 4629 3736
rect 4618 3703 4621 3726
rect 4626 3696 4629 3733
rect 4618 3693 4629 3696
rect 4562 3603 4573 3606
rect 4578 3603 4589 3606
rect 4594 3603 4597 3626
rect 4550 3593 4557 3596
rect 4554 3573 4557 3593
rect 4538 3553 4549 3556
rect 4530 3506 4533 3526
rect 4522 3503 4533 3506
rect 4522 3386 4525 3503
rect 4546 3496 4549 3553
rect 4570 3533 4573 3603
rect 4594 3523 4597 3546
rect 4538 3493 4549 3496
rect 4522 3383 4533 3386
rect 4530 3363 4533 3383
rect 4498 3333 4501 3346
rect 4514 3213 4517 3326
rect 4530 3296 4533 3316
rect 4526 3293 4533 3296
rect 4410 3103 4413 3126
rect 4426 3123 4437 3126
rect 4446 3153 4453 3156
rect 4426 3033 4429 3123
rect 4446 3096 4449 3153
rect 4446 3093 4453 3096
rect 4450 3073 4453 3093
rect 4466 3026 4469 3166
rect 4490 3163 4493 3206
rect 4526 3176 4529 3293
rect 4526 3173 4533 3176
rect 4530 3146 4533 3173
rect 4538 3166 4541 3493
rect 4602 3456 4605 3686
rect 4610 3613 4613 3626
rect 4618 3566 4621 3693
rect 4626 3606 4629 3686
rect 4634 3613 4637 3833
rect 4642 3793 4645 3806
rect 4650 3763 4653 3816
rect 4642 3683 4645 3746
rect 4666 3723 4669 3936
rect 4682 3933 4685 4023
rect 4698 3766 4701 4206
rect 4706 4173 4709 4236
rect 4714 4153 4717 4216
rect 4722 4203 4725 4326
rect 4730 4213 4741 4216
rect 4722 4123 4725 4146
rect 4722 3923 4725 3946
rect 4722 3793 4725 3816
rect 4690 3763 4701 3766
rect 4626 3603 4637 3606
rect 4642 3603 4645 3626
rect 4650 3603 4653 3616
rect 4614 3563 4621 3566
rect 4634 3566 4637 3603
rect 4634 3563 4641 3566
rect 4614 3466 4617 3563
rect 4638 3506 4641 3563
rect 4658 3536 4661 3616
rect 4666 3603 4669 3716
rect 4674 3623 4677 3726
rect 4690 3636 4693 3763
rect 4730 3736 4733 4176
rect 4738 4163 4741 4206
rect 4746 4113 4749 4216
rect 4754 4163 4757 4206
rect 4762 4193 4765 4216
rect 4770 4183 4773 4536
rect 4778 4413 4781 4426
rect 4778 4306 4781 4326
rect 4778 4303 4789 4306
rect 4786 4226 4789 4303
rect 4778 4223 4789 4226
rect 4778 4203 4781 4223
rect 4778 4123 4781 4166
rect 4762 3936 4765 3956
rect 4762 3933 4769 3936
rect 4766 3886 4769 3933
rect 4778 3923 4781 4006
rect 4794 3906 4797 3976
rect 4762 3883 4769 3886
rect 4786 3903 4797 3906
rect 4762 3856 4765 3883
rect 4762 3853 4769 3856
rect 4766 3776 4769 3853
rect 4786 3836 4789 3903
rect 4786 3833 4797 3836
rect 4762 3773 4769 3776
rect 4762 3736 4765 3773
rect 4726 3733 4733 3736
rect 4758 3733 4765 3736
rect 4778 3733 4781 3816
rect 4794 3776 4797 3833
rect 4794 3773 4801 3776
rect 4714 3713 4717 3726
rect 4726 3686 4729 3733
rect 4722 3683 4729 3686
rect 4690 3633 4701 3636
rect 4674 3613 4693 3616
rect 4674 3603 4677 3613
rect 4658 3533 4669 3536
rect 4698 3533 4701 3633
rect 4722 3576 4725 3683
rect 4738 3586 4741 3726
rect 4758 3676 4761 3733
rect 4754 3673 4761 3676
rect 4754 3596 4757 3673
rect 4770 3603 4773 3726
rect 4786 3723 4789 3766
rect 4798 3716 4801 3773
rect 4794 3713 4801 3716
rect 4754 3593 4765 3596
rect 4738 3583 4745 3586
rect 4722 3573 4733 3576
rect 4634 3503 4641 3506
rect 4634 3486 4637 3503
rect 4626 3483 4637 3486
rect 4614 3463 4621 3466
rect 4594 3453 4605 3456
rect 4554 3383 4557 3406
rect 4578 3396 4581 3416
rect 4570 3393 4581 3396
rect 4546 3323 4549 3336
rect 4554 3333 4557 3366
rect 4570 3333 4573 3393
rect 4594 3376 4597 3453
rect 4594 3373 4605 3376
rect 4578 3326 4581 3356
rect 4562 3313 4565 3326
rect 4570 3296 4573 3326
rect 4578 3323 4597 3326
rect 4602 3316 4605 3373
rect 4610 3323 4613 3336
rect 4562 3293 4573 3296
rect 4562 3236 4565 3293
rect 4562 3233 4573 3236
rect 4570 3213 4573 3233
rect 4538 3163 4549 3166
rect 4490 3123 4493 3146
rect 4530 3143 4537 3146
rect 4410 3013 4413 3026
rect 4458 3023 4469 3026
rect 4426 3013 4445 3016
rect 4394 2993 4397 3006
rect 4402 2973 4405 3006
rect 4386 2923 4389 2936
rect 4378 2913 4389 2916
rect 4402 2913 4405 2956
rect 4418 2946 4421 3006
rect 4426 2993 4429 3013
rect 4434 2983 4437 3006
rect 4458 2976 4461 3023
rect 4458 2973 4469 2976
rect 4418 2943 4429 2946
rect 4426 2923 4429 2943
rect 4326 2833 4333 2836
rect 4290 2803 4301 2806
rect 4290 2723 4293 2803
rect 4314 2723 4317 2826
rect 4326 2786 4329 2833
rect 4346 2803 4349 2856
rect 4370 2813 4373 2836
rect 4326 2783 4333 2786
rect 4262 2643 4269 2646
rect 4250 2623 4253 2636
rect 4178 2603 4181 2616
rect 4178 2566 4181 2596
rect 4226 2566 4229 2616
rect 4170 2563 4181 2566
rect 4170 2506 4173 2563
rect 4194 2533 4197 2566
rect 4218 2563 4229 2566
rect 4218 2546 4221 2563
rect 4218 2543 4229 2546
rect 4170 2503 4181 2506
rect 4170 2413 4173 2426
rect 4114 2323 4117 2346
rect 4018 2203 4029 2206
rect 4058 2203 4069 2206
rect 4114 2203 4117 2216
rect 3978 2083 3981 2123
rect 3970 2073 3989 2076
rect 4026 2073 4029 2136
rect 3986 2013 3989 2073
rect 4034 2043 4037 2146
rect 4050 2133 4061 2136
rect 4042 2086 4045 2126
rect 4042 2083 4053 2086
rect 3850 1933 3853 1946
rect 3874 1923 3877 1936
rect 3826 1893 3837 1896
rect 3834 1846 3837 1893
rect 3890 1886 3893 1963
rect 3962 1943 3965 2006
rect 4034 2003 4037 2026
rect 4042 2013 4045 2076
rect 4050 2013 4053 2083
rect 4050 1993 4053 2006
rect 4058 1953 4061 2126
rect 4066 2116 4069 2203
rect 4162 2166 4165 2336
rect 4178 2283 4181 2503
rect 4226 2496 4229 2543
rect 4242 2523 4245 2546
rect 4262 2526 4265 2643
rect 4298 2636 4301 2716
rect 4330 2713 4333 2783
rect 4346 2723 4349 2776
rect 4386 2733 4389 2913
rect 4426 2876 4429 2916
rect 4418 2873 4429 2876
rect 4418 2816 4421 2873
rect 4418 2813 4429 2816
rect 4434 2813 4437 2926
rect 4466 2913 4469 2973
rect 4442 2813 4445 2906
rect 4474 2903 4477 3016
rect 4482 2923 4485 3006
rect 4426 2796 4429 2813
rect 4306 2693 4309 2706
rect 4362 2693 4365 2726
rect 4274 2613 4277 2636
rect 4290 2633 4301 2636
rect 4262 2523 4269 2526
rect 4274 2523 4277 2586
rect 4290 2556 4293 2633
rect 4306 2616 4309 2626
rect 4338 2623 4341 2636
rect 4346 2633 4349 2656
rect 4306 2613 4317 2616
rect 4306 2583 4309 2606
rect 4314 2596 4317 2613
rect 4314 2593 4321 2596
rect 4290 2553 4301 2556
rect 4282 2533 4293 2536
rect 4218 2493 4229 2496
rect 4194 2323 4197 2336
rect 4218 2323 4221 2493
rect 4242 2413 4245 2516
rect 4266 2506 4269 2523
rect 4282 2513 4285 2526
rect 4266 2503 4277 2506
rect 4274 2446 4277 2503
rect 4274 2443 4285 2446
rect 4258 2413 4261 2426
rect 4234 2353 4237 2406
rect 4250 2366 4253 2406
rect 4266 2403 4269 2416
rect 4274 2413 4277 2426
rect 4242 2363 4253 2366
rect 4242 2323 4245 2363
rect 4274 2323 4277 2406
rect 4282 2313 4285 2443
rect 4290 2413 4293 2533
rect 4298 2506 4301 2553
rect 4306 2523 4309 2536
rect 4318 2516 4321 2593
rect 4330 2523 4333 2616
rect 4354 2613 4357 2626
rect 4354 2603 4373 2606
rect 4338 2533 4341 2546
rect 4354 2533 4357 2603
rect 4362 2533 4365 2556
rect 4314 2513 4321 2516
rect 4346 2513 4349 2526
rect 4298 2503 4305 2506
rect 4302 2406 4305 2503
rect 4298 2403 4305 2406
rect 4314 2403 4317 2513
rect 4338 2433 4341 2466
rect 4298 2346 4301 2403
rect 4294 2343 4301 2346
rect 4282 2293 4285 2306
rect 4226 2233 4237 2236
rect 4226 2193 4229 2226
rect 4250 2223 4253 2286
rect 4294 2276 4297 2343
rect 4322 2336 4325 2426
rect 4306 2333 4325 2336
rect 4338 2333 4341 2426
rect 4346 2413 4349 2436
rect 4306 2323 4309 2333
rect 4290 2273 4297 2276
rect 4290 2196 4293 2273
rect 4306 2233 4309 2316
rect 4322 2223 4349 2226
rect 4306 2203 4309 2216
rect 4330 2213 4341 2216
rect 4346 2213 4349 2223
rect 4354 2213 4357 2416
rect 4362 2376 4365 2426
rect 4378 2413 4381 2726
rect 4402 2653 4405 2766
rect 4410 2696 4413 2746
rect 4418 2723 4421 2796
rect 4426 2793 4445 2796
rect 4434 2773 4437 2786
rect 4442 2696 4445 2793
rect 4450 2783 4453 2816
rect 4466 2813 4485 2816
rect 4490 2813 4493 3036
rect 4498 3003 4501 3116
rect 4534 3076 4537 3143
rect 4530 3073 4537 3076
rect 4530 3053 4533 3073
rect 4546 3056 4549 3163
rect 4570 3103 4573 3126
rect 4578 3123 4581 3316
rect 4602 3313 4613 3316
rect 4586 3286 4589 3306
rect 4586 3283 4597 3286
rect 4594 3226 4597 3283
rect 4586 3223 4597 3226
rect 4586 3086 4589 3223
rect 4594 3183 4597 3206
rect 4594 3113 4597 3136
rect 4538 3053 4549 3056
rect 4578 3083 4589 3086
rect 4538 3033 4541 3053
rect 4578 3036 4581 3083
rect 4578 3033 4589 3036
rect 4538 3013 4557 3016
rect 4458 2746 4461 2806
rect 4474 2793 4477 2806
rect 4482 2803 4485 2813
rect 4506 2766 4509 2936
rect 4530 2923 4533 3006
rect 4546 2926 4549 3006
rect 4554 3003 4557 3013
rect 4546 2923 4553 2926
rect 4506 2763 4513 2766
rect 4458 2743 4469 2746
rect 4466 2723 4469 2743
rect 4510 2716 4513 2763
rect 4522 2726 4525 2806
rect 4530 2803 4533 2816
rect 4538 2803 4541 2916
rect 4550 2856 4553 2923
rect 4546 2853 4553 2856
rect 4546 2793 4549 2853
rect 4586 2836 4589 3033
rect 4602 3013 4605 3126
rect 4594 2993 4597 3006
rect 4610 2976 4613 3313
rect 4618 3303 4621 3463
rect 4626 3203 4629 3483
rect 4634 3333 4637 3416
rect 4642 3413 4645 3426
rect 4650 3403 4653 3526
rect 4666 3436 4669 3533
rect 4658 3433 4669 3436
rect 4658 3413 4661 3433
rect 4658 3363 4661 3406
rect 4682 3403 4685 3516
rect 4722 3513 4725 3526
rect 4730 3486 4733 3573
rect 4722 3483 4733 3486
rect 4690 3413 4709 3416
rect 4690 3393 4693 3413
rect 4722 3396 4725 3483
rect 4742 3476 4745 3583
rect 4762 3576 4765 3593
rect 4762 3573 4769 3576
rect 4766 3486 4769 3573
rect 4738 3473 4745 3476
rect 4762 3483 4769 3486
rect 4738 3403 4741 3473
rect 4722 3393 4733 3396
rect 4634 3306 4637 3326
rect 4634 3303 4645 3306
rect 4642 3226 4645 3303
rect 4634 3223 4645 3226
rect 4618 3133 4621 3146
rect 4626 3123 4629 3156
rect 4602 2973 4613 2976
rect 4602 2856 4605 2973
rect 4602 2853 4609 2856
rect 4554 2813 4557 2836
rect 4586 2833 4597 2836
rect 4562 2813 4573 2816
rect 4522 2723 4541 2726
rect 4510 2713 4525 2716
rect 4410 2693 4421 2696
rect 4418 2636 4421 2693
rect 4410 2633 4421 2636
rect 4434 2693 4445 2696
rect 4434 2636 4437 2693
rect 4434 2633 4445 2636
rect 4402 2606 4405 2626
rect 4394 2603 4405 2606
rect 4394 2546 4397 2603
rect 4394 2543 4405 2546
rect 4402 2523 4405 2543
rect 4410 2533 4413 2633
rect 4418 2506 4421 2526
rect 4410 2503 4421 2506
rect 4378 2393 4381 2406
rect 4410 2376 4413 2503
rect 4426 2413 4429 2606
rect 4434 2543 4437 2616
rect 4442 2613 4445 2633
rect 4450 2603 4453 2656
rect 4466 2613 4469 2696
rect 4490 2603 4493 2616
rect 4506 2586 4509 2676
rect 4498 2583 4509 2586
rect 4442 2456 4445 2536
rect 4442 2453 4449 2456
rect 4446 2396 4449 2453
rect 4458 2413 4461 2536
rect 4466 2533 4469 2546
rect 4498 2466 4501 2583
rect 4498 2463 4509 2466
rect 4474 2403 4477 2446
rect 4442 2393 4449 2396
rect 4442 2376 4445 2393
rect 4362 2373 4389 2376
rect 4386 2323 4389 2373
rect 4402 2373 4413 2376
rect 4426 2373 4445 2376
rect 4402 2316 4405 2373
rect 4362 2293 4365 2316
rect 4378 2313 4405 2316
rect 4410 2313 4413 2336
rect 4418 2333 4421 2356
rect 4426 2326 4429 2373
rect 4434 2333 4437 2346
rect 4418 2323 4429 2326
rect 4378 2213 4381 2313
rect 4418 2306 4421 2323
rect 4442 2313 4445 2326
rect 4410 2303 4421 2306
rect 4290 2193 4301 2196
rect 4154 2163 4165 2166
rect 4066 2113 4077 2116
rect 4074 2046 4077 2113
rect 4154 2053 4157 2163
rect 4178 2123 4181 2136
rect 4258 2133 4261 2146
rect 4250 2113 4253 2126
rect 4298 2056 4301 2193
rect 4066 2043 4077 2046
rect 4066 2023 4069 2043
rect 4066 2013 4093 2016
rect 4066 1993 4069 2006
rect 4074 2003 4085 2006
rect 4162 1993 4165 2016
rect 4210 1993 4213 2056
rect 4298 2053 4309 2056
rect 4282 2013 4285 2026
rect 4234 1993 4237 2006
rect 4306 1976 4309 2053
rect 4330 2013 4333 2206
rect 4362 2113 4365 2126
rect 4370 2023 4373 2136
rect 4386 2133 4389 2216
rect 4394 2203 4397 2226
rect 4410 2213 4413 2303
rect 4450 2296 4453 2336
rect 4442 2293 4453 2296
rect 4442 2226 4445 2293
rect 4426 2213 4429 2226
rect 4442 2223 4453 2226
rect 4378 2103 4381 2126
rect 4298 1973 4309 1976
rect 4298 1956 4301 1973
rect 4294 1953 4301 1956
rect 3890 1883 3901 1886
rect 3826 1843 3837 1846
rect 3626 1746 3629 1806
rect 3626 1743 3637 1746
rect 3602 1633 3605 1736
rect 3634 1696 3637 1743
rect 3650 1723 3653 1736
rect 3626 1693 3637 1696
rect 3626 1653 3629 1693
rect 3554 1593 3565 1596
rect 3534 1513 3541 1516
rect 3402 1403 3413 1406
rect 3378 1333 3381 1356
rect 3386 1343 3389 1366
rect 3418 1353 3421 1416
rect 3522 1413 3525 1466
rect 3534 1456 3537 1513
rect 3534 1453 3541 1456
rect 3506 1383 3509 1396
rect 3514 1393 3517 1406
rect 3530 1383 3533 1436
rect 3474 1296 3477 1326
rect 3370 1293 3381 1296
rect 3378 1166 3381 1293
rect 3458 1293 3477 1296
rect 3458 1206 3461 1293
rect 3482 1213 3485 1376
rect 3490 1323 3493 1356
rect 3522 1256 3525 1346
rect 3538 1343 3541 1453
rect 3546 1403 3549 1506
rect 3554 1413 3557 1516
rect 3570 1453 3573 1586
rect 3578 1513 3581 1526
rect 3586 1433 3589 1596
rect 3610 1433 3613 1576
rect 3650 1446 3653 1616
rect 3658 1613 3661 1626
rect 3666 1543 3669 1746
rect 3730 1716 3733 1816
rect 3746 1803 3749 1826
rect 3754 1773 3757 1806
rect 3770 1793 3773 1806
rect 3778 1766 3781 1816
rect 3794 1813 3797 1826
rect 3826 1823 3829 1843
rect 3762 1763 3781 1766
rect 3738 1733 3741 1756
rect 3746 1733 3757 1736
rect 3674 1536 3677 1616
rect 3706 1613 3709 1636
rect 3682 1593 3685 1606
rect 3666 1533 3677 1536
rect 3650 1443 3661 1446
rect 3562 1393 3565 1416
rect 3650 1393 3653 1416
rect 3658 1403 3661 1443
rect 3666 1423 3669 1533
rect 3546 1346 3549 1366
rect 3546 1343 3553 1346
rect 3550 1296 3553 1343
rect 3562 1306 3565 1386
rect 3570 1313 3573 1326
rect 3650 1316 3653 1336
rect 3642 1313 3653 1316
rect 3562 1303 3573 1306
rect 3506 1253 3525 1256
rect 3546 1293 3553 1296
rect 3458 1203 3477 1206
rect 3506 1203 3509 1253
rect 3370 1163 3381 1166
rect 3370 1136 3373 1163
rect 3346 1043 3357 1046
rect 3362 1133 3373 1136
rect 3378 1133 3381 1146
rect 3386 1133 3389 1146
rect 3474 1143 3477 1203
rect 3346 1026 3349 1043
rect 3338 1023 3349 1026
rect 3322 963 3325 1006
rect 3338 996 3341 1023
rect 3346 1003 3349 1016
rect 3354 1013 3357 1036
rect 3362 996 3365 1133
rect 3370 1113 3373 1126
rect 3338 993 3349 996
rect 3322 883 3325 946
rect 3330 813 3333 926
rect 3338 923 3341 936
rect 3346 933 3349 993
rect 3358 993 3365 996
rect 3358 906 3361 993
rect 3370 933 3373 1016
rect 3474 1013 3477 1126
rect 3482 1113 3485 1126
rect 3490 1043 3493 1156
rect 3498 1133 3509 1136
rect 3482 1013 3485 1026
rect 3458 993 3461 1006
rect 3482 993 3485 1006
rect 3358 903 3365 906
rect 3362 883 3365 903
rect 3370 893 3373 926
rect 3386 923 3389 946
rect 3474 896 3477 926
rect 3466 893 3477 896
rect 3482 893 3485 926
rect 3354 813 3357 826
rect 3330 793 3333 806
rect 3354 766 3357 786
rect 3282 713 3285 726
rect 3306 723 3309 766
rect 3354 763 3361 766
rect 3378 763 3381 806
rect 3386 793 3389 806
rect 3322 686 3325 736
rect 3346 723 3349 746
rect 3358 696 3361 763
rect 3354 693 3361 696
rect 3322 683 3333 686
rect 3266 596 3269 676
rect 3274 613 3277 636
rect 3282 603 3285 626
rect 3298 613 3301 636
rect 3258 593 3277 596
rect 3250 573 3261 576
rect 3146 503 3153 506
rect 3138 413 3141 426
rect 3114 373 3117 406
rect 3050 323 3077 326
rect 3026 313 3045 316
rect 2866 113 2869 126
rect 2874 123 2885 126
rect 2898 123 2901 146
rect 2930 133 2933 216
rect 2938 183 2941 216
rect 2986 123 2989 136
rect 3034 123 3037 246
rect 3042 213 3045 306
rect 3082 243 3085 366
rect 3106 283 3109 336
rect 3114 323 3117 336
rect 3146 303 3149 503
rect 3178 456 3181 546
rect 3202 513 3205 526
rect 3258 486 3261 573
rect 3290 523 3293 536
rect 3306 533 3309 566
rect 3330 563 3333 683
rect 3354 673 3357 693
rect 3354 613 3357 646
rect 3394 633 3397 886
rect 3418 763 3421 846
rect 3466 836 3469 893
rect 3466 833 3477 836
rect 3474 813 3477 833
rect 3490 813 3493 936
rect 3498 913 3501 936
rect 3506 836 3509 1126
rect 3522 1026 3525 1186
rect 3546 1123 3549 1293
rect 3570 1256 3573 1303
rect 3570 1253 3581 1256
rect 3554 1213 3557 1226
rect 3578 1176 3581 1253
rect 3642 1246 3645 1313
rect 3642 1243 3653 1246
rect 3570 1173 3581 1176
rect 3562 1103 3565 1116
rect 3518 1023 3525 1026
rect 3518 926 3521 1023
rect 3530 933 3533 1016
rect 3518 923 3525 926
rect 3506 833 3517 836
rect 3498 796 3501 816
rect 3494 793 3501 796
rect 3410 713 3413 726
rect 3410 603 3413 616
rect 3426 563 3429 736
rect 3450 673 3453 726
rect 3494 716 3497 793
rect 3506 723 3509 806
rect 3514 793 3517 833
rect 3494 713 3501 716
rect 3514 713 3517 736
rect 3450 613 3453 636
rect 3498 613 3501 713
rect 3522 576 3525 923
rect 3538 906 3541 1026
rect 3546 1013 3565 1016
rect 3546 993 3549 1006
rect 3570 993 3573 1173
rect 3586 1106 3589 1136
rect 3594 1133 3597 1216
rect 3602 1183 3605 1206
rect 3602 1123 3605 1176
rect 3618 1106 3621 1216
rect 3626 1203 3629 1226
rect 3634 1203 3637 1216
rect 3650 1183 3653 1243
rect 3658 1166 3661 1396
rect 3666 1373 3669 1416
rect 3674 1366 3677 1526
rect 3690 1493 3693 1536
rect 3698 1533 3701 1606
rect 3714 1603 3717 1616
rect 3722 1593 3725 1716
rect 3730 1713 3741 1716
rect 3738 1636 3741 1713
rect 3762 1676 3765 1763
rect 3786 1756 3789 1806
rect 3826 1793 3829 1816
rect 3874 1803 3877 1816
rect 3890 1813 3893 1826
rect 3898 1803 3901 1883
rect 3930 1876 3933 1926
rect 3938 1906 3941 1926
rect 3938 1903 3949 1906
rect 3922 1873 3933 1876
rect 3778 1753 3789 1756
rect 3778 1723 3781 1753
rect 3786 1733 3789 1746
rect 3730 1633 3741 1636
rect 3754 1673 3765 1676
rect 3730 1613 3733 1633
rect 3754 1616 3757 1673
rect 3746 1613 3757 1616
rect 3746 1556 3749 1613
rect 3746 1553 3753 1556
rect 3682 1393 3685 1426
rect 3670 1363 3677 1366
rect 3690 1363 3693 1436
rect 3706 1423 3709 1536
rect 3714 1513 3717 1526
rect 3730 1523 3733 1536
rect 3670 1236 3673 1363
rect 3650 1163 3661 1166
rect 3666 1233 3673 1236
rect 3586 1103 3597 1106
rect 3578 933 3581 1016
rect 3594 1006 3597 1103
rect 3610 1103 3621 1106
rect 3610 1036 3613 1103
rect 3610 1033 3621 1036
rect 3618 1013 3621 1033
rect 3586 1003 3597 1006
rect 3538 903 3549 906
rect 3546 836 3549 903
rect 3538 833 3549 836
rect 3530 813 3533 826
rect 3538 813 3541 833
rect 3530 793 3533 806
rect 3330 523 3333 556
rect 3386 533 3397 536
rect 3426 523 3429 546
rect 3450 523 3453 536
rect 3250 483 3261 486
rect 3178 453 3189 456
rect 3186 396 3189 453
rect 3210 413 3213 426
rect 3178 393 3189 396
rect 3178 376 3181 393
rect 3170 373 3181 376
rect 3226 373 3229 406
rect 3154 293 3157 326
rect 3082 213 3085 236
rect 3146 213 3149 226
rect 3066 193 3069 206
rect 3170 193 3173 373
rect 3250 356 3253 483
rect 3258 413 3261 436
rect 3314 403 3317 426
rect 3330 386 3333 416
rect 3338 393 3341 416
rect 3362 413 3365 426
rect 3362 393 3365 406
rect 3378 403 3381 416
rect 3394 413 3397 446
rect 3402 406 3405 416
rect 3410 413 3413 426
rect 3450 413 3453 516
rect 3386 403 3405 406
rect 3242 353 3253 356
rect 3322 383 3333 386
rect 3194 303 3197 326
rect 3242 306 3245 353
rect 3258 343 3277 346
rect 3258 333 3261 343
rect 3258 313 3261 326
rect 3242 303 3261 306
rect 3274 303 3277 326
rect 3282 323 3285 336
rect 3322 326 3325 383
rect 3290 313 3293 326
rect 3322 323 3333 326
rect 3330 303 3333 323
rect 3258 213 3261 303
rect 3346 213 3349 356
rect 3354 323 3357 336
rect 3354 303 3357 316
rect 3050 123 3053 156
rect 3186 133 3189 196
rect 3234 133 3237 206
rect 3162 113 3165 126
rect 3258 113 3261 206
rect 3330 203 3349 206
rect 3330 133 3333 156
rect 3362 153 3365 336
rect 3370 306 3373 326
rect 3386 323 3389 403
rect 3394 316 3397 336
rect 3402 323 3405 346
rect 3386 313 3397 316
rect 3370 303 3377 306
rect 3374 236 3377 303
rect 3370 233 3377 236
rect 3370 133 3373 233
rect 3378 203 3381 216
rect 3386 213 3389 306
rect 3394 166 3397 216
rect 3402 206 3405 226
rect 3410 213 3413 336
rect 3402 203 3413 206
rect 3386 163 3397 166
rect 3362 103 3365 126
rect 3386 123 3389 163
rect 3394 133 3397 146
rect 3394 113 3405 116
rect 3410 103 3413 203
rect 3418 113 3421 406
rect 3426 313 3429 336
rect 3442 313 3445 406
rect 3458 336 3461 536
rect 3482 533 3485 576
rect 3514 573 3525 576
rect 3490 533 3493 546
rect 3466 353 3469 526
rect 3474 513 3485 516
rect 3474 423 3477 513
rect 3514 496 3517 573
rect 3546 566 3549 816
rect 3570 803 3573 926
rect 3586 853 3589 1003
rect 3594 923 3597 936
rect 3586 733 3589 816
rect 3602 736 3605 936
rect 3610 923 3613 986
rect 3626 873 3629 1106
rect 3650 1096 3653 1163
rect 3666 1103 3669 1233
rect 3674 1203 3677 1216
rect 3682 1133 3685 1326
rect 3690 1313 3693 1336
rect 3698 1286 3701 1326
rect 3694 1283 3701 1286
rect 3694 1166 3697 1283
rect 3706 1213 3709 1336
rect 3722 1226 3725 1416
rect 3722 1223 3729 1226
rect 3706 1173 3709 1206
rect 3694 1163 3701 1166
rect 3650 1093 3669 1096
rect 3634 816 3637 1086
rect 3642 1016 3645 1036
rect 3642 1013 3649 1016
rect 3658 1013 3661 1026
rect 3666 1013 3669 1093
rect 3646 946 3649 1013
rect 3674 983 3677 1006
rect 3642 943 3649 946
rect 3642 923 3645 943
rect 3658 913 3661 936
rect 3618 813 3637 816
rect 3602 733 3613 736
rect 3578 693 3581 726
rect 3538 563 3549 566
rect 3538 503 3541 563
rect 3562 533 3565 606
rect 3578 603 3581 616
rect 3594 613 3597 726
rect 3610 716 3613 733
rect 3606 713 3613 716
rect 3606 646 3609 713
rect 3602 643 3609 646
rect 3586 583 3589 606
rect 3602 603 3605 643
rect 3610 613 3613 626
rect 3602 566 3605 586
rect 3602 563 3609 566
rect 3514 493 3525 496
rect 3546 493 3549 526
rect 3482 413 3485 456
rect 3506 423 3509 436
rect 3482 393 3485 406
rect 3490 346 3493 416
rect 3522 413 3525 493
rect 3562 473 3565 526
rect 3578 456 3581 536
rect 3606 496 3609 563
rect 3618 516 3621 813
rect 3626 716 3629 806
rect 3642 733 3645 856
rect 3626 713 3637 716
rect 3634 626 3637 713
rect 3626 623 3637 626
rect 3650 623 3653 816
rect 3666 793 3669 936
rect 3682 933 3685 1056
rect 3698 956 3701 1163
rect 3714 1156 3717 1216
rect 3710 1153 3717 1156
rect 3710 1076 3713 1153
rect 3726 1146 3729 1223
rect 3722 1143 3729 1146
rect 3710 1073 3717 1076
rect 3714 1053 3717 1073
rect 3722 973 3725 1143
rect 3738 1126 3741 1536
rect 3750 1436 3753 1553
rect 3762 1446 3765 1666
rect 3794 1663 3797 1776
rect 3802 1676 3805 1726
rect 3818 1723 3821 1736
rect 3866 1723 3869 1736
rect 3802 1673 3821 1676
rect 3770 1613 3773 1646
rect 3786 1613 3789 1656
rect 3762 1443 3769 1446
rect 3750 1433 3757 1436
rect 3754 1413 3757 1433
rect 3746 1383 3749 1406
rect 3754 1366 3757 1406
rect 3750 1363 3757 1366
rect 3750 1186 3753 1363
rect 3766 1356 3769 1443
rect 3778 1413 3781 1606
rect 3794 1603 3797 1616
rect 3818 1556 3821 1673
rect 3906 1656 3909 1816
rect 3922 1803 3925 1873
rect 3946 1826 3949 1903
rect 3938 1823 3949 1826
rect 3906 1653 3917 1656
rect 3874 1613 3877 1636
rect 3866 1593 3869 1606
rect 3802 1553 3821 1556
rect 3794 1516 3797 1536
rect 3790 1513 3797 1516
rect 3790 1396 3793 1513
rect 3802 1406 3805 1553
rect 3810 1523 3813 1536
rect 3874 1533 3877 1566
rect 3882 1533 3885 1606
rect 3890 1603 3893 1616
rect 3898 1613 3901 1646
rect 3914 1606 3917 1653
rect 3906 1603 3917 1606
rect 3906 1533 3909 1603
rect 3930 1593 3933 1816
rect 3938 1803 3941 1823
rect 3946 1773 3949 1806
rect 3978 1803 3981 1926
rect 3986 1756 3989 1816
rect 4026 1813 4029 1946
rect 4074 1933 4077 1946
rect 4154 1933 4173 1936
rect 4202 1933 4205 1946
rect 4122 1913 4125 1926
rect 4154 1923 4157 1933
rect 4162 1906 4165 1926
rect 4154 1903 4165 1906
rect 4154 1836 4157 1903
rect 4154 1833 4165 1836
rect 3994 1783 3997 1806
rect 3954 1733 3957 1756
rect 3978 1753 3989 1756
rect 3962 1733 3973 1736
rect 3946 1626 3949 1726
rect 3978 1656 3981 1753
rect 3986 1733 3989 1746
rect 4010 1733 4013 1756
rect 4042 1733 4045 1806
rect 4066 1796 4069 1816
rect 4058 1793 4069 1796
rect 3994 1686 3997 1706
rect 3994 1683 4005 1686
rect 4050 1683 4053 1776
rect 4058 1733 4061 1793
rect 4074 1773 4077 1826
rect 4098 1756 4101 1776
rect 3938 1623 3949 1626
rect 3938 1603 3941 1623
rect 3962 1613 3965 1656
rect 3978 1653 3989 1656
rect 3978 1613 3981 1646
rect 3826 1513 3829 1526
rect 3842 1513 3845 1526
rect 3818 1413 3821 1426
rect 3802 1403 3821 1406
rect 3790 1393 3797 1396
rect 3762 1353 3769 1356
rect 3762 1196 3765 1353
rect 3794 1346 3797 1393
rect 3794 1343 3805 1346
rect 3778 1333 3789 1336
rect 3770 1306 3773 1326
rect 3770 1303 3777 1306
rect 3774 1236 3777 1303
rect 3786 1253 3789 1326
rect 3770 1233 3777 1236
rect 3770 1213 3773 1233
rect 3802 1226 3805 1343
rect 3818 1313 3821 1403
rect 3834 1353 3837 1416
rect 3842 1413 3845 1466
rect 3874 1463 3877 1526
rect 3906 1503 3909 1526
rect 3922 1406 3925 1536
rect 3930 1533 3933 1556
rect 3954 1516 3957 1606
rect 3970 1593 3973 1606
rect 3938 1513 3957 1516
rect 3938 1413 3941 1513
rect 3954 1413 3957 1426
rect 3866 1363 3869 1406
rect 3890 1346 3893 1406
rect 3826 1323 3845 1326
rect 3858 1323 3861 1336
rect 3842 1296 3845 1323
rect 3794 1223 3805 1226
rect 3834 1293 3845 1296
rect 3834 1226 3837 1293
rect 3834 1223 3845 1226
rect 3762 1193 3773 1196
rect 3750 1183 3757 1186
rect 3734 1123 3741 1126
rect 3734 1036 3737 1123
rect 3730 1033 3737 1036
rect 3730 1013 3733 1033
rect 3730 983 3733 1006
rect 3738 1003 3741 1026
rect 3746 1013 3749 1126
rect 3754 1013 3757 1183
rect 3770 1106 3773 1193
rect 3794 1156 3797 1223
rect 3794 1153 3805 1156
rect 3762 1103 3773 1106
rect 3762 1083 3765 1103
rect 3762 1013 3765 1026
rect 3690 953 3701 956
rect 3690 833 3693 953
rect 3698 923 3701 946
rect 3706 896 3709 966
rect 3714 913 3717 926
rect 3706 893 3717 896
rect 3626 566 3629 623
rect 3666 616 3669 736
rect 3674 703 3677 726
rect 3666 613 3673 616
rect 3682 613 3685 816
rect 3690 803 3693 826
rect 3634 593 3637 606
rect 3626 563 3645 566
rect 3626 523 3629 546
rect 3618 513 3629 516
rect 3562 453 3581 456
rect 3602 493 3609 496
rect 3546 416 3549 436
rect 3514 393 3517 406
rect 3482 343 3493 346
rect 3458 333 3469 336
rect 3434 223 3437 296
rect 3434 173 3437 206
rect 3442 193 3445 206
rect 3442 133 3445 186
rect 3450 113 3453 226
rect 3466 223 3469 316
rect 3482 303 3485 343
rect 3514 333 3517 376
rect 3522 333 3525 346
rect 3514 293 3517 316
rect 3474 213 3477 226
rect 3466 133 3469 146
rect 3490 113 3493 286
rect 3522 223 3525 326
rect 3530 323 3533 416
rect 3538 413 3549 416
rect 3538 293 3541 413
rect 3546 383 3549 406
rect 3562 363 3565 453
rect 3570 333 3573 346
rect 3554 293 3557 316
rect 3538 213 3541 226
rect 3578 213 3581 336
rect 3578 183 3581 206
rect 3514 123 3517 146
rect 3586 123 3589 216
rect 3602 213 3605 493
rect 3626 456 3629 513
rect 3626 453 3633 456
rect 3610 393 3613 416
rect 3630 406 3633 453
rect 3626 403 3633 406
rect 3626 383 3629 403
rect 3610 316 3613 336
rect 3642 323 3645 563
rect 3650 536 3653 606
rect 3658 583 3661 606
rect 3670 556 3673 613
rect 3690 603 3693 796
rect 3698 716 3701 816
rect 3714 813 3717 893
rect 3722 823 3725 936
rect 3730 823 3733 936
rect 3738 923 3741 996
rect 3746 906 3749 1006
rect 3754 943 3757 1006
rect 3770 983 3773 1006
rect 3754 913 3757 926
rect 3746 903 3757 906
rect 3706 733 3709 806
rect 3738 756 3741 836
rect 3754 826 3757 903
rect 3754 823 3761 826
rect 3722 753 3741 756
rect 3698 713 3709 716
rect 3706 636 3709 713
rect 3698 633 3709 636
rect 3698 613 3701 633
rect 3706 556 3709 606
rect 3666 553 3673 556
rect 3650 533 3661 536
rect 3658 416 3661 533
rect 3666 513 3669 553
rect 3658 413 3665 416
rect 3650 343 3653 406
rect 3662 356 3665 413
rect 3658 353 3665 356
rect 3610 313 3621 316
rect 3618 256 3621 313
rect 3610 253 3621 256
rect 3610 203 3613 253
rect 3634 213 3637 236
rect 3650 223 3653 336
rect 3658 333 3661 353
rect 3658 303 3661 326
rect 3626 143 3629 206
rect 3666 203 3669 336
rect 3674 233 3677 536
rect 3690 516 3693 556
rect 3698 553 3709 556
rect 3722 556 3725 753
rect 3738 566 3741 746
rect 3746 703 3749 816
rect 3758 756 3761 823
rect 3754 753 3761 756
rect 3754 733 3757 753
rect 3762 713 3765 726
rect 3770 706 3773 976
rect 3778 923 3781 1046
rect 3786 993 3789 1136
rect 3794 1023 3797 1126
rect 3802 1006 3805 1153
rect 3810 1133 3813 1216
rect 3842 1203 3845 1223
rect 3858 1216 3861 1316
rect 3858 1213 3865 1216
rect 3810 1013 3813 1126
rect 3794 936 3797 1006
rect 3802 1003 3813 1006
rect 3790 933 3797 936
rect 3778 803 3781 866
rect 3790 826 3793 933
rect 3802 903 3805 926
rect 3810 896 3813 1003
rect 3818 983 3821 1126
rect 3826 1083 3829 1136
rect 3802 893 3813 896
rect 3790 823 3797 826
rect 3786 793 3789 806
rect 3762 703 3773 706
rect 3738 563 3749 566
rect 3722 553 3733 556
rect 3698 523 3701 553
rect 3706 533 3709 546
rect 3714 523 3717 536
rect 3686 513 3693 516
rect 3686 436 3689 513
rect 3686 433 3693 436
rect 3682 193 3685 416
rect 3690 403 3693 433
rect 3690 306 3693 336
rect 3698 323 3701 516
rect 3706 393 3709 406
rect 3690 303 3697 306
rect 3714 303 3717 496
rect 3722 403 3725 536
rect 3730 493 3733 553
rect 3730 393 3733 476
rect 3746 456 3749 563
rect 3738 453 3749 456
rect 3722 333 3725 386
rect 3738 326 3741 453
rect 3762 436 3765 703
rect 3770 476 3773 536
rect 3778 523 3781 736
rect 3786 733 3789 746
rect 3786 683 3789 726
rect 3786 533 3789 556
rect 3794 533 3797 823
rect 3802 803 3805 893
rect 3802 696 3805 796
rect 3810 713 3813 816
rect 3818 723 3821 786
rect 3826 733 3829 1016
rect 3842 1013 3845 1136
rect 3850 1106 3853 1206
rect 3862 1166 3865 1213
rect 3858 1163 3865 1166
rect 3858 1133 3861 1163
rect 3866 1113 3869 1126
rect 3850 1103 3857 1106
rect 3854 1026 3857 1103
rect 3874 1046 3877 1346
rect 3882 1343 3893 1346
rect 3906 1343 3909 1406
rect 3922 1403 3933 1406
rect 3962 1403 3965 1516
rect 3970 1403 3973 1416
rect 3882 1323 3885 1343
rect 3906 1256 3909 1336
rect 3930 1333 3933 1403
rect 3986 1366 3989 1653
rect 4002 1626 4005 1683
rect 3994 1623 4005 1626
rect 3994 1576 3997 1623
rect 4034 1613 4037 1656
rect 4010 1593 4013 1606
rect 3994 1573 4005 1576
rect 4002 1466 4005 1573
rect 4026 1513 4029 1606
rect 4042 1603 4045 1616
rect 4050 1593 4053 1606
rect 4058 1603 4061 1616
rect 4066 1603 4069 1726
rect 4074 1716 4077 1756
rect 4094 1753 4101 1756
rect 4074 1713 4085 1716
rect 4082 1656 4085 1713
rect 4094 1706 4097 1753
rect 4106 1716 4109 1746
rect 4122 1733 4125 1816
rect 4130 1773 4133 1816
rect 4162 1813 4165 1833
rect 4138 1793 4141 1806
rect 4170 1803 4173 1916
rect 4178 1813 4181 1826
rect 4130 1733 4133 1756
rect 4146 1733 4157 1736
rect 4162 1733 4165 1746
rect 4106 1713 4117 1716
rect 4094 1703 4101 1706
rect 4074 1653 4085 1656
rect 4074 1593 4077 1653
rect 4090 1613 4093 1636
rect 3994 1463 4005 1466
rect 3994 1386 3997 1463
rect 4018 1413 4021 1446
rect 4002 1393 4005 1406
rect 3994 1383 4013 1386
rect 3986 1363 3997 1366
rect 3914 1286 3917 1306
rect 3914 1283 3925 1286
rect 3850 1023 3857 1026
rect 3866 1043 3877 1046
rect 3890 1253 3909 1256
rect 3850 1003 3853 1023
rect 3866 976 3869 1043
rect 3890 1003 3893 1253
rect 3922 1176 3925 1283
rect 3978 1276 3981 1326
rect 3994 1303 3997 1363
rect 3978 1273 3997 1276
rect 3914 1173 3925 1176
rect 3938 1176 3941 1216
rect 3938 1173 3957 1176
rect 3898 1123 3901 1136
rect 3906 1133 3909 1166
rect 3906 1013 3909 1036
rect 3850 933 3853 976
rect 3866 973 3885 976
rect 3858 933 3861 966
rect 3834 783 3837 816
rect 3874 813 3877 836
rect 3834 723 3837 736
rect 3842 723 3845 736
rect 3802 693 3813 696
rect 3810 526 3813 693
rect 3786 513 3789 526
rect 3802 523 3813 526
rect 3770 473 3789 476
rect 3746 433 3765 436
rect 3746 376 3749 433
rect 3786 413 3789 473
rect 3746 373 3753 376
rect 3722 323 3741 326
rect 3626 113 3629 136
rect 3674 123 3677 136
rect 3694 106 3697 303
rect 3706 213 3709 256
rect 3690 103 3697 106
rect 3690 86 3693 103
rect 2370 0 2389 3
rect 2530 83 2541 86
rect 3682 83 3693 86
rect 2530 0 2533 83
rect 2666 0 2669 16
rect 3682 0 3685 83
rect 3706 0 3709 196
rect 3714 133 3717 206
rect 3722 193 3725 323
rect 3750 316 3753 373
rect 3762 366 3765 406
rect 3762 363 3773 366
rect 3770 333 3773 363
rect 3746 313 3753 316
rect 3746 253 3749 313
rect 3730 213 3733 226
rect 3802 213 3805 523
rect 3826 466 3829 696
rect 3834 526 3837 606
rect 3834 523 3845 526
rect 3842 506 3845 523
rect 3842 503 3849 506
rect 3826 463 3833 466
rect 3830 376 3833 463
rect 3846 436 3849 503
rect 3842 433 3849 436
rect 3830 373 3837 376
rect 3818 323 3821 346
rect 3730 183 3733 206
rect 3762 203 3781 206
rect 3754 123 3757 196
rect 3810 183 3813 206
rect 3778 113 3781 146
rect 3818 113 3821 216
rect 3834 213 3837 373
rect 3826 123 3829 206
rect 3842 76 3845 433
rect 3850 116 3853 406
rect 3858 323 3861 806
rect 3866 793 3869 806
rect 3882 803 3885 973
rect 3898 873 3901 916
rect 3890 733 3893 826
rect 3906 813 3909 836
rect 3890 613 3893 716
rect 3882 593 3885 606
rect 3898 603 3901 796
rect 3906 783 3909 806
rect 3914 776 3917 1173
rect 3954 1133 3957 1173
rect 3970 1143 3973 1216
rect 3978 1203 3981 1216
rect 3946 1113 3949 1126
rect 3970 1083 3973 1136
rect 3954 1013 3957 1056
rect 3962 1006 3965 1026
rect 3930 993 3933 1006
rect 3922 916 3925 936
rect 3946 933 3949 1006
rect 3958 1003 3965 1006
rect 3958 926 3961 1003
rect 3954 923 3961 926
rect 3922 913 3933 916
rect 3930 826 3933 913
rect 3922 823 3933 826
rect 3922 793 3925 823
rect 3938 803 3949 806
rect 3954 803 3957 923
rect 3962 786 3965 826
rect 3970 816 3973 936
rect 3978 923 3981 946
rect 3970 813 3981 816
rect 3978 796 3981 813
rect 3946 783 3965 786
rect 3970 793 3981 796
rect 3914 773 3925 776
rect 3922 716 3925 773
rect 3914 713 3925 716
rect 3906 613 3909 706
rect 3914 693 3917 713
rect 3946 666 3949 783
rect 3970 736 3973 793
rect 3962 733 3973 736
rect 3986 736 3989 1236
rect 3994 1203 3997 1273
rect 4010 1226 4013 1383
rect 4002 1223 4013 1226
rect 4002 1136 4005 1223
rect 4010 1183 4013 1206
rect 3998 1133 4005 1136
rect 4018 1133 4021 1146
rect 3998 996 4001 1133
rect 4010 1003 4013 1126
rect 4018 1013 4021 1046
rect 4026 1023 4029 1336
rect 4034 1286 4037 1536
rect 4050 1523 4053 1536
rect 4050 1436 4053 1516
rect 4066 1513 4069 1526
rect 4046 1433 4053 1436
rect 4046 1346 4049 1433
rect 4046 1343 4053 1346
rect 4042 1303 4045 1326
rect 4050 1323 4053 1343
rect 4034 1283 4045 1286
rect 4042 1226 4045 1283
rect 4042 1223 4053 1226
rect 4034 1133 4037 1166
rect 4034 1013 4037 1066
rect 3998 993 4005 996
rect 3994 903 3997 926
rect 4002 836 4005 993
rect 4026 943 4029 1006
rect 4042 993 4045 1216
rect 4050 986 4053 1223
rect 4058 1003 4061 1426
rect 4066 1333 4069 1426
rect 4074 1423 4077 1536
rect 4082 1533 4085 1606
rect 4098 1603 4101 1703
rect 4114 1646 4117 1713
rect 4138 1696 4141 1726
rect 4106 1643 4117 1646
rect 4130 1693 4141 1696
rect 4130 1646 4133 1693
rect 4130 1643 4141 1646
rect 4074 1313 4077 1416
rect 4082 1316 4085 1336
rect 4090 1333 4093 1596
rect 4098 1523 4101 1536
rect 4106 1373 4109 1643
rect 4114 1603 4117 1616
rect 4114 1523 4117 1536
rect 4122 1423 4125 1536
rect 4130 1533 4133 1626
rect 4138 1603 4141 1643
rect 4146 1556 4149 1726
rect 4154 1703 4157 1726
rect 4178 1723 4181 1806
rect 4186 1783 4189 1806
rect 4194 1793 4197 1806
rect 4202 1723 4205 1736
rect 4210 1703 4213 1836
rect 4226 1813 4229 1826
rect 4234 1803 4237 1926
rect 4242 1813 4245 1836
rect 4258 1796 4261 1826
rect 4242 1793 4261 1796
rect 4242 1706 4245 1793
rect 4266 1783 4269 1806
rect 4282 1803 4285 1926
rect 4294 1786 4297 1953
rect 4322 1926 4325 1946
rect 4338 1943 4341 2016
rect 4354 2013 4373 2016
rect 4362 1993 4365 2006
rect 4370 2003 4373 2013
rect 4394 1993 4397 2196
rect 4418 2193 4421 2206
rect 4290 1783 4297 1786
rect 4258 1733 4277 1736
rect 4258 1723 4261 1733
rect 4266 1713 4269 1726
rect 4242 1703 4253 1706
rect 4162 1613 4165 1636
rect 4138 1553 4149 1556
rect 4130 1513 4133 1526
rect 4114 1403 4117 1416
rect 4122 1333 4125 1406
rect 4138 1403 4141 1553
rect 4146 1523 4149 1546
rect 4154 1533 4157 1606
rect 4170 1593 4173 1606
rect 4178 1603 4181 1616
rect 4186 1613 4189 1646
rect 4194 1533 4197 1546
rect 4202 1456 4205 1686
rect 4234 1613 4237 1656
rect 4250 1636 4253 1703
rect 4242 1633 4253 1636
rect 4226 1546 4229 1606
rect 4242 1593 4245 1633
rect 4290 1626 4293 1783
rect 4306 1643 4309 1926
rect 4322 1923 4333 1926
rect 4330 1866 4333 1923
rect 4322 1863 4333 1866
rect 4322 1803 4325 1863
rect 4386 1856 4389 1946
rect 4386 1853 4397 1856
rect 4330 1733 4333 1756
rect 4346 1733 4349 1816
rect 4394 1776 4397 1853
rect 4386 1773 4397 1776
rect 4290 1623 4301 1626
rect 4250 1603 4253 1616
rect 4290 1593 4293 1606
rect 4218 1543 4229 1546
rect 4218 1526 4221 1543
rect 4226 1533 4237 1536
rect 4242 1533 4245 1566
rect 4218 1523 4229 1526
rect 4202 1453 4209 1456
rect 4162 1403 4165 1416
rect 4082 1313 4093 1316
rect 4066 1286 4069 1306
rect 4066 1283 4077 1286
rect 4074 1226 4077 1283
rect 4066 1223 4077 1226
rect 4066 1203 4069 1223
rect 4090 1206 4093 1313
rect 4114 1296 4117 1326
rect 4082 1203 4093 1206
rect 4106 1293 4117 1296
rect 4082 1183 4085 1203
rect 4066 1086 4069 1176
rect 4082 1133 4085 1166
rect 4106 1156 4109 1293
rect 4122 1236 4125 1326
rect 4130 1303 4133 1326
rect 4118 1233 4125 1236
rect 4118 1186 4121 1233
rect 4138 1213 4141 1376
rect 4206 1366 4209 1453
rect 4202 1363 4209 1366
rect 4202 1346 4205 1363
rect 4194 1343 4205 1346
rect 4218 1343 4221 1416
rect 4226 1413 4229 1523
rect 4234 1406 4237 1426
rect 4146 1313 4149 1326
rect 4170 1323 4181 1326
rect 4194 1266 4197 1343
rect 4226 1336 4229 1406
rect 4234 1403 4241 1406
rect 4210 1333 4229 1336
rect 4194 1263 4205 1266
rect 4118 1183 4125 1186
rect 4106 1153 4113 1156
rect 4074 1103 4077 1126
rect 4066 1083 4073 1086
rect 4070 996 4073 1083
rect 4090 1066 4093 1126
rect 4098 1123 4101 1136
rect 4082 1063 4093 1066
rect 4082 1003 4085 1063
rect 4110 1056 4113 1153
rect 4122 1066 4125 1183
rect 4122 1063 4129 1066
rect 4090 1013 4093 1056
rect 4110 1053 4117 1056
rect 4106 1013 4109 1036
rect 4114 1013 4117 1053
rect 4126 1006 4129 1063
rect 4034 983 4053 986
rect 4066 993 4073 996
rect 4010 843 4013 926
rect 4002 833 4013 836
rect 4010 816 4013 833
rect 4010 813 4017 816
rect 3986 733 3993 736
rect 3962 686 3965 733
rect 3962 683 3973 686
rect 3946 663 3965 666
rect 3962 613 3965 663
rect 3914 583 3917 606
rect 3882 533 3885 546
rect 3890 443 3893 526
rect 3898 413 3901 536
rect 3914 456 3917 556
rect 3922 523 3925 606
rect 3970 603 3973 683
rect 3978 613 3981 726
rect 3990 616 3993 733
rect 3990 613 3997 616
rect 3938 566 3941 586
rect 3986 583 3989 606
rect 3934 563 3941 566
rect 3934 506 3937 563
rect 3946 516 3949 536
rect 3962 516 3965 546
rect 3970 533 3973 556
rect 3946 513 3957 516
rect 3962 513 3973 516
rect 3934 503 3941 506
rect 3938 456 3941 503
rect 3914 453 3921 456
rect 3938 453 3945 456
rect 3906 406 3909 446
rect 3858 203 3861 226
rect 3874 153 3877 406
rect 3898 403 3909 406
rect 3890 333 3893 356
rect 3898 213 3901 403
rect 3918 396 3921 453
rect 3914 393 3921 396
rect 3914 353 3917 393
rect 3942 376 3945 453
rect 3922 346 3925 376
rect 3906 333 3909 346
rect 3914 343 3925 346
rect 3938 373 3945 376
rect 3914 323 3917 343
rect 3930 306 3933 336
rect 3922 303 3933 306
rect 3922 226 3925 303
rect 3922 223 3933 226
rect 3906 193 3909 206
rect 3922 183 3925 206
rect 3930 166 3933 223
rect 3938 213 3941 373
rect 3946 333 3949 346
rect 3954 333 3957 513
rect 3970 446 3973 513
rect 3994 503 3997 613
rect 4002 506 4005 806
rect 4014 636 4017 813
rect 4010 633 4017 636
rect 4010 613 4013 633
rect 4026 623 4029 826
rect 4034 803 4037 983
rect 4042 933 4045 956
rect 4050 816 4053 936
rect 4058 923 4061 946
rect 4050 813 4061 816
rect 4042 803 4053 806
rect 4058 796 4061 813
rect 4050 793 4061 796
rect 4010 513 4013 526
rect 4002 503 4009 506
rect 3962 443 3973 446
rect 3962 343 3965 443
rect 4006 406 4009 503
rect 4018 413 4021 536
rect 3978 363 3981 406
rect 4006 403 4013 406
rect 4026 403 4029 616
rect 4042 613 4045 626
rect 4034 556 4037 606
rect 4050 603 4053 793
rect 4066 776 4069 993
rect 4098 943 4101 1006
rect 4106 986 4109 1006
rect 4122 1003 4129 1006
rect 4106 983 4113 986
rect 4110 936 4113 983
rect 4106 933 4113 936
rect 4074 873 4077 916
rect 4090 893 4093 926
rect 4082 813 4085 836
rect 4098 813 4101 826
rect 4062 773 4069 776
rect 4062 656 4065 773
rect 4062 653 4069 656
rect 4058 613 4061 636
rect 4034 553 4045 556
rect 4034 533 4037 546
rect 4042 456 4045 553
rect 4050 513 4053 526
rect 4042 453 4049 456
rect 3954 313 3957 326
rect 3962 236 3965 336
rect 3978 333 3981 356
rect 4002 313 4005 326
rect 4010 296 4013 403
rect 3954 233 3965 236
rect 4006 293 4013 296
rect 3954 186 3957 233
rect 4006 216 4009 293
rect 3954 183 3965 186
rect 3922 163 3933 166
rect 3858 133 3877 136
rect 3858 123 3861 133
rect 3850 113 3861 116
rect 3866 113 3869 126
rect 3834 73 3845 76
rect 3834 16 3837 73
rect 3834 13 3845 16
rect 3842 0 3845 13
rect 3858 0 3861 113
rect 3922 106 3925 163
rect 3938 133 3941 156
rect 3962 123 3965 183
rect 3970 143 3973 206
rect 3994 193 3997 216
rect 4006 213 4013 216
rect 4010 193 4013 213
rect 4018 133 4021 336
rect 4026 323 4029 396
rect 4046 346 4049 453
rect 4034 333 4037 346
rect 4042 343 4049 346
rect 4042 326 4045 343
rect 4034 323 4045 326
rect 4018 113 4021 126
rect 4034 123 4037 323
rect 4058 236 4061 536
rect 4066 383 4069 653
rect 4074 493 4077 806
rect 4082 716 4085 806
rect 4106 803 4109 933
rect 4122 903 4125 1003
rect 4114 786 4117 836
rect 4122 813 4125 886
rect 4110 783 4117 786
rect 4082 713 4089 716
rect 4086 556 4089 713
rect 4082 553 4089 556
rect 4082 523 4085 553
rect 4090 506 4093 536
rect 4086 503 4093 506
rect 4086 436 4089 503
rect 4098 456 4101 736
rect 4110 726 4113 783
rect 4122 733 4125 806
rect 4110 723 4117 726
rect 4114 633 4117 723
rect 4122 613 4125 646
rect 4106 593 4109 606
rect 4114 583 4117 606
rect 4130 603 4133 926
rect 4138 916 4141 1206
rect 4162 1163 4165 1216
rect 4202 1166 4205 1263
rect 4194 1163 4205 1166
rect 4146 993 4149 1006
rect 4162 1003 4165 1126
rect 4194 1086 4197 1163
rect 4194 1083 4205 1086
rect 4170 1013 4173 1046
rect 4186 1013 4189 1066
rect 4194 1013 4197 1036
rect 4178 946 4181 1006
rect 4194 993 4197 1006
rect 4146 933 4149 946
rect 4162 943 4181 946
rect 4138 913 4145 916
rect 4142 796 4145 913
rect 4154 803 4157 926
rect 4162 923 4165 943
rect 4162 913 4181 916
rect 4162 903 4165 913
rect 4142 793 4157 796
rect 4138 613 4141 726
rect 4154 686 4157 793
rect 4170 703 4173 816
rect 4178 733 4181 906
rect 4186 823 4189 936
rect 4194 933 4197 946
rect 4194 813 4197 916
rect 4202 836 4205 1083
rect 4210 903 4213 1333
rect 4238 1326 4241 1403
rect 4234 1323 4241 1326
rect 4250 1323 4253 1426
rect 4258 1403 4261 1516
rect 4266 1493 4269 1516
rect 4298 1513 4301 1623
rect 4314 1613 4317 1636
rect 4306 1536 4309 1606
rect 4330 1603 4333 1726
rect 4354 1693 4357 1726
rect 4370 1713 4373 1726
rect 4386 1666 4389 1773
rect 4394 1733 4397 1746
rect 4410 1733 4413 1816
rect 4382 1663 4389 1666
rect 4338 1613 4341 1646
rect 4338 1593 4341 1606
rect 4370 1603 4373 1626
rect 4382 1616 4385 1663
rect 4378 1613 4385 1616
rect 4394 1613 4397 1656
rect 4306 1533 4317 1536
rect 4314 1523 4317 1533
rect 4258 1323 4261 1336
rect 4218 1143 4221 1216
rect 4234 1193 4237 1323
rect 4266 1313 4269 1336
rect 4218 1133 4229 1136
rect 4258 1133 4261 1216
rect 4218 986 4221 1133
rect 4226 1096 4229 1126
rect 4266 1103 4269 1306
rect 4274 1146 4277 1416
rect 4282 1333 4285 1406
rect 4322 1356 4325 1536
rect 4330 1533 4333 1556
rect 4370 1503 4373 1516
rect 4378 1473 4381 1613
rect 4386 1523 4389 1606
rect 4402 1603 4405 1726
rect 4394 1456 4397 1536
rect 4402 1503 4405 1516
rect 4418 1513 4421 2186
rect 4434 2173 4437 2206
rect 4450 2203 4453 2223
rect 4442 2133 4445 2146
rect 4458 2136 4461 2296
rect 4466 2286 4469 2386
rect 4490 2323 4493 2346
rect 4466 2283 4477 2286
rect 4474 2203 4477 2283
rect 4506 2253 4509 2463
rect 4522 2443 4525 2713
rect 4546 2646 4549 2786
rect 4554 2743 4557 2806
rect 4562 2766 4565 2806
rect 4562 2763 4581 2766
rect 4554 2703 4557 2736
rect 4546 2643 4553 2646
rect 4550 2596 4553 2643
rect 4562 2613 4565 2756
rect 4570 2613 4573 2736
rect 4578 2726 4581 2763
rect 4586 2736 4589 2796
rect 4594 2753 4597 2833
rect 4606 2806 4609 2853
rect 4618 2813 4621 3056
rect 4626 3013 4629 3026
rect 4626 2923 4629 2996
rect 4634 2906 4637 3223
rect 4642 3186 4645 3206
rect 4674 3196 4677 3386
rect 4706 3333 4709 3386
rect 4730 3276 4733 3393
rect 4762 3366 4765 3483
rect 4778 3403 4781 3526
rect 4762 3363 4773 3366
rect 4770 3346 4773 3363
rect 4770 3343 4777 3346
rect 4722 3273 4733 3276
rect 4682 3203 4685 3226
rect 4722 3216 4725 3273
rect 4738 3223 4741 3326
rect 4690 3213 4709 3216
rect 4722 3213 4733 3216
rect 4674 3193 4685 3196
rect 4642 3183 4653 3186
rect 4650 3036 4653 3183
rect 4682 3133 4685 3193
rect 4690 3173 4693 3213
rect 4698 3193 4701 3206
rect 4730 3166 4733 3213
rect 4746 3203 4749 3316
rect 4774 3286 4777 3343
rect 4786 3313 4789 3326
rect 4770 3283 4777 3286
rect 4770 3216 4773 3283
rect 4722 3163 4733 3166
rect 4706 3123 4709 3146
rect 4630 2903 4637 2906
rect 4642 3033 4653 3036
rect 4630 2826 4633 2903
rect 4626 2823 4633 2826
rect 4606 2803 4613 2806
rect 4610 2743 4613 2803
rect 4626 2763 4629 2823
rect 4642 2773 4645 3033
rect 4586 2733 4605 2736
rect 4578 2723 4597 2726
rect 4602 2706 4605 2733
rect 4594 2703 4605 2706
rect 4610 2733 4629 2736
rect 4594 2636 4597 2703
rect 4594 2633 4605 2636
rect 4594 2596 4597 2616
rect 4546 2593 4553 2596
rect 4590 2593 4597 2596
rect 4546 2523 4549 2593
rect 4554 2533 4557 2546
rect 4562 2506 4565 2526
rect 4554 2503 4565 2506
rect 4522 2413 4525 2426
rect 4554 2416 4557 2503
rect 4570 2423 4573 2536
rect 4554 2413 4573 2416
rect 4578 2413 4581 2576
rect 4590 2506 4593 2593
rect 4602 2513 4605 2633
rect 4610 2613 4613 2733
rect 4618 2706 4621 2726
rect 4618 2703 4629 2706
rect 4642 2703 4645 2736
rect 4626 2646 4629 2703
rect 4650 2696 4653 3016
rect 4658 2993 4661 3006
rect 4666 3003 4669 3116
rect 4690 3013 4709 3016
rect 4658 2823 4661 2936
rect 4666 2913 4669 2926
rect 4658 2733 4661 2746
rect 4666 2723 4669 2806
rect 4650 2693 4661 2696
rect 4618 2643 4629 2646
rect 4590 2503 4597 2506
rect 4586 2413 4589 2426
rect 4562 2313 4565 2326
rect 4570 2323 4573 2413
rect 4498 2193 4501 2216
rect 4570 2213 4573 2226
rect 4578 2213 4581 2396
rect 4594 2393 4597 2503
rect 4618 2456 4621 2643
rect 4634 2613 4637 2626
rect 4642 2613 4653 2616
rect 4626 2593 4629 2606
rect 4642 2573 4645 2606
rect 4626 2533 4637 2536
rect 4602 2386 4605 2456
rect 4618 2453 4629 2456
rect 4610 2413 4613 2436
rect 4586 2233 4589 2386
rect 4594 2383 4605 2386
rect 4594 2333 4597 2383
rect 4610 2333 4613 2346
rect 4602 2313 4605 2326
rect 4618 2323 4621 2426
rect 4626 2383 4629 2453
rect 4626 2306 4629 2336
rect 4634 2333 4637 2516
rect 4642 2453 4645 2566
rect 4650 2543 4653 2606
rect 4622 2303 4629 2306
rect 4586 2156 4589 2206
rect 4594 2203 4597 2216
rect 4602 2203 4605 2226
rect 4610 2213 4613 2236
rect 4622 2226 4625 2303
rect 4622 2223 4629 2226
rect 4586 2153 4597 2156
rect 4450 2133 4461 2136
rect 4474 2133 4477 2146
rect 4498 2133 4525 2136
rect 4586 2133 4589 2146
rect 4450 2116 4453 2133
rect 4498 2126 4501 2133
rect 4442 2113 4453 2116
rect 4442 2026 4445 2113
rect 4458 2096 4461 2126
rect 4482 2123 4501 2126
rect 4458 2093 4469 2096
rect 4466 2036 4469 2093
rect 4458 2033 4469 2036
rect 4442 2023 4453 2026
rect 4450 2003 4453 2023
rect 4458 2013 4461 2033
rect 4466 1933 4485 1936
rect 4434 1886 4437 1926
rect 4466 1923 4469 1933
rect 4434 1883 4445 1886
rect 4426 1783 4429 1806
rect 4426 1733 4429 1756
rect 4434 1693 4437 1816
rect 4442 1803 4445 1883
rect 4442 1676 4445 1726
rect 4434 1673 4445 1676
rect 4434 1626 4437 1673
rect 4434 1623 4445 1626
rect 4450 1623 4453 1816
rect 4458 1803 4461 1826
rect 4474 1813 4477 1926
rect 4490 1816 4493 2016
rect 4522 2003 4525 2126
rect 4538 2113 4541 2126
rect 4554 2016 4557 2126
rect 4594 2106 4597 2153
rect 4602 2116 4605 2136
rect 4618 2133 4621 2156
rect 4626 2143 4629 2223
rect 4634 2123 4637 2316
rect 4642 2203 4645 2446
rect 4650 2296 4653 2516
rect 4658 2503 4661 2693
rect 4666 2603 4669 2716
rect 4674 2696 4677 2986
rect 4682 2953 4685 3006
rect 4690 2993 4693 3013
rect 4698 2983 4701 3006
rect 4722 2976 4725 3163
rect 4754 3153 4757 3216
rect 4770 3213 4781 3216
rect 4762 3123 4765 3206
rect 4778 3106 4781 3213
rect 4770 3103 4781 3106
rect 4722 2973 4729 2976
rect 4690 2886 4693 2946
rect 4714 2923 4717 2956
rect 4690 2883 4701 2886
rect 4698 2766 4701 2883
rect 4726 2846 4729 2973
rect 4738 2856 4741 3086
rect 4762 3006 4765 3096
rect 4770 3083 4773 3103
rect 4758 3003 4765 3006
rect 4758 2946 4761 3003
rect 4758 2943 4765 2946
rect 4762 2923 4765 2943
rect 4770 2923 4773 2996
rect 4778 2933 4789 2936
rect 4738 2853 4745 2856
rect 4726 2843 4733 2846
rect 4722 2813 4725 2826
rect 4690 2763 4701 2766
rect 4674 2693 4681 2696
rect 4678 2626 4681 2693
rect 4674 2623 4681 2626
rect 4690 2623 4693 2763
rect 4714 2723 4717 2746
rect 4730 2713 4733 2843
rect 4742 2776 4745 2853
rect 4738 2773 4745 2776
rect 4674 2536 4677 2623
rect 4690 2613 4709 2616
rect 4682 2543 4685 2606
rect 4690 2593 4693 2613
rect 4698 2556 4701 2606
rect 4690 2553 4701 2556
rect 4690 2536 4693 2553
rect 4658 2413 4661 2446
rect 4666 2433 4669 2536
rect 4674 2533 4693 2536
rect 4674 2443 4677 2526
rect 4690 2483 4693 2533
rect 4706 2456 4709 2606
rect 4738 2563 4741 2773
rect 4778 2766 4781 2926
rect 4786 2913 4789 2926
rect 4794 2896 4797 3713
rect 4790 2893 4797 2896
rect 4790 2806 4793 2893
rect 4802 2813 4805 2936
rect 4790 2803 4797 2806
rect 4770 2763 4781 2766
rect 4770 2576 4773 2763
rect 4786 2723 4789 2736
rect 4794 2616 4797 2803
rect 4794 2613 4801 2616
rect 4770 2573 4777 2576
rect 4730 2523 4733 2546
rect 4774 2516 4777 2573
rect 4786 2523 4789 2606
rect 4798 2536 4801 2613
rect 4794 2533 4801 2536
rect 4774 2513 4781 2516
rect 4794 2513 4797 2533
rect 4730 2486 4733 2506
rect 4690 2453 4709 2456
rect 4674 2403 4677 2426
rect 4690 2383 4693 2453
rect 4714 2413 4717 2436
rect 4706 2366 4709 2396
rect 4702 2363 4709 2366
rect 4666 2323 4669 2336
rect 4690 2323 4693 2346
rect 4650 2293 4657 2296
rect 4654 2226 4657 2293
rect 4702 2246 4705 2363
rect 4714 2256 4717 2406
rect 4722 2393 4725 2486
rect 4730 2483 4737 2486
rect 4734 2366 4737 2483
rect 4770 2413 4773 2426
rect 4754 2366 4757 2386
rect 4734 2363 4741 2366
rect 4738 2286 4741 2363
rect 4750 2363 4757 2366
rect 4750 2316 4753 2363
rect 4762 2323 4765 2336
rect 4750 2313 4757 2316
rect 4730 2283 4741 2286
rect 4714 2253 4721 2256
rect 4702 2243 4709 2246
rect 4650 2223 4657 2226
rect 4650 2153 4653 2223
rect 4666 2213 4669 2236
rect 4682 2213 4685 2226
rect 4698 2213 4701 2226
rect 4666 2186 4669 2206
rect 4662 2183 4669 2186
rect 4662 2126 4665 2183
rect 4674 2133 4677 2206
rect 4706 2203 4709 2243
rect 4718 2206 4721 2253
rect 4730 2233 4733 2283
rect 4714 2203 4721 2206
rect 4714 2183 4717 2203
rect 4698 2133 4701 2166
rect 4662 2123 4669 2126
rect 4722 2123 4725 2136
rect 4602 2113 4613 2116
rect 4586 2103 4597 2106
rect 4586 2036 4589 2103
rect 4610 2056 4613 2113
rect 4602 2053 4613 2056
rect 4586 2033 4597 2036
rect 4602 2033 4605 2053
rect 4546 2013 4557 2016
rect 4594 2013 4597 2033
rect 4546 1946 4549 2013
rect 4570 1966 4573 2006
rect 4570 1963 4577 1966
rect 4506 1933 4509 1946
rect 4546 1943 4557 1946
rect 4482 1813 4493 1816
rect 4458 1733 4461 1796
rect 4466 1783 4469 1806
rect 4474 1733 4477 1746
rect 4482 1736 4485 1813
rect 4498 1786 4501 1816
rect 4506 1803 4509 1916
rect 4530 1913 4533 1926
rect 4554 1856 4557 1943
rect 4574 1886 4577 1963
rect 4586 1933 4605 1936
rect 4586 1923 4589 1933
rect 4546 1853 4557 1856
rect 4570 1883 4577 1886
rect 4514 1806 4517 1826
rect 4522 1813 4525 1846
rect 4514 1803 4525 1806
rect 4498 1783 4509 1786
rect 4482 1733 4493 1736
rect 4466 1703 4469 1726
rect 4442 1603 4445 1623
rect 4458 1616 4461 1656
rect 4450 1613 4461 1616
rect 4466 1613 4469 1646
rect 4442 1533 4453 1536
rect 4458 1523 4461 1606
rect 4474 1593 4477 1606
rect 4482 1603 4485 1726
rect 4490 1686 4493 1733
rect 4506 1726 4509 1783
rect 4530 1733 4533 1816
rect 4498 1723 4509 1726
rect 4498 1703 4501 1723
rect 4538 1716 4541 1846
rect 4530 1713 4541 1716
rect 4490 1683 4501 1686
rect 4498 1596 4501 1683
rect 4530 1636 4533 1713
rect 4514 1613 4517 1636
rect 4530 1633 4541 1636
rect 4490 1593 4501 1596
rect 4474 1533 4477 1546
rect 4490 1526 4493 1593
rect 4370 1453 4397 1456
rect 4354 1403 4357 1416
rect 4370 1396 4373 1453
rect 4370 1393 4381 1396
rect 4314 1353 4325 1356
rect 4282 1173 4285 1316
rect 4290 1303 4293 1326
rect 4314 1236 4317 1353
rect 4314 1233 4325 1236
rect 4274 1143 4293 1146
rect 4282 1113 4285 1126
rect 4226 1093 4237 1096
rect 4234 1026 4237 1093
rect 4290 1086 4293 1143
rect 4298 1133 4301 1156
rect 4314 1133 4317 1216
rect 4322 1123 4325 1233
rect 4330 1203 4333 1336
rect 4346 1333 4349 1376
rect 4378 1336 4381 1393
rect 4402 1373 4405 1406
rect 4418 1393 4421 1406
rect 4378 1333 4385 1336
rect 4370 1276 4373 1326
rect 4362 1273 4373 1276
rect 4330 1133 4333 1156
rect 4282 1083 4293 1086
rect 4226 1023 4237 1026
rect 4226 1003 4229 1023
rect 4218 983 4229 986
rect 4202 833 4213 836
rect 4186 733 4197 736
rect 4154 683 4165 686
rect 4146 613 4149 636
rect 4146 576 4149 606
rect 4162 576 4165 683
rect 4186 643 4189 726
rect 4186 593 4189 606
rect 4142 573 4149 576
rect 4154 573 4165 576
rect 4114 523 4117 536
rect 4142 506 4145 573
rect 4154 506 4157 573
rect 4162 523 4165 546
rect 4142 503 4149 506
rect 4154 503 4161 506
rect 4098 453 4109 456
rect 4086 433 4093 436
rect 4090 416 4093 433
rect 4106 426 4109 453
rect 4106 423 4117 426
rect 4074 413 4093 416
rect 4074 306 4077 336
rect 4082 323 4085 406
rect 4106 376 4109 416
rect 4090 373 4109 376
rect 4090 333 4093 373
rect 4050 233 4061 236
rect 4070 303 4077 306
rect 4070 236 4073 303
rect 4070 233 4077 236
rect 4050 226 4053 233
rect 4042 223 4053 226
rect 4042 106 4045 223
rect 4050 206 4053 216
rect 4058 213 4061 226
rect 4050 203 4069 206
rect 4074 203 4077 233
rect 4082 213 4085 306
rect 4050 123 4053 196
rect 4090 193 4093 206
rect 4106 183 4109 336
rect 4114 323 4117 423
rect 4122 213 4125 486
rect 4130 323 4133 496
rect 4146 483 4149 503
rect 4158 446 4161 503
rect 4154 443 4161 446
rect 4154 393 4157 443
rect 4162 333 4165 346
rect 4154 313 4157 326
rect 4170 323 4173 426
rect 4194 423 4197 726
rect 4202 603 4205 826
rect 4210 733 4213 833
rect 4226 826 4229 983
rect 4242 923 4245 1006
rect 4250 993 4253 1056
rect 4282 1026 4285 1083
rect 4282 1023 4293 1026
rect 4290 1003 4293 1023
rect 4298 986 4301 1106
rect 4294 983 4301 986
rect 4306 983 4309 1046
rect 4222 823 4229 826
rect 4250 823 4253 936
rect 4258 923 4261 936
rect 4222 756 4225 823
rect 4218 753 4225 756
rect 4210 633 4213 726
rect 4210 613 4213 626
rect 4218 573 4221 753
rect 4234 746 4237 806
rect 4250 803 4253 816
rect 4258 776 4261 816
rect 4250 773 4261 776
rect 4234 743 4241 746
rect 4226 546 4229 736
rect 4238 696 4241 743
rect 4250 713 4253 773
rect 4238 693 4245 696
rect 4242 636 4245 693
rect 4234 633 4245 636
rect 4234 593 4237 633
rect 4258 616 4261 746
rect 4266 733 4269 806
rect 4274 733 4277 926
rect 4282 903 4285 916
rect 4282 813 4285 836
rect 4294 806 4297 983
rect 4306 813 4309 936
rect 4314 933 4317 1006
rect 4322 986 4325 1026
rect 4330 1003 4333 1126
rect 4338 996 4341 1126
rect 4346 1103 4349 1136
rect 4354 1123 4357 1236
rect 4362 1203 4365 1273
rect 4382 1266 4385 1333
rect 4378 1263 4385 1266
rect 4378 1216 4381 1263
rect 4378 1213 4389 1216
rect 4378 1173 4381 1206
rect 4362 1113 4365 1136
rect 4370 1133 4381 1136
rect 4346 1013 4349 1036
rect 4370 1003 4373 1126
rect 4386 1116 4389 1213
rect 4382 1113 4389 1116
rect 4382 1036 4385 1113
rect 4382 1033 4389 1036
rect 4394 1033 4397 1346
rect 4434 1333 4437 1366
rect 4442 1326 4445 1516
rect 4474 1506 4477 1526
rect 4490 1523 4497 1526
rect 4466 1503 4477 1506
rect 4466 1426 4469 1503
rect 4466 1423 4477 1426
rect 4482 1423 4485 1516
rect 4494 1446 4497 1523
rect 4490 1443 4497 1446
rect 4458 1346 4461 1366
rect 4386 1013 4389 1033
rect 4338 993 4349 996
rect 4322 983 4333 986
rect 4322 933 4325 966
rect 4330 943 4333 983
rect 4346 926 4349 993
rect 4330 923 4349 926
rect 4362 923 4365 936
rect 4378 926 4381 1006
rect 4386 933 4389 1006
rect 4394 963 4397 1016
rect 4402 1003 4405 1216
rect 4426 1203 4429 1326
rect 4434 1323 4445 1326
rect 4434 1313 4437 1323
rect 4418 1133 4421 1196
rect 4442 1193 4445 1323
rect 4454 1343 4461 1346
rect 4454 1226 4457 1343
rect 4450 1223 4457 1226
rect 4442 1113 4445 1126
rect 4410 1013 4413 1026
rect 4418 1006 4421 1036
rect 4410 1003 4421 1006
rect 4394 933 4397 956
rect 4378 923 4389 926
rect 4410 923 4413 1003
rect 4418 933 4429 936
rect 4434 933 4437 1006
rect 4314 893 4317 916
rect 4330 856 4333 923
rect 4370 903 4373 916
rect 4322 853 4333 856
rect 4294 803 4301 806
rect 4298 783 4301 803
rect 4306 776 4309 806
rect 4322 803 4325 853
rect 4306 773 4313 776
rect 4282 623 4285 766
rect 4290 723 4293 736
rect 4298 733 4301 746
rect 4298 703 4301 726
rect 4310 696 4313 773
rect 4322 716 4325 786
rect 4330 763 4333 836
rect 4338 783 4341 806
rect 4346 733 4349 826
rect 4354 793 4357 806
rect 4322 713 4333 716
rect 4354 713 4357 726
rect 4306 693 4313 696
rect 4250 613 4261 616
rect 4218 543 4229 546
rect 4218 446 4221 543
rect 4242 453 4245 536
rect 4250 523 4253 613
rect 4258 533 4261 546
rect 4218 443 4229 446
rect 4226 413 4229 443
rect 4266 426 4269 526
rect 4290 513 4293 546
rect 4298 516 4301 536
rect 4306 526 4309 693
rect 4330 636 4333 713
rect 4322 633 4333 636
rect 4314 533 4317 546
rect 4306 523 4317 526
rect 4298 513 4309 516
rect 4306 496 4309 513
rect 4298 493 4309 496
rect 4298 436 4301 493
rect 4298 433 4309 436
rect 4262 423 4269 426
rect 4226 393 4229 406
rect 4250 366 4253 416
rect 4262 376 4265 423
rect 4274 393 4277 416
rect 4306 413 4309 433
rect 4314 413 4317 523
rect 4262 373 4269 376
rect 4242 363 4253 366
rect 4178 323 4181 336
rect 4138 143 4141 216
rect 4162 193 4165 216
rect 4202 213 4205 336
rect 4226 323 4229 346
rect 4242 286 4245 363
rect 4242 283 4253 286
rect 4266 283 4269 373
rect 4218 206 4221 216
rect 4226 213 4229 226
rect 4250 213 4253 283
rect 4274 276 4277 366
rect 4322 363 4325 633
rect 4330 533 4333 546
rect 4338 523 4341 616
rect 4330 383 4333 456
rect 4346 453 4349 536
rect 4362 426 4365 736
rect 4378 703 4381 816
rect 4386 803 4389 923
rect 4394 713 4397 816
rect 4410 813 4413 846
rect 4418 823 4421 933
rect 4426 913 4429 926
rect 4402 766 4405 806
rect 4402 763 4409 766
rect 4406 706 4409 763
rect 4402 703 4409 706
rect 4378 603 4397 606
rect 4378 523 4381 603
rect 4402 566 4405 703
rect 4418 686 4421 736
rect 4434 733 4437 926
rect 4442 923 4445 1026
rect 4450 993 4453 1223
rect 4458 983 4461 1216
rect 4466 1213 4469 1406
rect 4474 1343 4477 1423
rect 4482 1383 4485 1406
rect 4490 1393 4493 1443
rect 4474 1296 4477 1336
rect 4482 1323 4485 1336
rect 4498 1333 4501 1426
rect 4506 1363 4509 1536
rect 4514 1413 4517 1536
rect 4522 1533 4525 1606
rect 4530 1603 4533 1616
rect 4538 1593 4541 1633
rect 4546 1556 4549 1853
rect 4562 1793 4565 1816
rect 4570 1786 4573 1883
rect 4594 1843 4597 1926
rect 4618 1833 4621 2016
rect 4626 2003 4629 2026
rect 4634 2003 4653 2006
rect 4666 2003 4669 2123
rect 4690 2013 4693 2036
rect 4634 1923 4637 2003
rect 4738 1996 4741 2256
rect 4754 2163 4757 2313
rect 4778 2216 4781 2513
rect 4770 2213 4781 2216
rect 4770 2116 4773 2213
rect 4786 2123 4789 2206
rect 4770 2113 4781 2116
rect 4746 2013 4749 2026
rect 4738 1993 4749 1996
rect 4666 1886 4669 1926
rect 4650 1883 4669 1886
rect 4562 1783 4573 1786
rect 4554 1713 4557 1736
rect 4538 1553 4549 1556
rect 4522 1423 4525 1436
rect 4538 1416 4541 1553
rect 4546 1533 4549 1546
rect 4554 1423 4557 1646
rect 4562 1633 4565 1783
rect 4610 1776 4613 1816
rect 4610 1773 4617 1776
rect 4626 1773 4629 1826
rect 4534 1413 4541 1416
rect 4474 1293 4485 1296
rect 4482 1236 4485 1293
rect 4474 1233 4485 1236
rect 4474 1203 4477 1233
rect 4466 1023 4469 1196
rect 4482 1166 4485 1216
rect 4498 1203 4501 1326
rect 4522 1323 4525 1396
rect 4534 1346 4537 1413
rect 4534 1343 4541 1346
rect 4482 1163 4489 1166
rect 4486 1106 4489 1163
rect 4506 1136 4509 1216
rect 4514 1203 4517 1226
rect 4522 1213 4525 1256
rect 4506 1133 4513 1136
rect 4482 1103 4489 1106
rect 4482 1086 4485 1103
rect 4474 1083 4485 1086
rect 4450 913 4453 936
rect 4458 923 4461 956
rect 4466 933 4469 1016
rect 4474 916 4477 1083
rect 4498 1036 4501 1126
rect 4510 1036 4513 1133
rect 4490 1033 4501 1036
rect 4506 1033 4513 1036
rect 4482 973 4485 1016
rect 4490 1003 4493 1033
rect 4498 1013 4501 1026
rect 4506 1003 4509 1033
rect 4482 926 4485 936
rect 4482 923 4493 926
rect 4458 913 4477 916
rect 4442 793 4445 806
rect 4450 803 4453 816
rect 4458 803 4461 913
rect 4482 893 4485 916
rect 4490 863 4493 923
rect 4466 813 4469 836
rect 4474 783 4477 806
rect 4482 746 4485 806
rect 4466 733 4469 746
rect 4474 743 4485 746
rect 4426 713 4429 726
rect 4442 703 4445 726
rect 4418 683 4429 686
rect 4394 563 4405 566
rect 4394 546 4397 563
rect 4426 556 4429 683
rect 4474 613 4477 743
rect 4482 723 4485 736
rect 4490 723 4493 836
rect 4498 733 4501 996
rect 4506 813 4509 986
rect 4514 893 4517 1016
rect 4506 723 4509 806
rect 4514 796 4517 816
rect 4522 803 4525 1206
rect 4530 1203 4533 1326
rect 4538 1323 4541 1343
rect 4546 1306 4549 1406
rect 4554 1403 4557 1416
rect 4562 1333 4565 1536
rect 4570 1533 4573 1736
rect 4578 1643 4581 1726
rect 4586 1713 4589 1726
rect 4578 1526 4581 1636
rect 4594 1603 4597 1736
rect 4602 1733 4605 1756
rect 4614 1726 4617 1773
rect 4642 1746 4645 1836
rect 4650 1803 4653 1883
rect 4658 1763 4661 1816
rect 4666 1783 4669 1806
rect 4682 1793 4685 1826
rect 4714 1823 4717 1936
rect 4746 1916 4749 1993
rect 4738 1913 4749 1916
rect 4738 1893 4741 1913
rect 4634 1743 4645 1746
rect 4610 1723 4617 1726
rect 4586 1533 4589 1556
rect 4594 1533 4597 1596
rect 4570 1523 4581 1526
rect 4602 1523 4605 1616
rect 4610 1613 4613 1723
rect 4610 1543 4613 1606
rect 4570 1436 4573 1523
rect 4610 1506 4613 1536
rect 4602 1503 4613 1506
rect 4602 1436 4605 1503
rect 4570 1433 4581 1436
rect 4570 1366 4573 1426
rect 4578 1386 4581 1433
rect 4586 1406 4589 1436
rect 4602 1433 4613 1436
rect 4610 1416 4613 1433
rect 4594 1413 4613 1416
rect 4618 1416 4621 1636
rect 4626 1603 4629 1726
rect 4634 1593 4637 1743
rect 4626 1533 4629 1556
rect 4634 1516 4637 1546
rect 4630 1513 4637 1516
rect 4630 1436 4633 1513
rect 4630 1433 4637 1436
rect 4618 1413 4629 1416
rect 4634 1413 4637 1433
rect 4586 1403 4605 1406
rect 4578 1383 4589 1386
rect 4570 1363 4577 1366
rect 4542 1303 4549 1306
rect 4542 1236 4545 1303
rect 4542 1233 4549 1236
rect 4538 1186 4541 1216
rect 4546 1213 4549 1233
rect 4554 1206 4557 1276
rect 4530 1183 4541 1186
rect 4546 1203 4557 1206
rect 4562 1203 4565 1326
rect 4574 1256 4577 1363
rect 4570 1253 4577 1256
rect 4546 1183 4549 1203
rect 4530 1133 4533 1183
rect 4538 1023 4541 1166
rect 4546 1106 4549 1136
rect 4570 1126 4573 1253
rect 4586 1236 4589 1383
rect 4602 1346 4605 1403
rect 4578 1233 4589 1236
rect 4598 1343 4605 1346
rect 4598 1236 4601 1343
rect 4618 1336 4621 1406
rect 4610 1333 4621 1336
rect 4598 1233 4605 1236
rect 4578 1163 4581 1233
rect 4586 1193 4589 1206
rect 4578 1133 4581 1156
rect 4586 1133 4589 1146
rect 4570 1123 4581 1126
rect 4578 1106 4581 1123
rect 4586 1113 4589 1126
rect 4594 1106 4597 1216
rect 4546 1103 4557 1106
rect 4554 1046 4557 1103
rect 4546 1043 4557 1046
rect 4570 1103 4581 1106
rect 4586 1103 4597 1106
rect 4570 1046 4573 1103
rect 4570 1043 4581 1046
rect 4546 1013 4549 1043
rect 4530 906 4533 1006
rect 4554 1003 4557 1016
rect 4562 1013 4565 1026
rect 4578 1013 4581 1043
rect 4586 1006 4589 1103
rect 4538 923 4541 936
rect 4546 923 4549 946
rect 4562 936 4565 1006
rect 4570 943 4573 1006
rect 4578 1003 4589 1006
rect 4530 903 4541 906
rect 4538 846 4541 903
rect 4554 893 4557 936
rect 4562 933 4573 936
rect 4562 913 4565 926
rect 4578 906 4581 1003
rect 4594 953 4597 1016
rect 4602 946 4605 1233
rect 4610 983 4613 1333
rect 4618 1203 4621 1326
rect 4618 1006 4621 1136
rect 4626 1116 4629 1413
rect 4634 1273 4637 1406
rect 4642 1403 4645 1734
rect 4650 1506 4653 1746
rect 4658 1633 4661 1736
rect 4674 1733 4677 1746
rect 4666 1683 4669 1726
rect 4682 1643 4685 1786
rect 4698 1746 4701 1766
rect 4694 1743 4701 1746
rect 4694 1676 4697 1743
rect 4714 1733 4717 1816
rect 4762 1813 4765 1826
rect 4730 1736 4733 1776
rect 4730 1733 4741 1736
rect 4706 1683 4709 1726
rect 4722 1703 4725 1726
rect 4730 1713 4733 1726
rect 4738 1723 4741 1733
rect 4746 1733 4765 1736
rect 4694 1673 4701 1676
rect 4698 1646 4701 1673
rect 4698 1643 4705 1646
rect 4666 1543 4669 1616
rect 4690 1613 4693 1636
rect 4702 1586 4705 1643
rect 4730 1626 4733 1646
rect 4730 1623 4737 1626
rect 4698 1583 4705 1586
rect 4698 1563 4701 1583
rect 4658 1533 4669 1536
rect 4666 1513 4669 1526
rect 4674 1523 4677 1536
rect 4650 1503 4657 1506
rect 4654 1446 4657 1503
rect 4650 1443 4657 1446
rect 4650 1383 4653 1443
rect 4666 1403 4669 1426
rect 4690 1423 4693 1546
rect 4714 1523 4717 1536
rect 4722 1513 4725 1566
rect 4734 1506 4737 1623
rect 4746 1613 4749 1733
rect 4754 1613 4757 1646
rect 4730 1503 4737 1506
rect 4730 1456 4733 1503
rect 4730 1453 4737 1456
rect 4658 1216 4661 1346
rect 4666 1333 4669 1396
rect 4690 1393 4693 1416
rect 4674 1313 4677 1326
rect 4682 1233 4685 1386
rect 4734 1376 4737 1453
rect 4746 1406 4749 1416
rect 4762 1413 4765 1726
rect 4770 1703 4773 1816
rect 4778 1786 4781 2113
rect 4786 1803 4789 1826
rect 4778 1783 4789 1786
rect 4786 1576 4789 1783
rect 4778 1573 4789 1576
rect 4770 1513 4773 1526
rect 4746 1403 4765 1406
rect 4730 1373 4737 1376
rect 4690 1316 4693 1336
rect 4730 1333 4733 1373
rect 4770 1343 4773 1416
rect 4690 1313 4709 1316
rect 4706 1226 4709 1313
rect 4730 1236 4733 1256
rect 4690 1223 4709 1226
rect 4722 1233 4733 1236
rect 4634 1133 4637 1206
rect 4626 1113 4633 1116
rect 4630 1046 4633 1113
rect 4626 1043 4633 1046
rect 4642 1043 4645 1216
rect 4658 1213 4669 1216
rect 4650 1153 4653 1206
rect 4666 1146 4669 1213
rect 4658 1143 4669 1146
rect 4658 1066 4661 1143
rect 4650 1063 4661 1066
rect 4626 1023 4629 1043
rect 4618 1003 4629 1006
rect 4594 943 4605 946
rect 4574 903 4581 906
rect 4530 843 4541 846
rect 4530 823 4533 843
rect 4574 836 4577 903
rect 4574 833 4581 836
rect 4530 813 4541 816
rect 4514 793 4525 796
rect 4514 616 4517 746
rect 4522 703 4525 793
rect 4530 713 4533 813
rect 4538 766 4541 806
rect 4538 763 4545 766
rect 4542 706 4545 763
rect 4562 726 4565 826
rect 4578 813 4581 833
rect 4570 733 4573 746
rect 4586 733 4589 926
rect 4594 883 4597 943
rect 4602 803 4605 936
rect 4610 903 4613 936
rect 4626 896 4629 1003
rect 4642 993 4645 1006
rect 4650 1003 4653 1063
rect 4618 893 4629 896
rect 4618 793 4621 893
rect 4538 703 4545 706
rect 4538 623 4541 703
rect 4514 613 4525 616
rect 4418 553 4429 556
rect 4390 543 4397 546
rect 4346 423 4365 426
rect 4282 333 4301 336
rect 4282 323 4285 333
rect 4290 313 4293 326
rect 4314 323 4317 336
rect 4266 273 4277 276
rect 4266 213 4269 273
rect 4282 213 4285 226
rect 4322 213 4325 286
rect 4346 213 4349 423
rect 4378 416 4381 516
rect 4390 486 4393 543
rect 4410 523 4413 546
rect 4390 483 4397 486
rect 4354 393 4357 406
rect 4362 373 4365 416
rect 4370 413 4381 416
rect 4370 403 4373 413
rect 4378 383 4381 406
rect 4394 383 4397 483
rect 4418 416 4421 553
rect 4458 523 4461 536
rect 4410 413 4421 416
rect 4362 323 4365 346
rect 4410 323 4413 413
rect 4426 353 4429 416
rect 4434 393 4437 406
rect 4450 403 4453 456
rect 4458 413 4461 436
rect 4474 403 4477 526
rect 4506 523 4509 606
rect 4514 453 4517 606
rect 4522 433 4525 613
rect 4530 566 4533 606
rect 4538 573 4541 616
rect 4554 613 4557 726
rect 4562 723 4569 726
rect 4566 626 4569 723
rect 4566 623 4573 626
rect 4530 563 4541 566
rect 4538 523 4541 563
rect 4546 513 4549 606
rect 4554 593 4557 606
rect 4570 603 4573 623
rect 4578 613 4581 716
rect 4594 713 4597 726
rect 4602 636 4605 736
rect 4610 733 4613 746
rect 4618 716 4621 786
rect 4614 713 4621 716
rect 4614 656 4617 713
rect 4614 653 4621 656
rect 4602 633 4613 636
rect 4586 603 4589 616
rect 4594 593 4597 606
rect 4554 506 4557 576
rect 4586 523 4589 536
rect 4546 503 4557 506
rect 4498 393 4501 416
rect 4434 356 4437 376
rect 4434 353 4441 356
rect 4426 306 4429 336
rect 4418 303 4429 306
rect 4418 226 4421 303
rect 4438 296 4441 353
rect 4434 293 4441 296
rect 4418 223 4429 226
rect 4218 203 4237 206
rect 4242 173 4245 206
rect 4258 166 4261 206
rect 4282 193 4285 206
rect 4250 163 4261 166
rect 4058 113 4061 136
rect 4082 123 4101 126
rect 4114 123 4117 136
rect 4162 133 4165 156
rect 4202 133 4205 156
rect 4250 123 4253 163
rect 4298 123 4301 206
rect 4306 193 4309 206
rect 4314 133 4317 156
rect 4330 146 4333 206
rect 4346 173 4349 206
rect 4330 143 4341 146
rect 4338 123 4341 143
rect 4394 123 4397 206
rect 4402 193 4405 206
rect 4426 173 4429 223
rect 4434 213 4437 293
rect 4450 213 4453 386
rect 4458 333 4461 346
rect 4466 323 4469 356
rect 4442 146 4445 206
rect 4458 173 4461 206
rect 4474 193 4477 386
rect 4530 306 4533 326
rect 4522 303 4533 306
rect 4522 226 4525 303
rect 4522 223 4533 226
rect 4426 133 4429 146
rect 4442 143 4453 146
rect 4450 123 4453 143
rect 4506 123 4509 206
rect 4514 193 4517 206
rect 4530 133 4533 223
rect 4546 213 4549 503
rect 4602 496 4605 626
rect 4598 493 4605 496
rect 4554 406 4557 416
rect 4562 413 4565 436
rect 4598 426 4601 493
rect 4586 413 4589 426
rect 4598 423 4605 426
rect 4554 403 4573 406
rect 4562 356 4565 396
rect 4578 383 4581 406
rect 4558 353 4565 356
rect 4558 306 4561 353
rect 4594 346 4597 406
rect 4602 393 4605 423
rect 4610 413 4613 633
rect 4618 523 4621 653
rect 4626 506 4629 806
rect 4634 733 4637 836
rect 4642 803 4645 986
rect 4658 963 4661 1026
rect 4674 1013 4677 1046
rect 4658 816 4661 936
rect 4666 923 4669 1006
rect 4682 993 4685 1006
rect 4690 1003 4693 1223
rect 4722 1176 4725 1233
rect 4738 1186 4741 1316
rect 4746 1253 4749 1326
rect 4738 1183 4745 1186
rect 4706 996 4709 1176
rect 4722 1173 4733 1176
rect 4730 1076 4733 1173
rect 4742 1126 4745 1183
rect 4690 993 4709 996
rect 4722 1073 4733 1076
rect 4738 1123 4745 1126
rect 4754 1123 4757 1336
rect 4762 1213 4765 1326
rect 4690 933 4693 993
rect 4722 916 4725 1073
rect 4738 973 4741 1123
rect 4746 966 4749 1006
rect 4754 993 4757 1016
rect 4770 1003 4773 1336
rect 4778 1316 4781 1573
rect 4786 1513 4789 1536
rect 4794 1523 4797 1556
rect 4786 1333 4789 1416
rect 4778 1313 4789 1316
rect 4786 1226 4789 1313
rect 4778 1223 4789 1226
rect 4778 1106 4781 1223
rect 4786 1123 4789 1206
rect 4778 1103 4789 1106
rect 4786 1016 4789 1103
rect 4778 1013 4789 1016
rect 4738 963 4749 966
rect 4738 923 4741 963
rect 4754 956 4757 976
rect 4754 953 4761 956
rect 4722 913 4733 916
rect 4634 613 4637 726
rect 4642 706 4645 796
rect 4650 723 4653 816
rect 4658 813 4669 816
rect 4666 796 4669 813
rect 4658 793 4669 796
rect 4658 733 4661 793
rect 4674 783 4677 896
rect 4730 826 4733 913
rect 4758 886 4761 953
rect 4770 913 4773 926
rect 4754 883 4761 886
rect 4754 856 4757 883
rect 4750 853 4757 856
rect 4730 823 4741 826
rect 4642 703 4653 706
rect 4650 646 4653 703
rect 4642 643 4653 646
rect 4642 603 4645 643
rect 4666 626 4669 736
rect 4674 723 4677 736
rect 4682 706 4685 746
rect 4706 736 4709 806
rect 4678 703 4685 706
rect 4678 636 4681 703
rect 4678 633 4685 636
rect 4650 623 4669 626
rect 4650 613 4653 623
rect 4658 603 4661 616
rect 4666 596 4669 616
rect 4682 613 4685 633
rect 4658 593 4669 596
rect 4622 503 4629 506
rect 4622 436 4625 503
rect 4622 433 4629 436
rect 4626 413 4629 433
rect 4634 413 4637 526
rect 4642 483 4645 536
rect 4650 486 4653 586
rect 4658 523 4661 593
rect 4666 533 4669 546
rect 4674 506 4677 536
rect 4670 503 4677 506
rect 4650 483 4661 486
rect 4610 373 4613 406
rect 4650 386 4653 406
rect 4658 403 4661 483
rect 4670 416 4673 503
rect 4682 446 4685 606
rect 4690 583 4693 736
rect 4698 733 4709 736
rect 4730 733 4733 816
rect 4698 466 4701 733
rect 4706 696 4709 726
rect 4738 706 4741 823
rect 4750 796 4753 853
rect 4778 826 4781 1013
rect 4786 913 4789 936
rect 4794 923 4797 996
rect 4774 823 4781 826
rect 4750 793 4757 796
rect 4754 776 4757 793
rect 4774 776 4777 823
rect 4754 773 4765 776
rect 4774 773 4781 776
rect 4762 756 4765 773
rect 4762 753 4769 756
rect 4730 703 4741 706
rect 4706 693 4717 696
rect 4714 646 4717 693
rect 4706 643 4717 646
rect 4706 593 4709 643
rect 4730 626 4733 703
rect 4722 623 4733 626
rect 4722 566 4725 623
rect 4738 586 4741 616
rect 4746 603 4749 736
rect 4754 713 4757 726
rect 4766 706 4769 753
rect 4778 716 4781 773
rect 4786 733 4789 816
rect 4778 713 4789 716
rect 4762 703 4769 706
rect 4738 583 4745 586
rect 4722 563 4733 566
rect 4722 523 4725 546
rect 4698 463 4709 466
rect 4682 443 4693 446
rect 4666 413 4673 416
rect 4682 413 4685 426
rect 4666 386 4669 413
rect 4674 393 4677 406
rect 4650 383 4661 386
rect 4666 383 4677 386
rect 4594 343 4605 346
rect 4578 323 4581 336
rect 4602 323 4605 343
rect 4658 323 4661 383
rect 4666 333 4669 376
rect 4674 326 4677 383
rect 4666 323 4677 326
rect 4666 306 4669 323
rect 4682 306 4685 406
rect 4690 403 4693 443
rect 4706 403 4709 463
rect 4730 423 4733 563
rect 4742 446 4745 583
rect 4762 533 4765 703
rect 4786 626 4789 713
rect 4778 623 4789 626
rect 4778 606 4781 623
rect 4774 603 4781 606
rect 4738 443 4745 446
rect 4730 393 4733 416
rect 4558 303 4565 306
rect 4562 213 4565 303
rect 4658 303 4669 306
rect 4678 303 4685 306
rect 4658 236 4661 303
rect 4678 236 4681 303
rect 4658 233 4669 236
rect 4678 233 4685 236
rect 4554 123 4557 206
rect 4570 173 4573 206
rect 4586 193 4589 216
rect 4666 213 4669 233
rect 4610 123 4613 206
rect 4626 173 4629 206
rect 4642 133 4645 146
rect 4674 123 4677 206
rect 3922 103 3941 106
rect 4042 103 4061 106
rect 3938 0 3941 103
rect 4058 0 4061 103
rect 4082 0 4085 116
rect 4098 76 4101 123
rect 4682 113 4685 233
rect 4690 173 4693 336
rect 4698 323 4701 336
rect 4706 223 4709 336
rect 4714 323 4717 376
rect 4722 333 4725 386
rect 4738 323 4741 443
rect 4746 373 4749 426
rect 4774 406 4777 603
rect 4786 523 4789 606
rect 4786 413 4789 486
rect 4774 403 4781 406
rect 4778 346 4781 403
rect 4770 343 4781 346
rect 4770 266 4773 343
rect 4770 263 4781 266
rect 4730 213 4733 226
rect 4706 143 4709 206
rect 4778 203 4781 263
rect 4786 213 4789 336
rect 4722 133 4741 136
rect 4722 123 4725 133
rect 4730 113 4733 126
rect 4098 73 4109 76
rect 4106 16 4109 73
rect 4809 37 4829 4703
rect 4098 13 4109 16
rect 4833 13 4853 4727
rect 4098 0 4101 13
<< metal3 >>
rect 1649 4732 3126 4737
rect 1169 4702 2798 4707
rect 2017 4682 2478 4687
rect 1865 4672 2006 4677
rect 2001 4667 2006 4672
rect 2489 4672 3166 4677
rect 2489 4667 2494 4672
rect 2001 4662 2494 4667
rect 1569 4642 2878 4647
rect 3569 4642 3662 4647
rect 3569 4637 3574 4642
rect 3481 4632 3574 4637
rect 3657 4637 3662 4642
rect 3657 4632 3822 4637
rect 545 4622 590 4627
rect 689 4622 734 4627
rect 1025 4622 1070 4627
rect 1801 4622 1846 4627
rect 2169 4622 2214 4627
rect 2537 4622 2582 4627
rect 2673 4622 2718 4627
rect 2849 4622 2894 4627
rect 3617 4622 3646 4627
rect 4473 4622 4550 4627
rect 4473 4617 4478 4622
rect 3585 4612 3958 4617
rect 4449 4612 4478 4617
rect 4545 4617 4550 4622
rect 4545 4612 4686 4617
rect 377 4602 430 4607
rect 857 4602 886 4607
rect 1369 4602 1446 4607
rect 3033 4602 3102 4607
rect 3161 4602 3246 4607
rect 3265 4602 3310 4607
rect 3433 4602 3518 4607
rect 3729 4602 3758 4607
rect 3937 4602 4006 4607
rect 4081 4602 4126 4607
rect 4497 4602 4534 4607
rect 3161 4597 3166 4602
rect 89 4592 710 4597
rect 809 4592 838 4597
rect 897 4592 1262 4597
rect 1345 4592 1590 4597
rect 1793 4592 1846 4597
rect 1953 4592 2030 4597
rect 2185 4592 2502 4597
rect 2553 4592 2710 4597
rect 2729 4592 2822 4597
rect 2841 4592 2918 4597
rect 2985 4592 3014 4597
rect 3105 4592 3166 4597
rect 3241 4597 3246 4602
rect 3241 4592 3286 4597
rect 3457 4592 3486 4597
rect 3529 4592 3638 4597
rect 4049 4592 4118 4597
rect 4217 4592 4454 4597
rect 4681 4592 4710 4597
rect 833 4587 902 4592
rect 1953 4587 1958 4592
rect 1817 4582 1958 4587
rect 2025 4587 2030 4592
rect 2705 4587 2710 4592
rect 2841 4587 2846 4592
rect 2025 4582 2054 4587
rect 2705 4582 2846 4587
rect 2913 4587 2918 4592
rect 3009 4587 3110 4592
rect 2913 4582 2942 4587
rect 3129 4582 3590 4587
rect 3625 4582 3790 4587
rect 3809 4582 3846 4587
rect 4329 4582 4366 4587
rect 1513 4572 1774 4577
rect 1513 4567 1518 4572
rect 449 4562 518 4567
rect 537 4562 558 4567
rect 961 4562 1038 4567
rect 449 4557 454 4562
rect 273 4552 454 4557
rect 513 4557 518 4562
rect 961 4557 966 4562
rect 513 4552 558 4557
rect 937 4552 966 4557
rect 1033 4557 1038 4562
rect 1289 4562 1470 4567
rect 1489 4562 1518 4567
rect 1769 4567 1774 4572
rect 2121 4572 2214 4577
rect 2121 4567 2126 4572
rect 1769 4562 1870 4567
rect 1897 4562 2126 4567
rect 2209 4567 2214 4572
rect 2273 4572 2446 4577
rect 2273 4567 2278 4572
rect 2209 4562 2238 4567
rect 2249 4562 2278 4567
rect 2441 4567 2446 4572
rect 2529 4572 2654 4577
rect 2673 4572 2782 4577
rect 2801 4572 2846 4577
rect 2873 4572 3286 4577
rect 3505 4572 3630 4577
rect 3649 4572 3830 4577
rect 3865 4572 4126 4577
rect 2529 4567 2534 4572
rect 2441 4562 2534 4567
rect 2649 4567 2654 4572
rect 2801 4567 2806 4572
rect 3865 4567 3870 4572
rect 2649 4562 2806 4567
rect 2825 4562 2982 4567
rect 3425 4562 3870 4567
rect 4121 4567 4126 4572
rect 4385 4572 4550 4577
rect 4385 4567 4390 4572
rect 4121 4562 4390 4567
rect 4545 4567 4550 4572
rect 4545 4562 4574 4567
rect 4593 4562 4670 4567
rect 1289 4557 1294 4562
rect 1033 4552 1062 4557
rect 1265 4552 1294 4557
rect 1465 4557 1470 4562
rect 3121 4557 3262 4562
rect 3889 4557 4006 4562
rect 4593 4557 4598 4562
rect 1465 4552 1662 4557
rect 2137 4552 2358 4557
rect 2377 4552 2430 4557
rect 2425 4547 2430 4552
rect 2545 4552 2758 4557
rect 2849 4552 2894 4557
rect 2545 4547 2550 4552
rect 2889 4547 2894 4552
rect 2977 4552 3126 4557
rect 3257 4552 3486 4557
rect 3601 4552 3894 4557
rect 4001 4552 4110 4557
rect 4345 4552 4550 4557
rect 4561 4552 4598 4557
rect 4665 4557 4670 4562
rect 4665 4552 4782 4557
rect 2977 4547 2982 4552
rect 169 4542 190 4547
rect 393 4542 494 4547
rect 681 4542 782 4547
rect 1001 4542 1086 4547
rect 1105 4542 1246 4547
rect 1305 4542 1510 4547
rect 1689 4542 1822 4547
rect 1833 4542 1910 4547
rect 1937 4542 2030 4547
rect 1105 4537 1110 4542
rect 529 4532 654 4537
rect 713 4532 950 4537
rect 1009 4532 1110 4537
rect 1241 4537 1246 4542
rect 1241 4532 1270 4537
rect 1401 4532 1534 4537
rect 1593 4532 1678 4537
rect 1897 4532 1974 4537
rect 2057 4532 2134 4537
rect 1265 4527 1406 4532
rect 1673 4527 1902 4532
rect 177 4522 230 4527
rect 265 4522 310 4527
rect 793 4522 838 4527
rect 913 4522 1094 4527
rect 1113 4522 1214 4527
rect 1425 4522 1654 4527
rect 1921 4522 2070 4527
rect 2161 4522 2166 4547
rect 2225 4542 2270 4547
rect 2425 4542 2550 4547
rect 2569 4542 2638 4547
rect 2681 4542 2718 4547
rect 2761 4542 2862 4547
rect 2889 4542 2982 4547
rect 3001 4542 3030 4547
rect 3137 4542 3246 4547
rect 3529 4542 3654 4547
rect 3729 4542 3934 4547
rect 3953 4542 4310 4547
rect 4337 4542 4430 4547
rect 4545 4542 4742 4547
rect 3025 4537 3142 4542
rect 2193 4532 2406 4537
rect 2585 4532 2750 4537
rect 2793 4532 2870 4537
rect 3161 4532 3278 4537
rect 3289 4532 3790 4537
rect 3897 4532 4094 4537
rect 4321 4532 4446 4537
rect 4521 4532 4598 4537
rect 3785 4527 3902 4532
rect 2521 4522 2606 4527
rect 2641 4522 2686 4527
rect 2697 4522 2790 4527
rect 3097 4522 3190 4527
rect 3201 4522 3766 4527
rect 3921 4522 4038 4527
rect 4097 4522 4198 4527
rect 4265 4522 4350 4527
rect 4657 4522 4702 4527
rect 3201 4517 3206 4522
rect 3761 4517 3766 4522
rect 169 4512 198 4517
rect 193 4507 198 4512
rect 273 4512 326 4517
rect 369 4512 406 4517
rect 489 4512 718 4517
rect 777 4512 822 4517
rect 937 4512 1078 4517
rect 1137 4512 1198 4517
rect 1257 4512 1438 4517
rect 1481 4512 1630 4517
rect 1737 4512 1782 4517
rect 1857 4512 2150 4517
rect 2241 4512 2350 4517
rect 2433 4512 2510 4517
rect 2569 4512 2598 4517
rect 2841 4512 2934 4517
rect 2969 4512 3094 4517
rect 3153 4512 3206 4517
rect 3257 4512 3286 4517
rect 3401 4512 3542 4517
rect 3641 4512 3686 4517
rect 3761 4512 3966 4517
rect 4001 4512 4094 4517
rect 4225 4512 4294 4517
rect 4409 4512 4558 4517
rect 4673 4512 4726 4517
rect 273 4507 278 4512
rect 193 4502 278 4507
rect 321 4507 326 4512
rect 1073 4507 1078 4512
rect 2505 4507 2574 4512
rect 321 4502 510 4507
rect 1073 4502 1158 4507
rect 1233 4502 1286 4507
rect 2009 4502 2158 4507
rect 2177 4502 2318 4507
rect 2937 4502 3022 4507
rect 3569 4502 3758 4507
rect 529 4497 718 4502
rect 473 4492 534 4497
rect 713 4492 1030 4497
rect 1065 4492 1166 4497
rect 1889 4492 1998 4497
rect 2057 4492 2086 4497
rect 2265 4492 2390 4497
rect 2409 4492 2654 4497
rect 2777 4492 2926 4497
rect 3033 4492 3422 4497
rect 3473 4492 3550 4497
rect 3961 4492 4630 4497
rect 1201 4487 1294 4492
rect 1993 4487 2062 4492
rect 2409 4487 2414 4492
rect 465 4482 702 4487
rect 1065 4482 1206 4487
rect 1289 4482 1814 4487
rect 2153 4482 2414 4487
rect 2649 4487 2654 4492
rect 2921 4487 3038 4492
rect 3473 4487 3478 4492
rect 3545 4487 3630 4492
rect 2649 4482 2678 4487
rect 3433 4482 3478 4487
rect 3625 4482 3950 4487
rect 721 4477 870 4482
rect 961 4477 1070 4482
rect 1809 4477 1814 4482
rect 2433 4477 2542 4482
rect 3945 4477 3950 4482
rect 4369 4482 4398 4487
rect 449 4472 486 4477
rect 609 4472 726 4477
rect 865 4472 966 4477
rect 1089 4472 1134 4477
rect 1217 4472 1278 4477
rect 1809 4472 1918 4477
rect 1129 4467 1222 4472
rect 1913 4467 1918 4472
rect 2057 4472 2438 4477
rect 2537 4472 2718 4477
rect 2961 4472 3014 4477
rect 3033 4472 3278 4477
rect 3489 4472 3518 4477
rect 3713 4472 3742 4477
rect 3945 4472 4222 4477
rect 2057 4467 2062 4472
rect 3033 4467 3038 4472
rect 585 4462 1110 4467
rect 1105 4457 1110 4462
rect 1241 4462 1798 4467
rect 1241 4457 1246 4462
rect 481 4452 1014 4457
rect 1105 4452 1246 4457
rect 1793 4457 1798 4462
rect 1865 4462 1894 4467
rect 1913 4462 2062 4467
rect 2081 4462 2110 4467
rect 1865 4457 1870 4462
rect 1793 4452 1870 4457
rect 2105 4457 2110 4462
rect 2233 4462 2438 4467
rect 2497 4462 2526 4467
rect 2729 4462 3038 4467
rect 3273 4467 3278 4472
rect 3513 4467 3614 4472
rect 3713 4467 3718 4472
rect 4217 4467 4222 4472
rect 4369 4467 4374 4482
rect 3273 4462 3422 4467
rect 3609 4462 3718 4467
rect 3753 4462 3838 4467
rect 4217 4462 4374 4467
rect 4433 4462 4590 4467
rect 2233 4457 2238 4462
rect 2521 4457 2734 4462
rect 3057 4457 3150 4462
rect 2105 4452 2238 4457
rect 2313 4452 2430 4457
rect 2993 4452 3062 4457
rect 3145 4452 3262 4457
rect 3505 4452 3590 4457
rect 3857 4452 4110 4457
rect 3857 4447 3862 4452
rect 217 4442 462 4447
rect 753 4442 886 4447
rect 1265 4442 1302 4447
rect 1321 4442 1502 4447
rect 2545 4442 2622 4447
rect 457 4437 662 4442
rect 937 4437 1086 4442
rect 1265 4437 1270 4442
rect 1321 4437 1326 4442
rect 161 4432 270 4437
rect 657 4432 782 4437
rect 777 4427 782 4432
rect 841 4432 942 4437
rect 1081 4432 1110 4437
rect 1233 4432 1270 4437
rect 1289 4432 1326 4437
rect 1497 4437 1502 4442
rect 2281 4437 2350 4442
rect 2401 4437 2478 4442
rect 2545 4437 2550 4442
rect 1497 4432 1694 4437
rect 1809 4432 1838 4437
rect 2257 4432 2286 4437
rect 2345 4432 2406 4437
rect 2473 4432 2550 4437
rect 2617 4437 2622 4442
rect 2681 4442 2758 4447
rect 2897 4442 3134 4447
rect 3273 4442 3430 4447
rect 3497 4442 3526 4447
rect 3601 4442 3862 4447
rect 4105 4447 4110 4452
rect 4105 4442 4198 4447
rect 2681 4437 2686 4442
rect 2617 4432 2686 4437
rect 2753 4437 2758 4442
rect 3129 4437 3278 4442
rect 3521 4437 3606 4442
rect 2753 4432 2854 4437
rect 2873 4432 3006 4437
rect 3073 4432 3110 4437
rect 3473 4432 3502 4437
rect 841 4427 846 4432
rect 3497 4427 3502 4432
rect 3641 4432 3670 4437
rect 3865 4432 3950 4437
rect 4217 4432 4414 4437
rect 3641 4427 3646 4432
rect 129 4422 174 4427
rect 257 4422 286 4427
rect 353 4422 430 4427
rect 449 4422 646 4427
rect 777 4422 846 4427
rect 953 4422 1310 4427
rect 1321 4422 1486 4427
rect 1625 4422 1710 4427
rect 353 4417 358 4422
rect 121 4412 214 4417
rect 329 4412 358 4417
rect 425 4417 430 4422
rect 1745 4417 1750 4427
rect 1769 4422 1830 4427
rect 1881 4422 1974 4427
rect 1993 4422 2030 4427
rect 2049 4422 2166 4427
rect 2185 4422 2270 4427
rect 2289 4422 2334 4427
rect 2417 4422 2462 4427
rect 2561 4422 2606 4427
rect 2697 4422 2742 4427
rect 2825 4422 2918 4427
rect 2985 4422 3030 4427
rect 3089 4422 3262 4427
rect 3497 4422 3646 4427
rect 3721 4422 3886 4427
rect 3921 4422 3966 4427
rect 4017 4422 4094 4427
rect 4449 4422 4502 4427
rect 4601 4422 4782 4427
rect 1881 4417 1886 4422
rect 425 4412 462 4417
rect 633 4412 662 4417
rect 681 4412 758 4417
rect 889 4412 950 4417
rect 1041 4412 1094 4417
rect 1105 4412 1166 4417
rect 1257 4412 1342 4417
rect 1497 4412 1614 4417
rect 1697 4412 1726 4417
rect 1745 4412 1774 4417
rect 1857 4412 1886 4417
rect 1969 4417 1974 4422
rect 2049 4417 2054 4422
rect 1969 4412 2054 4417
rect 2161 4417 2166 4422
rect 4113 4417 4254 4422
rect 2161 4412 2254 4417
rect 481 4407 614 4412
rect 681 4407 686 4412
rect 257 4402 486 4407
rect 609 4402 686 4407
rect 753 4407 758 4412
rect 1161 4407 1262 4412
rect 1337 4407 1502 4412
rect 1609 4407 1702 4412
rect 1769 4407 1862 4412
rect 2249 4407 2254 4412
rect 2345 4412 2406 4417
rect 2345 4407 2350 4412
rect 753 4402 798 4407
rect 1049 4402 1078 4407
rect 1089 4402 1142 4407
rect 1281 4402 1318 4407
rect 1985 4402 2030 4407
rect 2041 4402 2070 4407
rect 2249 4402 2350 4407
rect 2401 4407 2406 4412
rect 2473 4412 2550 4417
rect 2473 4407 2478 4412
rect 2401 4402 2478 4407
rect 2545 4407 2550 4412
rect 2617 4412 2942 4417
rect 2617 4407 2622 4412
rect 2937 4407 2942 4412
rect 3033 4412 3070 4417
rect 3225 4412 3462 4417
rect 3033 4407 3038 4412
rect 2545 4402 2622 4407
rect 2641 4402 2830 4407
rect 833 4397 990 4402
rect 1089 4397 1094 4402
rect 2825 4397 2830 4402
rect 2889 4402 2918 4407
rect 2937 4402 3038 4407
rect 3457 4407 3462 4412
rect 3673 4412 4118 4417
rect 4249 4412 4278 4417
rect 3673 4407 3678 4412
rect 4369 4407 4374 4417
rect 4409 4412 4542 4417
rect 3457 4402 3678 4407
rect 3697 4402 4430 4407
rect 4441 4402 4526 4407
rect 4561 4402 4622 4407
rect 2889 4397 2894 4402
rect 217 4392 246 4397
rect 449 4392 518 4397
rect 545 4392 654 4397
rect 809 4392 838 4397
rect 985 4392 1094 4397
rect 1161 4392 1262 4397
rect 1385 4392 1494 4397
rect 1593 4392 1702 4397
rect 1801 4392 1830 4397
rect 241 4387 366 4392
rect 449 4387 454 4392
rect 361 4382 454 4387
rect 513 4387 518 4392
rect 649 4387 742 4392
rect 809 4387 814 4392
rect 1161 4387 1166 4392
rect 513 4382 574 4387
rect 585 4382 630 4387
rect 737 4382 814 4387
rect 857 4382 974 4387
rect 1097 4382 1166 4387
rect 1257 4387 1262 4392
rect 1825 4387 1830 4392
rect 1897 4392 2022 4397
rect 2033 4392 2230 4397
rect 2825 4392 2894 4397
rect 3081 4392 3166 4397
rect 3265 4392 3350 4397
rect 3729 4392 4014 4397
rect 4113 4392 4142 4397
rect 4161 4392 4254 4397
rect 4273 4392 4462 4397
rect 4609 4392 4694 4397
rect 1897 4387 1902 4392
rect 2681 4387 2782 4392
rect 3265 4387 3270 4392
rect 1257 4382 1302 4387
rect 1825 4382 1902 4387
rect 2273 4382 2326 4387
rect 2345 4382 2622 4387
rect 2657 4382 2686 4387
rect 2777 4382 2806 4387
rect 3057 4382 3270 4387
rect 3345 4387 3350 4392
rect 3345 4382 3406 4387
rect 3945 4382 4422 4387
rect 1977 4377 2254 4382
rect 2345 4377 2350 4382
rect 273 4372 342 4377
rect 273 4367 278 4372
rect 233 4362 278 4367
rect 337 4367 342 4372
rect 649 4372 718 4377
rect 1001 4372 1270 4377
rect 1545 4372 1622 4377
rect 1921 4372 1982 4377
rect 2249 4372 2350 4377
rect 2617 4377 2622 4382
rect 3769 4377 3918 4382
rect 2617 4372 2798 4377
rect 2865 4372 3046 4377
rect 3209 4372 3334 4377
rect 649 4367 654 4372
rect 337 4362 654 4367
rect 713 4367 718 4372
rect 873 4367 982 4372
rect 3041 4367 3046 4372
rect 3113 4367 3214 4372
rect 3329 4367 3334 4372
rect 3417 4372 3774 4377
rect 3913 4372 3942 4377
rect 4169 4372 4606 4377
rect 3417 4367 3422 4372
rect 713 4362 878 4367
rect 977 4362 1350 4367
rect 1345 4357 1350 4362
rect 1361 4362 1502 4367
rect 1993 4362 2262 4367
rect 2385 4362 2438 4367
rect 3041 4362 3118 4367
rect 3233 4362 3310 4367
rect 3329 4362 3422 4367
rect 3785 4362 3894 4367
rect 4009 4362 4086 4367
rect 4129 4362 4446 4367
rect 1361 4357 1366 4362
rect 289 4352 326 4357
rect 889 4352 982 4357
rect 1233 4352 1278 4357
rect 1345 4352 1366 4357
rect 1497 4357 1502 4362
rect 2585 4357 2678 4362
rect 4009 4357 4014 4362
rect 1497 4352 1782 4357
rect 1905 4352 2590 4357
rect 2673 4352 2934 4357
rect 3137 4352 3310 4357
rect 3641 4352 3902 4357
rect 3985 4352 4014 4357
rect 4081 4357 4086 4362
rect 4081 4352 4302 4357
rect 321 4347 326 4352
rect 513 4347 702 4352
rect 889 4347 894 4352
rect 1145 4347 1214 4352
rect 321 4342 518 4347
rect 697 4342 894 4347
rect 913 4342 998 4347
rect 1081 4342 1150 4347
rect 1209 4342 1270 4347
rect 1377 4342 1486 4347
rect 1753 4342 1854 4347
rect 1969 4342 2054 4347
rect 2129 4342 2158 4347
rect 2257 4342 2310 4347
rect 2425 4342 2494 4347
rect 2601 4342 2662 4347
rect 2889 4342 2926 4347
rect 3089 4342 3142 4347
rect 3569 4342 3614 4347
rect 3761 4342 3886 4347
rect 4001 4342 4070 4347
rect 4153 4342 4230 4347
rect 2153 4337 2262 4342
rect 3657 4337 3742 4342
rect 265 4332 302 4337
rect 537 4332 614 4337
rect 1161 4332 1206 4337
rect 1721 4332 1766 4337
rect 2281 4332 2342 4337
rect 2361 4327 2478 4332
rect 2497 4327 2502 4337
rect 2561 4332 2678 4337
rect 2689 4332 2734 4337
rect 3065 4332 3558 4337
rect 3625 4332 3662 4337
rect 3737 4332 4150 4337
rect 4289 4332 4326 4337
rect 4353 4332 4398 4337
rect 409 4322 486 4327
rect 617 4322 678 4327
rect 833 4322 862 4327
rect 897 4322 1014 4327
rect 1025 4322 1078 4327
rect 1313 4322 1470 4327
rect 1513 4322 1598 4327
rect 1009 4317 1014 4322
rect 1513 4317 1518 4322
rect 137 4312 182 4317
rect 505 4312 550 4317
rect 585 4312 614 4317
rect 881 4312 926 4317
rect 1009 4312 1102 4317
rect 1305 4312 1518 4317
rect 1593 4317 1598 4322
rect 1793 4322 2102 4327
rect 2217 4322 2246 4327
rect 2329 4322 2366 4327
rect 2473 4322 2502 4327
rect 2529 4322 2614 4327
rect 2625 4322 2878 4327
rect 2937 4322 2974 4327
rect 3089 4322 3094 4332
rect 3553 4327 3630 4332
rect 3673 4322 4270 4327
rect 4417 4322 4454 4327
rect 1793 4317 1798 4322
rect 1593 4312 1798 4317
rect 2097 4317 2102 4322
rect 2097 4312 2830 4317
rect 3073 4312 3190 4317
rect 3241 4312 3334 4317
rect 3625 4312 4190 4317
rect 4313 4312 4350 4317
rect 4593 4312 4598 4337
rect 169 4302 254 4307
rect 577 4302 638 4307
rect 1113 4302 1174 4307
rect 1329 4302 1430 4307
rect 1529 4302 1582 4307
rect 1809 4302 1950 4307
rect 1993 4302 2086 4307
rect 2297 4302 2358 4307
rect 2473 4302 2934 4307
rect 3713 4302 4086 4307
rect 4297 4302 4398 4307
rect 2105 4297 2278 4302
rect 4105 4297 4190 4302
rect 1945 4292 2110 4297
rect 2273 4292 2334 4297
rect 2345 4292 2598 4297
rect 2593 4287 2598 4292
rect 2681 4292 2846 4297
rect 2953 4292 4110 4297
rect 4185 4292 4270 4297
rect 2681 4287 2686 4292
rect 1489 4282 1638 4287
rect 1673 4282 1734 4287
rect 1825 4282 1934 4287
rect 2073 4282 2574 4287
rect 2593 4282 2686 4287
rect 2705 4282 2758 4287
rect 3649 4282 4174 4287
rect 4377 4282 4414 4287
rect 1489 4277 1494 4282
rect 969 4272 1494 4277
rect 1633 4277 1638 4282
rect 1825 4277 1830 4282
rect 1929 4277 2078 4282
rect 1633 4272 1830 4277
rect 2201 4272 2390 4277
rect 2801 4272 3278 4277
rect 3585 4272 3614 4277
rect 3713 4272 3934 4277
rect 4089 4272 4134 4277
rect 4193 4272 4358 4277
rect 2097 4267 2206 4272
rect 2385 4267 2494 4272
rect 2801 4267 2806 4272
rect 3609 4267 3718 4272
rect 3929 4267 4094 4272
rect 4193 4267 4198 4272
rect 737 4262 950 4267
rect 1505 4262 1654 4267
rect 1945 4262 2102 4267
rect 2225 4262 2366 4267
rect 2489 4262 2806 4267
rect 3737 4262 3910 4267
rect 4113 4262 4198 4267
rect 4353 4267 4358 4272
rect 4353 4262 4430 4267
rect 737 4247 742 4262
rect 713 4242 742 4247
rect 945 4247 950 4262
rect 1737 4257 1902 4262
rect 1945 4257 1950 4262
rect 4257 4257 4334 4262
rect 1113 4252 1198 4257
rect 1473 4252 1526 4257
rect 1553 4252 1742 4257
rect 1897 4252 1950 4257
rect 2113 4252 2214 4257
rect 2329 4252 2470 4257
rect 2825 4252 2854 4257
rect 3593 4252 4262 4257
rect 4329 4252 4422 4257
rect 4449 4252 4542 4257
rect 1113 4247 1118 4252
rect 945 4242 1118 4247
rect 1193 4247 1198 4252
rect 2113 4247 2118 4252
rect 2209 4247 2334 4252
rect 4449 4247 4454 4252
rect 1193 4242 1566 4247
rect 1753 4242 2118 4247
rect 2929 4242 2998 4247
rect 1561 4237 1758 4242
rect 2929 4237 2934 4242
rect 441 4232 582 4237
rect 441 4227 446 4232
rect 129 4222 174 4227
rect 201 4222 262 4227
rect 281 4222 310 4227
rect 329 4222 374 4227
rect 417 4222 446 4227
rect 577 4227 582 4232
rect 625 4232 974 4237
rect 1129 4232 1182 4237
rect 1505 4232 1542 4237
rect 1777 4232 1886 4237
rect 2193 4232 2638 4237
rect 2857 4232 2934 4237
rect 2993 4237 2998 4242
rect 3033 4242 3430 4247
rect 3449 4242 3630 4247
rect 3865 4242 3926 4247
rect 4273 4242 4454 4247
rect 4537 4247 4542 4252
rect 4537 4242 4566 4247
rect 4585 4242 4686 4247
rect 3033 4237 3038 4242
rect 2993 4232 3038 4237
rect 3425 4237 3430 4242
rect 3649 4237 3750 4242
rect 3945 4237 4014 4242
rect 4105 4237 4222 4242
rect 4585 4237 4590 4242
rect 3425 4232 3654 4237
rect 3745 4232 3950 4237
rect 4009 4232 4110 4237
rect 4217 4232 4246 4237
rect 4361 4232 4590 4237
rect 4681 4237 4686 4242
rect 4681 4232 4710 4237
rect 625 4227 630 4232
rect 1257 4227 1326 4232
rect 2193 4227 2198 4232
rect 4241 4227 4246 4232
rect 577 4222 630 4227
rect 905 4222 950 4227
rect 1105 4222 1262 4227
rect 1321 4222 2198 4227
rect 2209 4222 2254 4227
rect 2737 4222 2782 4227
rect 681 4217 758 4222
rect 2841 4217 2846 4227
rect 3105 4222 3262 4227
rect 3361 4222 3390 4227
rect 3481 4222 3518 4227
rect 3617 4222 3646 4227
rect 3657 4222 3734 4227
rect 3833 4222 3862 4227
rect 3913 4222 3998 4227
rect 4121 4222 4222 4227
rect 4241 4222 4270 4227
rect 4353 4222 4414 4227
rect 4409 4217 4414 4222
rect 4497 4222 4526 4227
rect 4569 4222 4646 4227
rect 4673 4222 4702 4227
rect 4497 4217 4502 4222
rect 233 4207 238 4217
rect 281 4212 326 4217
rect 425 4212 470 4217
rect 481 4212 686 4217
rect 753 4212 822 4217
rect 1033 4212 1134 4217
rect 1273 4212 1310 4217
rect 1513 4212 1550 4217
rect 1801 4212 2318 4217
rect 2665 4212 2878 4217
rect 2945 4212 2982 4217
rect 3049 4212 3350 4217
rect 3369 4212 3598 4217
rect 4041 4212 4118 4217
rect 4145 4212 4366 4217
rect 4409 4212 4502 4217
rect 1649 4207 1766 4212
rect 4673 4207 4678 4222
rect 233 4202 262 4207
rect 585 4202 622 4207
rect 697 4202 974 4207
rect 1169 4202 1214 4207
rect 1497 4202 1654 4207
rect 1761 4202 2086 4207
rect 2329 4202 3718 4207
rect 3881 4202 3926 4207
rect 4193 4202 4318 4207
rect 4585 4202 4654 4207
rect 4673 4202 4702 4207
rect 2081 4197 2334 4202
rect 4585 4197 4590 4202
rect 161 4192 286 4197
rect 361 4192 646 4197
rect 665 4192 710 4197
rect 921 4192 950 4197
rect 1097 4192 1158 4197
rect 1249 4192 1278 4197
rect 1337 4192 1526 4197
rect 1665 4192 1750 4197
rect 1857 4192 1926 4197
rect 1977 4192 2062 4197
rect 2617 4192 2846 4197
rect 2889 4192 2998 4197
rect 3113 4192 3158 4197
rect 3185 4192 3254 4197
rect 3273 4192 3334 4197
rect 3345 4192 3446 4197
rect 3473 4192 3678 4197
rect 3825 4192 3870 4197
rect 4377 4192 4454 4197
rect 4561 4192 4590 4197
rect 4649 4197 4654 4202
rect 4737 4197 4742 4217
rect 4649 4192 4766 4197
rect 729 4187 902 4192
rect 969 4187 1070 4192
rect 1153 4187 1254 4192
rect 1545 4187 1646 4192
rect 1745 4187 1750 4192
rect 2521 4187 2598 4192
rect 3329 4187 3334 4192
rect 577 4182 734 4187
rect 897 4182 974 4187
rect 1065 4182 1094 4187
rect 1401 4182 1438 4187
rect 1481 4182 1550 4187
rect 1641 4182 1678 4187
rect 1745 4182 2526 4187
rect 2593 4182 2662 4187
rect 2921 4182 3230 4187
rect 3241 4182 3310 4187
rect 3329 4182 3550 4187
rect 3865 4182 4182 4187
rect 1297 4177 1382 4182
rect 2657 4177 2774 4182
rect 2921 4177 2926 4182
rect 4177 4177 4182 4182
rect 4273 4182 4302 4187
rect 4465 4182 4670 4187
rect 4737 4182 4774 4187
rect 4273 4177 4278 4182
rect 209 4172 1302 4177
rect 1377 4172 2070 4177
rect 2537 4172 2638 4177
rect 2769 4172 2926 4177
rect 3009 4172 3070 4177
rect 3153 4172 3198 4177
rect 3569 4172 3670 4177
rect 4177 4172 4278 4177
rect 4705 4172 4734 4177
rect 281 4162 310 4167
rect 817 4162 1126 4167
rect 1313 4162 1382 4167
rect 1401 4162 1590 4167
rect 1633 4162 1662 4167
rect 601 4157 718 4162
rect 1121 4157 1318 4162
rect 1657 4157 1662 4162
rect 1745 4162 1774 4167
rect 1745 4157 1750 4162
rect 273 4152 606 4157
rect 713 4152 838 4157
rect 961 4152 1102 4157
rect 1337 4152 1366 4157
rect 1521 4152 1630 4157
rect 1657 4152 1750 4157
rect 1817 4152 1870 4157
rect 1361 4147 1526 4152
rect 401 4142 430 4147
rect 617 4142 702 4147
rect 889 4142 1022 4147
rect 1161 4142 1286 4147
rect 1545 4142 1638 4147
rect 1785 4142 1886 4147
rect 1905 4142 1910 4172
rect 3217 4167 3350 4172
rect 3465 4167 3574 4172
rect 3665 4167 3670 4172
rect 3793 4167 3918 4172
rect 1937 4162 1990 4167
rect 2225 4162 2750 4167
rect 2745 4157 2750 4162
rect 2945 4162 3222 4167
rect 3345 4162 3374 4167
rect 3441 4162 3470 4167
rect 3665 4162 3798 4167
rect 3913 4162 3942 4167
rect 3953 4162 4006 4167
rect 4081 4162 4134 4167
rect 4673 4162 4742 4167
rect 4753 4162 4782 4167
rect 2945 4157 2950 4162
rect 2041 4152 2078 4157
rect 2105 4152 2206 4157
rect 2593 4152 2622 4157
rect 2745 4152 2950 4157
rect 2969 4152 3566 4157
rect 3601 4152 3846 4157
rect 3905 4152 4014 4157
rect 4633 4152 4718 4157
rect 2105 4147 2110 4152
rect 1977 4142 2030 4147
rect 2025 4137 2030 4142
rect 2089 4142 2110 4147
rect 2201 4147 2206 4152
rect 2369 4147 2574 4152
rect 2201 4142 2374 4147
rect 2569 4142 2694 4147
rect 3033 4142 3174 4147
rect 3217 4142 3846 4147
rect 2089 4137 2094 4142
rect 2689 4137 2694 4142
rect 3841 4137 3846 4142
rect 4025 4142 4198 4147
rect 4385 4142 4462 4147
rect 4641 4142 4726 4147
rect 4025 4137 4030 4142
rect 225 4132 454 4137
rect 553 4132 614 4137
rect 689 4132 910 4137
rect 905 4127 910 4132
rect 1001 4132 1030 4137
rect 1177 4132 1222 4137
rect 1289 4132 1334 4137
rect 1393 4132 1430 4137
rect 1457 4132 1646 4137
rect 1753 4132 1798 4137
rect 2025 4132 2094 4137
rect 2121 4132 2190 4137
rect 2385 4132 2486 4137
rect 2513 4132 2566 4137
rect 2689 4132 2726 4137
rect 3169 4132 3366 4137
rect 3457 4132 3486 4137
rect 1001 4127 1006 4132
rect 2185 4127 2390 4132
rect 2969 4127 3110 4132
rect 3481 4127 3486 4132
rect 3545 4132 3702 4137
rect 3713 4132 3822 4137
rect 3841 4132 4030 4137
rect 4185 4132 4318 4137
rect 3545 4127 3550 4132
rect 169 4122 262 4127
rect 481 4122 606 4127
rect 905 4122 1006 4127
rect 2409 4122 2774 4127
rect 2897 4122 2974 4127
rect 3105 4122 3422 4127
rect 3481 4122 3550 4127
rect 4193 4122 4598 4127
rect 161 4112 206 4117
rect 369 4112 414 4117
rect 497 4112 582 4117
rect 673 4112 886 4117
rect 881 4107 886 4112
rect 1041 4112 2422 4117
rect 2473 4112 2542 4117
rect 2617 4112 2662 4117
rect 2985 4112 3094 4117
rect 3177 4112 3270 4117
rect 3569 4112 3630 4117
rect 3785 4112 3894 4117
rect 3961 4112 4014 4117
rect 4113 4112 4214 4117
rect 4273 4112 4342 4117
rect 4361 4112 4398 4117
rect 4561 4112 4750 4117
rect 1041 4107 1046 4112
rect 3321 4107 3422 4112
rect 81 4102 182 4107
rect 401 4102 662 4107
rect 881 4102 1046 4107
rect 2409 4102 2438 4107
rect 2569 4102 2622 4107
rect 2713 4102 2902 4107
rect 2937 4102 2974 4107
rect 3057 4102 3190 4107
rect 3201 4102 3326 4107
rect 3417 4102 3502 4107
rect 3585 4102 3662 4107
rect 3777 4102 3806 4107
rect 2713 4097 2718 4102
rect 233 4092 286 4097
rect 553 4092 638 4097
rect 777 4092 862 4097
rect 2513 4092 2718 4097
rect 2897 4097 2902 4102
rect 3801 4097 3806 4102
rect 3889 4102 3918 4107
rect 4065 4102 4110 4107
rect 4281 4102 4318 4107
rect 3889 4097 3894 4102
rect 4337 4097 4342 4112
rect 4529 4102 4574 4107
rect 4529 4097 4534 4102
rect 2897 4092 3118 4097
rect 3337 4092 3406 4097
rect 3489 4092 3598 4097
rect 3801 4092 3894 4097
rect 4201 4092 4238 4097
rect 4337 4092 4534 4097
rect 4553 4092 4654 4097
rect 2753 4087 2862 4092
rect 3113 4087 3342 4092
rect 1073 4082 2502 4087
rect 2497 4077 2502 4082
rect 2729 4082 2758 4087
rect 2857 4082 2886 4087
rect 241 4072 302 4077
rect 2497 4072 2574 4077
rect 2569 4067 2574 4072
rect 2729 4067 2734 4082
rect 2953 4077 3094 4082
rect 3361 4077 3646 4082
rect 2753 4072 2782 4077
rect 1033 4062 1254 4067
rect 1281 4062 1342 4067
rect 1497 4062 1550 4067
rect 1865 4062 1958 4067
rect 2025 4062 2214 4067
rect 2569 4062 2734 4067
rect 2777 4067 2782 4072
rect 2841 4072 2958 4077
rect 3089 4072 3366 4077
rect 3641 4072 3766 4077
rect 3785 4072 3926 4077
rect 2841 4067 2846 4072
rect 3785 4067 3790 4072
rect 2777 4062 2846 4067
rect 2865 4062 2894 4067
rect 2889 4057 2894 4062
rect 2969 4062 3078 4067
rect 3377 4062 3614 4067
rect 3761 4062 3790 4067
rect 3921 4067 3926 4072
rect 3921 4062 4374 4067
rect 2969 4057 2974 4062
rect 3073 4057 3382 4062
rect 3609 4057 3766 4062
rect 241 4052 1086 4057
rect 1705 4052 1838 4057
rect 2393 4052 2526 4057
rect 2889 4052 2974 4057
rect 2993 4052 3054 4057
rect 3401 4052 3590 4057
rect 4049 4052 4078 4057
rect 1865 4047 2222 4052
rect 2393 4047 2398 4052
rect 137 4042 222 4047
rect 1705 4042 1734 4047
rect 137 4037 142 4042
rect 81 4032 142 4037
rect 217 4037 222 4042
rect 993 4037 1078 4042
rect 1729 4037 1734 4042
rect 1793 4042 1870 4047
rect 2217 4042 2398 4047
rect 2521 4047 2526 4052
rect 2521 4042 2550 4047
rect 2649 4042 2846 4047
rect 1793 4037 1798 4042
rect 2649 4037 2654 4042
rect 217 4032 326 4037
rect 641 4032 758 4037
rect 969 4032 998 4037
rect 1073 4032 1134 4037
rect 1257 4032 1294 4037
rect 1313 4032 1686 4037
rect 1729 4032 1798 4037
rect 1881 4032 1910 4037
rect 641 4027 646 4032
rect 153 4022 246 4027
rect 305 4022 358 4027
rect 489 4022 566 4027
rect 617 4022 646 4027
rect 753 4017 758 4032
rect 857 4022 950 4027
rect 977 4022 1062 4027
rect 1137 4022 1190 4027
rect 857 4017 862 4022
rect 641 4012 734 4017
rect 753 4012 862 4017
rect 945 4017 950 4022
rect 1313 4017 1318 4032
rect 1681 4017 1686 4032
rect 1905 4027 1910 4032
rect 1977 4032 2654 4037
rect 2841 4037 2846 4042
rect 3161 4042 3286 4047
rect 3441 4042 3910 4047
rect 3161 4037 3166 4042
rect 2841 4032 3166 4037
rect 3281 4037 3286 4042
rect 3281 4032 3382 4037
rect 3449 4032 3646 4037
rect 3985 4032 4022 4037
rect 4313 4032 4382 4037
rect 4577 4032 4670 4037
rect 1977 4027 1982 4032
rect 1817 4022 1862 4027
rect 1905 4022 1982 4027
rect 2001 4022 2046 4027
rect 2145 4022 2270 4027
rect 2281 4022 2342 4027
rect 2665 4022 2846 4027
rect 3177 4022 3270 4027
rect 3425 4022 3478 4027
rect 3497 4022 4214 4027
rect 4225 4022 4286 4027
rect 4369 4022 4406 4027
rect 4449 4022 4518 4027
rect 4553 4022 4662 4027
rect 945 4012 1318 4017
rect 1577 4012 1662 4017
rect 1681 4012 1710 4017
rect 2081 4012 2134 4017
rect 2593 4012 2678 4017
rect 2697 4012 2814 4017
rect 3105 4012 3198 4017
rect 3385 4012 3406 4017
rect 3969 4012 4046 4017
rect 4201 4012 4254 4017
rect 4273 4012 4358 4017
rect 1577 4007 1582 4012
rect 633 4002 766 4007
rect 873 4002 958 4007
rect 1129 4002 1582 4007
rect 1657 4007 1662 4012
rect 3545 4007 3654 4012
rect 4273 4007 4278 4012
rect 4497 4007 4614 4012
rect 1657 4002 2214 4007
rect 2225 4002 2294 4007
rect 2353 4002 2414 4007
rect 2433 4002 2510 4007
rect 2577 4002 2718 4007
rect 2865 4002 3086 4007
rect 3377 4002 3550 4007
rect 3649 4002 3678 4007
rect 4193 4002 4278 4007
rect 4377 4002 4502 4007
rect 4609 4002 4638 4007
rect 2209 3997 2214 4002
rect 2433 3997 2438 4002
rect 561 3992 662 3997
rect 961 3992 1166 3997
rect 1241 3992 1294 3997
rect 1593 3992 1678 3997
rect 1793 3992 1822 3997
rect 2081 3992 2182 3997
rect 2209 3992 2318 3997
rect 2369 3992 2438 3997
rect 2505 3997 2510 4002
rect 2865 3997 2870 4002
rect 2505 3992 2870 3997
rect 3081 3997 3086 4002
rect 3081 3992 3246 3997
rect 3561 3992 3654 3997
rect 3737 3992 3926 3997
rect 4153 3992 4254 3997
rect 4513 3992 4574 3997
rect 4649 3992 4678 3997
rect 4273 3987 4494 3992
rect 617 3982 646 3987
rect 713 3982 870 3987
rect 921 3982 950 3987
rect 945 3977 950 3982
rect 1017 3982 1110 3987
rect 2177 3982 2286 3987
rect 2313 3982 2630 3987
rect 2729 3982 2758 3987
rect 3025 3982 3350 3987
rect 3369 3982 3510 3987
rect 3585 3982 3702 3987
rect 3913 3982 4278 3987
rect 4489 3982 4702 3987
rect 1017 3977 1022 3982
rect 3369 3977 3374 3982
rect 145 3972 190 3977
rect 945 3972 1022 3977
rect 1457 3972 3230 3977
rect 3345 3972 3374 3977
rect 3505 3977 3510 3982
rect 3769 3977 3878 3982
rect 3505 3972 3646 3977
rect 3713 3972 3774 3977
rect 3873 3972 3902 3977
rect 3225 3967 3350 3972
rect 3641 3967 3718 3972
rect 3897 3967 3902 3972
rect 4025 3972 4054 3977
rect 4209 3972 4526 3977
rect 4609 3972 4798 3977
rect 4025 3967 4030 3972
rect 4521 3967 4614 3972
rect 217 3962 318 3967
rect 1265 3962 1350 3967
rect 2017 3962 2046 3967
rect 2145 3962 2254 3967
rect 2273 3962 2782 3967
rect 2961 3962 3046 3967
rect 3377 3962 3414 3967
rect 3449 3962 3494 3967
rect 3577 3962 3622 3967
rect 3785 3962 3862 3967
rect 3897 3962 4030 3967
rect 4393 3962 4438 3967
rect 217 3957 222 3962
rect 193 3952 222 3957
rect 313 3957 318 3962
rect 1881 3957 1998 3962
rect 2801 3957 2942 3962
rect 3065 3957 3206 3962
rect 4633 3957 4742 3962
rect 313 3952 446 3957
rect 977 3952 1014 3957
rect 1025 3952 1046 3957
rect 1089 3952 1214 3957
rect 1801 3952 1886 3957
rect 1993 3952 2038 3957
rect 2161 3952 2238 3957
rect 2321 3952 2382 3957
rect 2609 3952 2806 3957
rect 2937 3952 3070 3957
rect 3201 3952 3774 3957
rect 4049 3952 4382 3957
rect 4449 3952 4478 3957
rect 4553 3952 4638 3957
rect 4737 3952 4766 3957
rect 1089 3947 1094 3952
rect 177 3942 214 3947
rect 441 3942 518 3947
rect 993 3942 1094 3947
rect 1209 3947 1214 3952
rect 2401 3947 2590 3952
rect 3769 3947 3774 3952
rect 4377 3947 4454 3952
rect 1209 3942 1238 3947
rect 1465 3942 1654 3947
rect 1897 3942 1918 3947
rect 1969 3942 2030 3947
rect 2057 3942 2118 3947
rect 2225 3942 2406 3947
rect 2585 3942 2966 3947
rect 3009 3942 3142 3947
rect 161 3932 310 3937
rect 809 3932 854 3937
rect 1385 3932 1446 3937
rect 1465 3927 1470 3942
rect 145 3922 182 3927
rect 497 3922 590 3927
rect 633 3922 766 3927
rect 1105 3922 1222 3927
rect 1233 3922 1470 3927
rect 1649 3927 1654 3942
rect 3185 3937 3190 3947
rect 3385 3942 3494 3947
rect 3593 3942 3654 3947
rect 3665 3942 3750 3947
rect 3769 3942 4022 3947
rect 4225 3942 4278 3947
rect 4537 3942 4566 3947
rect 4649 3942 4726 3947
rect 3665 3937 3670 3942
rect 1713 3927 1718 3937
rect 1801 3932 1878 3937
rect 1929 3932 2886 3937
rect 3041 3932 3206 3937
rect 1801 3927 1806 3932
rect 1649 3922 1718 3927
rect 1745 3922 1806 3927
rect 1873 3927 1878 3932
rect 3041 3927 3046 3932
rect 1873 3922 2742 3927
rect 2873 3922 2926 3927
rect 3017 3922 3046 3927
rect 3201 3927 3206 3932
rect 3473 3932 3670 3937
rect 4361 3932 4494 3937
rect 4617 3932 4646 3937
rect 3473 3927 3478 3932
rect 4161 3927 4270 3932
rect 3201 3922 3478 3927
rect 3697 3922 3862 3927
rect 1233 3917 1238 3922
rect 1745 3917 1750 3922
rect 2737 3917 2878 3922
rect 2921 3917 3022 3922
rect 3857 3917 3862 3922
rect 4033 3922 4166 3927
rect 4265 3922 4518 3927
rect 4033 3917 4038 3922
rect 129 3912 174 3917
rect 409 3912 454 3917
rect 617 3912 662 3917
rect 737 3912 790 3917
rect 905 3912 950 3917
rect 969 3912 1086 3917
rect 969 3907 974 3912
rect 289 3902 398 3907
rect 393 3897 398 3902
rect 465 3902 526 3907
rect 609 3902 726 3907
rect 801 3902 974 3907
rect 1081 3907 1086 3912
rect 1137 3912 1238 3917
rect 1321 3912 1350 3917
rect 1137 3907 1142 3912
rect 1345 3907 1350 3912
rect 1481 3912 1638 3917
rect 1697 3912 1750 3917
rect 1817 3912 1886 3917
rect 2089 3912 2158 3917
rect 2273 3912 2294 3917
rect 2305 3912 2382 3917
rect 2497 3912 2566 3917
rect 2593 3912 2718 3917
rect 3065 3912 3134 3917
rect 3857 3912 4038 3917
rect 4177 3912 4254 3917
rect 4353 3912 4422 3917
rect 1481 3907 1486 3912
rect 1977 3907 2070 3912
rect 1081 3902 1142 3907
rect 1153 3902 1238 3907
rect 1345 3902 1486 3907
rect 1785 3902 1814 3907
rect 1897 3902 1982 3907
rect 2065 3902 2286 3907
rect 465 3897 470 3902
rect 609 3897 614 3902
rect 721 3897 806 3902
rect 1809 3897 1902 3902
rect 393 3892 470 3897
rect 489 3892 614 3897
rect 1993 3892 2182 3897
rect 2281 3887 2286 3902
rect 2513 3902 2662 3907
rect 2513 3887 2518 3902
rect 2657 3897 2662 3902
rect 2769 3902 2998 3907
rect 2769 3897 2774 3902
rect 2537 3892 2638 3897
rect 2657 3892 2774 3897
rect 2793 3892 2822 3897
rect 609 3882 1990 3887
rect 2105 3882 2190 3887
rect 2281 3882 2518 3887
rect 2817 3887 2822 3892
rect 2897 3892 2926 3897
rect 4257 3892 4278 3897
rect 2897 3887 2902 3892
rect 2817 3882 2902 3887
rect 3601 3882 3662 3887
rect 3841 3882 3926 3887
rect 4177 3882 4270 3887
rect 2201 3872 2262 3877
rect 865 3862 958 3867
rect 1009 3862 1294 3867
rect 1377 3862 1422 3867
rect 1809 3862 1838 3867
rect 1921 3862 1942 3867
rect 2569 3862 2710 3867
rect 865 3857 870 3862
rect 569 3852 870 3857
rect 953 3857 958 3862
rect 2265 3857 2342 3862
rect 953 3852 998 3857
rect 1305 3852 1366 3857
rect 1433 3852 1934 3857
rect 2033 3852 2270 3857
rect 2337 3852 2550 3857
rect 993 3847 998 3852
rect 1145 3847 1310 3852
rect 1361 3847 1438 3852
rect 2569 3847 2574 3862
rect 2705 3847 2710 3862
rect 3129 3862 3214 3867
rect 3761 3862 3846 3867
rect 3129 3857 3134 3862
rect 2825 3852 2878 3857
rect 3009 3852 3134 3857
rect 3209 3857 3214 3862
rect 3209 3852 3238 3857
rect 3881 3852 4014 3857
rect 4033 3852 4054 3857
rect 4217 3852 4334 3857
rect 3881 3847 3886 3852
rect 881 3842 942 3847
rect 993 3842 1150 3847
rect 2281 3842 2326 3847
rect 2521 3842 2574 3847
rect 2593 3842 2670 3847
rect 2705 3842 2734 3847
rect 2993 3842 3286 3847
rect 3473 3842 3542 3847
rect 3857 3842 3886 3847
rect 4009 3847 4014 3852
rect 4009 3842 4238 3847
rect 2345 3837 2502 3842
rect 2593 3837 2598 3842
rect 265 3832 326 3837
rect 481 3832 638 3837
rect 657 3832 790 3837
rect 809 3832 838 3837
rect 881 3832 926 3837
rect 945 3832 966 3837
rect 1169 3832 1198 3837
rect 657 3827 662 3832
rect 249 3822 310 3827
rect 385 3822 430 3827
rect 441 3822 494 3827
rect 577 3822 662 3827
rect 785 3827 790 3832
rect 1193 3827 1198 3832
rect 1281 3832 1774 3837
rect 1281 3827 1286 3832
rect 1769 3827 1774 3832
rect 1881 3832 2350 3837
rect 2497 3832 2598 3837
rect 2665 3837 2670 3842
rect 2897 3837 2974 3842
rect 2665 3832 2694 3837
rect 2801 3832 2902 3837
rect 2969 3832 3198 3837
rect 3297 3832 4038 3837
rect 4249 3832 4334 3837
rect 1881 3827 1886 3832
rect 2689 3827 2790 3832
rect 3193 3827 3302 3832
rect 4033 3827 4254 3832
rect 785 3822 974 3827
rect 1081 3822 1118 3827
rect 1193 3822 1286 3827
rect 1721 3822 1750 3827
rect 1769 3822 1886 3827
rect 2289 3822 2502 3827
rect 2609 3822 2654 3827
rect 2785 3822 2846 3827
rect 2913 3822 3022 3827
rect 3041 3822 3174 3827
rect 3457 3822 3486 3827
rect 3945 3822 4014 3827
rect 4273 3822 4342 3827
rect 4497 3822 4590 3827
rect 4497 3817 4502 3822
rect 201 3812 246 3817
rect 273 3812 302 3817
rect 313 3812 374 3817
rect 505 3812 926 3817
rect 953 3812 1038 3817
rect 1305 3812 1502 3817
rect 1569 3812 1646 3817
rect 241 3797 246 3812
rect 369 3807 510 3812
rect 1569 3807 1574 3812
rect 633 3802 870 3807
rect 1089 3802 1150 3807
rect 1441 3802 1574 3807
rect 1641 3807 1646 3812
rect 1905 3812 2006 3817
rect 2313 3812 2334 3817
rect 2457 3812 2510 3817
rect 2545 3812 2702 3817
rect 2785 3812 2926 3817
rect 3001 3812 3070 3817
rect 3193 3812 3286 3817
rect 1641 3802 1702 3807
rect 865 3797 966 3802
rect 1905 3797 1910 3812
rect 3193 3807 3198 3812
rect 1929 3802 2054 3807
rect 2065 3802 2446 3807
rect 2441 3797 2446 3802
rect 2601 3802 3198 3807
rect 3281 3807 3286 3812
rect 3825 3812 3926 3817
rect 4073 3812 4286 3817
rect 4473 3812 4502 3817
rect 4585 3817 4590 3822
rect 4585 3812 4614 3817
rect 3825 3807 3830 3812
rect 3921 3807 4054 3812
rect 3281 3802 3830 3807
rect 4049 3802 4142 3807
rect 4553 3802 4598 3807
rect 2601 3797 2606 3802
rect 185 3792 222 3797
rect 241 3792 406 3797
rect 417 3792 510 3797
rect 641 3792 678 3797
rect 785 3792 846 3797
rect 961 3792 1070 3797
rect 1169 3792 1198 3797
rect 1233 3792 1342 3797
rect 1361 3792 1518 3797
rect 1585 3792 1630 3797
rect 1777 3792 1910 3797
rect 1993 3792 2038 3797
rect 2441 3792 2606 3797
rect 2625 3792 2662 3797
rect 2705 3792 2814 3797
rect 2881 3792 2958 3797
rect 3025 3792 3110 3797
rect 3201 3792 3270 3797
rect 3377 3792 3406 3797
rect 3841 3792 3902 3797
rect 3913 3792 3966 3797
rect 3985 3792 4078 3797
rect 4513 3792 4598 3797
rect 4641 3792 4726 3797
rect 401 3787 406 3792
rect 545 3787 622 3792
rect 689 3787 790 3792
rect 1065 3787 1150 3792
rect 1233 3787 1238 3792
rect 401 3782 550 3787
rect 617 3782 694 3787
rect 809 3782 950 3787
rect 1145 3782 1238 3787
rect 1337 3787 1342 3792
rect 1337 3782 1798 3787
rect 1985 3782 2126 3787
rect 2169 3782 2198 3787
rect 2265 3782 2318 3787
rect 2753 3782 2790 3787
rect 2905 3782 2974 3787
rect 3361 3782 3470 3787
rect 3817 3782 3854 3787
rect 3889 3782 3918 3787
rect 313 3777 382 3782
rect 945 3777 950 3782
rect 3913 3777 3918 3782
rect 4089 3782 4182 3787
rect 4089 3777 4094 3782
rect 257 3772 318 3777
rect 377 3772 470 3777
rect 561 3772 926 3777
rect 945 3772 1438 3777
rect 1609 3772 1638 3777
rect 1769 3772 1830 3777
rect 2001 3772 2030 3777
rect 2057 3772 2078 3777
rect 2337 3772 2606 3777
rect 2945 3772 3190 3777
rect 465 3767 566 3772
rect 1433 3767 1534 3772
rect 1609 3767 1614 3772
rect 2337 3767 2342 3772
rect 145 3762 238 3767
rect 329 3762 446 3767
rect 585 3762 766 3767
rect 145 3757 150 3762
rect 89 3752 150 3757
rect 233 3757 238 3762
rect 761 3757 766 3762
rect 849 3762 1006 3767
rect 1049 3762 1222 3767
rect 1529 3762 1614 3767
rect 1889 3762 1998 3767
rect 2017 3762 2342 3767
rect 2601 3767 2606 3772
rect 3185 3767 3190 3772
rect 3281 3772 3374 3777
rect 3673 3772 3742 3777
rect 3761 3772 3790 3777
rect 3913 3772 4094 3777
rect 4529 3772 4582 3777
rect 3281 3767 3286 3772
rect 3673 3767 3678 3772
rect 2601 3762 2750 3767
rect 3185 3762 3286 3767
rect 3465 3762 3678 3767
rect 3737 3767 3742 3772
rect 3737 3762 3870 3767
rect 4417 3762 4502 3767
rect 4577 3762 4790 3767
rect 849 3757 854 3762
rect 233 3752 310 3757
rect 337 3752 518 3757
rect 585 3752 654 3757
rect 665 3752 742 3757
rect 761 3752 854 3757
rect 873 3752 974 3757
rect 1097 3752 1350 3757
rect 1457 3752 1510 3757
rect 1793 3752 2022 3757
rect 2033 3752 2070 3757
rect 3649 3752 3718 3757
rect 4113 3752 4190 3757
rect 4345 3752 4566 3757
rect 2529 3747 2622 3752
rect 4113 3747 4118 3752
rect 169 3742 214 3747
rect 385 3742 470 3747
rect 961 3742 1006 3747
rect 1225 3742 1334 3747
rect 1481 3742 1566 3747
rect 1585 3742 1678 3747
rect 1697 3742 2086 3747
rect 2097 3742 2158 3747
rect 2177 3742 2254 3747
rect 2305 3742 2534 3747
rect 2617 3742 2806 3747
rect 2841 3742 2870 3747
rect 2889 3742 3126 3747
rect 3449 3742 3478 3747
rect 3617 3742 4118 3747
rect 4185 3747 4190 3752
rect 4185 3742 4374 3747
rect 4521 3742 4550 3747
rect 4625 3742 4646 3747
rect 1353 3737 1462 3742
rect 1585 3737 1590 3742
rect 161 3732 494 3737
rect 841 3732 950 3737
rect 1017 3732 1358 3737
rect 1457 3732 1590 3737
rect 1673 3737 1678 3742
rect 2097 3737 2102 3742
rect 1673 3732 1702 3737
rect 1929 3732 2102 3737
rect 2129 3737 2134 3742
rect 2801 3737 2806 3742
rect 2129 3732 2190 3737
rect 2353 3732 2406 3737
rect 2545 3732 2606 3737
rect 2801 3732 2830 3737
rect 945 3727 1022 3732
rect 1697 3727 1934 3732
rect 2209 3727 2334 3732
rect 2889 3727 2894 3742
rect 3121 3727 3126 3742
rect 3617 3737 3622 3742
rect 4369 3737 4526 3742
rect 3385 3732 3622 3737
rect 3633 3732 3670 3737
rect 4129 3732 4174 3737
rect 3801 3727 3886 3732
rect 193 3722 222 3727
rect 217 3717 222 3722
rect 329 3722 646 3727
rect 657 3722 678 3727
rect 777 3722 822 3727
rect 1249 3722 1286 3727
rect 1321 3722 1550 3727
rect 2081 3722 2214 3727
rect 2329 3722 2894 3727
rect 2913 3722 2990 3727
rect 3121 3722 3150 3727
rect 3409 3722 3806 3727
rect 3881 3722 3910 3727
rect 329 3717 334 3722
rect 1953 3717 2086 3722
rect 2913 3717 2918 3722
rect 89 3712 190 3717
rect 217 3712 334 3717
rect 353 3712 398 3717
rect 489 3712 518 3717
rect 513 3707 518 3712
rect 641 3712 670 3717
rect 681 3712 798 3717
rect 881 3712 1166 3717
rect 1313 3712 1390 3717
rect 1425 3712 1454 3717
rect 641 3707 646 3712
rect 1449 3707 1454 3712
rect 1513 3712 1622 3717
rect 1665 3712 1958 3717
rect 2169 3712 2198 3717
rect 2233 3712 2358 3717
rect 2569 3712 2598 3717
rect 2641 3712 2686 3717
rect 2841 3712 2918 3717
rect 2985 3717 2990 3722
rect 4169 3717 4174 3732
rect 4321 3732 4350 3737
rect 4321 3717 4326 3732
rect 4441 3722 4478 3727
rect 4665 3722 4742 3727
rect 2985 3712 3286 3717
rect 3417 3712 3630 3717
rect 3641 3712 3718 3717
rect 3817 3712 3894 3717
rect 3969 3712 3998 3717
rect 4169 3712 4326 3717
rect 4481 3712 4542 3717
rect 4665 3712 4718 3717
rect 1513 3707 1518 3712
rect 513 3702 646 3707
rect 833 3702 894 3707
rect 1281 3702 1350 3707
rect 1449 3702 1518 3707
rect 1537 3702 1638 3707
rect 1969 3702 1998 3707
rect 2017 3702 2302 3707
rect 2369 3702 2470 3707
rect 2577 3702 2606 3707
rect 2713 3702 2782 3707
rect 2873 3702 2974 3707
rect 2297 3697 2374 3702
rect 2601 3697 2718 3702
rect 1033 3692 1262 3697
rect 1657 3692 1862 3697
rect 1881 3692 2190 3697
rect 2249 3692 2278 3697
rect 1657 3687 1662 3692
rect 1281 3682 1454 3687
rect 1473 3682 1502 3687
rect 1617 3682 1662 3687
rect 1857 3687 1862 3692
rect 2273 3687 2278 3692
rect 2425 3692 2454 3697
rect 2841 3692 2870 3697
rect 2425 3687 2430 3692
rect 2969 3687 2974 3702
rect 3297 3702 3406 3707
rect 3905 3702 4094 3707
rect 4513 3702 4622 3707
rect 3297 3687 3302 3702
rect 1857 3682 1902 3687
rect 2097 3682 2142 3687
rect 2273 3682 2430 3687
rect 2569 3682 2790 3687
rect 1169 3677 1286 3682
rect 1449 3677 1454 3682
rect 1921 3677 2046 3682
rect 2785 3677 2790 3682
rect 2921 3682 2950 3687
rect 2969 3682 3302 3687
rect 3401 3687 3406 3702
rect 3841 3697 3910 3702
rect 3841 3687 3846 3697
rect 3401 3682 3846 3687
rect 3865 3682 3990 3687
rect 4545 3682 4606 3687
rect 4625 3682 4646 3687
rect 2921 3677 2926 3682
rect 961 3672 1174 3677
rect 1449 3672 1926 3677
rect 2041 3672 2070 3677
rect 2081 3672 2222 3677
rect 2785 3672 2926 3677
rect 505 3662 590 3667
rect 505 3657 510 3662
rect 481 3652 510 3657
rect 585 3657 590 3662
rect 657 3662 942 3667
rect 1185 3662 1622 3667
rect 1809 3662 2166 3667
rect 657 3657 662 3662
rect 585 3652 614 3657
rect 633 3652 662 3657
rect 937 3657 942 3662
rect 1001 3657 1142 3662
rect 1185 3657 1190 3662
rect 1705 3657 1790 3662
rect 937 3652 1006 3657
rect 1137 3652 1190 3657
rect 1201 3652 1230 3657
rect 1329 3652 1358 3657
rect 1601 3652 1710 3657
rect 1785 3652 2030 3657
rect 2073 3652 2110 3657
rect 2129 3652 2382 3657
rect 2441 3652 2766 3657
rect 3897 3652 4190 3657
rect 4209 3652 4310 3657
rect 1225 3647 1334 3652
rect 1481 3647 1582 3652
rect 2129 3647 2134 3652
rect 2441 3647 2446 3652
rect 385 3642 462 3647
rect 1017 3642 1198 3647
rect 1457 3642 1486 3647
rect 1577 3642 1638 3647
rect 1721 3642 1798 3647
rect 1841 3642 1878 3647
rect 1977 3642 2062 3647
rect 2073 3642 2134 3647
rect 2185 3642 2342 3647
rect 2417 3642 2446 3647
rect 2761 3647 2766 3652
rect 4209 3647 4214 3652
rect 2761 3642 2790 3647
rect 3369 3642 3550 3647
rect 4097 3642 4214 3647
rect 4305 3647 4310 3652
rect 4345 3652 4438 3657
rect 4345 3647 4350 3652
rect 4305 3642 4350 3647
rect 4433 3647 4438 3652
rect 4433 3642 4590 3647
rect 385 3637 390 3642
rect 233 3632 390 3637
rect 457 3637 462 3642
rect 2465 3637 2638 3642
rect 3369 3637 3374 3642
rect 457 3632 966 3637
rect 977 3632 1014 3637
rect 1089 3632 1566 3637
rect 1649 3632 1710 3637
rect 1777 3632 1990 3637
rect 2113 3632 2470 3637
rect 2633 3632 2806 3637
rect 3345 3632 3374 3637
rect 3545 3637 3550 3642
rect 3545 3632 3774 3637
rect 4561 3632 4598 3637
rect 1561 3627 1654 3632
rect 1705 3627 1782 3632
rect 921 3622 1022 3627
rect 1033 3622 1070 3627
rect 1081 3622 1206 3627
rect 1801 3622 1878 3627
rect 2425 3622 2470 3627
rect 2489 3622 2534 3627
rect 2585 3622 2622 3627
rect 1473 3617 1542 3622
rect 2225 3617 2294 3622
rect 305 3612 334 3617
rect 329 3607 334 3612
rect 401 3612 718 3617
rect 809 3612 1110 3617
rect 1145 3612 1478 3617
rect 1537 3612 2230 3617
rect 2289 3612 2422 3617
rect 2449 3612 2478 3617
rect 2513 3612 2766 3617
rect 401 3607 406 3612
rect 2801 3607 2806 3632
rect 2977 3622 3126 3627
rect 3289 3622 3374 3627
rect 3409 3622 3438 3627
rect 3873 3622 4254 3627
rect 2825 3612 2918 3617
rect 2961 3612 2998 3617
rect 3425 3612 3534 3617
rect 4289 3607 4294 3627
rect 4361 3622 4422 3627
rect 4521 3622 4614 3627
rect 4641 3622 4678 3627
rect 4345 3612 4654 3617
rect 329 3602 406 3607
rect 425 3602 454 3607
rect 449 3597 454 3602
rect 729 3602 798 3607
rect 729 3597 734 3602
rect 449 3592 734 3597
rect 793 3597 798 3602
rect 921 3602 1094 3607
rect 1489 3602 1526 3607
rect 2241 3602 2270 3607
rect 2289 3602 2390 3607
rect 2433 3602 2542 3607
rect 2801 3602 2830 3607
rect 3369 3602 3502 3607
rect 3553 3602 3598 3607
rect 3769 3602 4126 3607
rect 4289 3602 4358 3607
rect 4585 3602 4678 3607
rect 921 3597 926 3602
rect 1745 3597 1822 3602
rect 1937 3597 2006 3602
rect 2129 3597 2222 3602
rect 793 3592 926 3597
rect 945 3592 990 3597
rect 1009 3592 1078 3597
rect 1193 3592 1270 3597
rect 1345 3592 1478 3597
rect 1537 3592 1750 3597
rect 1817 3592 1942 3597
rect 2001 3592 2134 3597
rect 2217 3592 2646 3597
rect 1009 3587 1014 3592
rect 1473 3587 1542 3592
rect 2641 3587 2646 3592
rect 2841 3592 2870 3597
rect 3041 3592 3134 3597
rect 3193 3592 3462 3597
rect 3481 3592 3558 3597
rect 3761 3592 3886 3597
rect 4041 3592 4094 3597
rect 4137 3592 4174 3597
rect 4337 3592 4374 3597
rect 2841 3587 2846 3592
rect 969 3582 1014 3587
rect 1761 3582 1806 3587
rect 1953 3582 1990 3587
rect 2145 3582 2438 3587
rect 2481 3582 2502 3587
rect 2585 3582 2622 3587
rect 2641 3582 2846 3587
rect 3665 3582 3742 3587
rect 3953 3582 4070 3587
rect 4113 3582 4294 3587
rect 4489 3582 4526 3587
rect 3665 3577 3670 3582
rect 681 3572 1726 3577
rect 1777 3572 2430 3577
rect 2441 3572 2486 3577
rect 2913 3572 3022 3577
rect 3081 3572 3198 3577
rect 3641 3572 3670 3577
rect 3737 3577 3742 3582
rect 3809 3577 3878 3582
rect 3737 3572 3814 3577
rect 3873 3572 3942 3577
rect 4041 3572 4086 3577
rect 4137 3572 4198 3577
rect 4489 3572 4558 3577
rect 2913 3567 2918 3572
rect 209 3562 246 3567
rect 457 3562 638 3567
rect 1961 3562 1990 3567
rect 2153 3562 2374 3567
rect 2417 3562 2470 3567
rect 2889 3562 2918 3567
rect 3017 3567 3022 3572
rect 3937 3567 4046 3572
rect 4217 3567 4326 3572
rect 3017 3562 3254 3567
rect 3433 3562 3526 3567
rect 3545 3562 3574 3567
rect 3825 3562 3862 3567
rect 4065 3562 4222 3567
rect 4321 3562 4382 3567
rect 209 3527 214 3562
rect 657 3557 726 3562
rect 849 3557 1038 3562
rect 1289 3557 1566 3562
rect 1609 3557 1678 3562
rect 1873 3557 1942 3562
rect 2009 3557 2134 3562
rect 3433 3557 3438 3562
rect 241 3552 342 3557
rect 633 3552 662 3557
rect 721 3552 854 3557
rect 1033 3552 1294 3557
rect 1561 3552 1614 3557
rect 1673 3552 1878 3557
rect 1937 3552 2014 3557
rect 2129 3552 2414 3557
rect 2449 3552 2510 3557
rect 2665 3552 2758 3557
rect 2905 3552 3158 3557
rect 3321 3552 3390 3557
rect 3409 3552 3438 3557
rect 3521 3557 3526 3562
rect 3521 3552 3782 3557
rect 3817 3552 3998 3557
rect 4089 3552 4398 3557
rect 4497 3552 4534 3557
rect 3321 3547 3326 3552
rect 225 3542 414 3547
rect 489 3542 526 3547
rect 601 3542 710 3547
rect 865 3542 934 3547
rect 993 3542 1022 3547
rect 1305 3542 1414 3547
rect 1425 3542 1550 3547
rect 1625 3542 1662 3547
rect 1889 3542 1974 3547
rect 2025 3542 2214 3547
rect 2433 3542 2574 3547
rect 2601 3542 2678 3547
rect 2689 3542 2710 3547
rect 3025 3542 3054 3547
rect 3169 3542 3326 3547
rect 3385 3547 3390 3552
rect 3385 3542 3822 3547
rect 3833 3542 3926 3547
rect 4161 3542 4206 3547
rect 4329 3542 4430 3547
rect 4513 3542 4598 3547
rect 1409 3537 1414 3542
rect 2305 3537 2374 3542
rect 2849 3537 2934 3542
rect 3025 3537 3030 3542
rect 3049 3537 3174 3542
rect 265 3532 334 3537
rect 785 3532 1214 3537
rect 1369 3532 1398 3537
rect 1409 3532 1670 3537
rect 1921 3532 2310 3537
rect 2369 3532 2550 3537
rect 2721 3532 2854 3537
rect 2929 3532 3030 3537
rect 3465 3532 3542 3537
rect 3777 3532 3870 3537
rect 209 3522 230 3527
rect 313 3522 414 3527
rect 737 3522 774 3527
rect 769 3517 774 3522
rect 897 3522 926 3527
rect 961 3522 990 3527
rect 897 3517 902 3522
rect 185 3512 214 3517
rect 209 3507 214 3512
rect 313 3512 342 3517
rect 465 3512 494 3517
rect 769 3512 902 3517
rect 985 3517 990 3522
rect 1225 3522 1318 3527
rect 1329 3522 1382 3527
rect 1225 3517 1230 3522
rect 1393 3517 1398 3532
rect 1665 3527 1670 3532
rect 2545 3527 2726 3532
rect 3865 3527 3870 3532
rect 3969 3532 3998 3537
rect 4049 3532 4118 3537
rect 4337 3532 4406 3537
rect 3969 3527 3974 3532
rect 1513 3522 1646 3527
rect 1665 3522 1750 3527
rect 1777 3522 1806 3527
rect 1817 3522 1846 3527
rect 1969 3522 2022 3527
rect 2121 3522 2254 3527
rect 2321 3522 2358 3527
rect 2457 3522 2526 3527
rect 2865 3522 2918 3527
rect 2993 3522 3078 3527
rect 3153 3522 3198 3527
rect 3337 3522 3622 3527
rect 3865 3522 3974 3527
rect 2017 3517 2126 3522
rect 2353 3517 2358 3522
rect 985 3512 1230 3517
rect 1369 3512 1398 3517
rect 2289 3512 2342 3517
rect 2353 3512 2390 3517
rect 2449 3512 2518 3517
rect 2545 3512 2710 3517
rect 2969 3512 3086 3517
rect 3185 3512 3214 3517
rect 3257 3512 3350 3517
rect 3513 3512 3606 3517
rect 3617 3512 3622 3522
rect 4025 3512 4054 3517
rect 313 3507 318 3512
rect 1713 3507 1798 3512
rect 209 3502 318 3507
rect 385 3502 414 3507
rect 409 3497 414 3502
rect 489 3502 518 3507
rect 1281 3502 1318 3507
rect 1441 3502 1542 3507
rect 1609 3502 1718 3507
rect 1793 3502 1926 3507
rect 1937 3502 1990 3507
rect 2057 3502 2102 3507
rect 2225 3502 2246 3507
rect 2329 3502 2366 3507
rect 489 3497 494 3502
rect 2385 3497 2390 3512
rect 4049 3507 4054 3512
rect 4129 3512 4294 3517
rect 4681 3512 4726 3517
rect 4129 3507 4134 3512
rect 2401 3502 2510 3507
rect 2593 3502 2646 3507
rect 2673 3502 2710 3507
rect 3049 3502 3126 3507
rect 3321 3502 3502 3507
rect 3633 3502 3782 3507
rect 4049 3502 4134 3507
rect 4337 3502 4374 3507
rect 2593 3497 2598 3502
rect 3145 3497 3302 3502
rect 3497 3497 3638 3502
rect 409 3492 494 3497
rect 793 3492 1270 3497
rect 1553 3492 1598 3497
rect 1729 3492 1782 3497
rect 1929 3492 1958 3497
rect 2273 3492 2326 3497
rect 2385 3492 2598 3497
rect 2729 3492 2950 3497
rect 2985 3492 3150 3497
rect 3297 3492 3350 3497
rect 1265 3487 1366 3492
rect 1473 3487 1558 3492
rect 1593 3487 1734 3492
rect 2617 3487 2734 3492
rect 2945 3487 2950 3492
rect 3369 3487 3478 3492
rect 1361 3482 1478 3487
rect 2281 3482 2358 3487
rect 2409 3482 2622 3487
rect 2945 3482 2974 3487
rect 3001 3482 3374 3487
rect 3473 3482 3566 3487
rect 1033 3472 1062 3477
rect 1105 3472 1342 3477
rect 1497 3472 1534 3477
rect 1601 3472 1814 3477
rect 1977 3472 2254 3477
rect 2417 3472 2982 3477
rect 2993 3472 3294 3477
rect 3377 3472 3462 3477
rect 1977 3467 1982 3472
rect 2249 3467 2398 3472
rect 3289 3467 3382 3472
rect 3457 3467 3462 3472
rect 3553 3472 3630 3477
rect 3553 3467 3558 3472
rect 289 3462 326 3467
rect 1081 3462 1110 3467
rect 1617 3462 1646 3467
rect 1785 3462 1982 3467
rect 2393 3462 2478 3467
rect 2873 3462 2974 3467
rect 3057 3462 3270 3467
rect 3401 3462 3438 3467
rect 3457 3462 3558 3467
rect 1641 3457 1790 3462
rect 2001 3457 2230 3462
rect 2473 3457 2878 3462
rect 2969 3457 3062 3462
rect 473 3452 558 3457
rect 681 3452 734 3457
rect 1025 3452 1214 3457
rect 1945 3452 2006 3457
rect 2225 3452 2454 3457
rect 2897 3452 2950 3457
rect 3081 3452 3302 3457
rect 473 3447 478 3452
rect 449 3442 478 3447
rect 553 3447 558 3452
rect 1809 3447 1926 3452
rect 3321 3447 3494 3452
rect 553 3442 582 3447
rect 705 3442 798 3447
rect 1153 3442 1254 3447
rect 1361 3442 1598 3447
rect 1361 3437 1366 3442
rect 529 3432 582 3437
rect 721 3432 774 3437
rect 1057 3432 1150 3437
rect 1193 3432 1366 3437
rect 1593 3437 1598 3442
rect 1617 3442 1686 3447
rect 1705 3442 1774 3447
rect 1785 3442 1814 3447
rect 1921 3442 2406 3447
rect 2473 3442 2878 3447
rect 2969 3442 3326 3447
rect 3489 3442 3726 3447
rect 3937 3442 3974 3447
rect 4217 3442 4238 3447
rect 1617 3437 1622 3442
rect 1593 3432 1622 3437
rect 1681 3437 1686 3442
rect 2473 3437 2478 3442
rect 1681 3432 2478 3437
rect 2873 3437 2878 3442
rect 2873 3432 2974 3437
rect 3337 3432 3478 3437
rect 4065 3432 4142 3437
rect 2753 3427 2854 3432
rect 2969 3427 3342 3432
rect 3905 3427 4022 3432
rect 4065 3427 4070 3432
rect 89 3422 326 3427
rect 337 3422 382 3427
rect 473 3422 526 3427
rect 681 3422 718 3427
rect 1233 3422 1278 3427
rect 1633 3422 1758 3427
rect 1969 3422 2014 3427
rect 2113 3422 2158 3427
rect 2193 3422 2494 3427
rect 2505 3422 2558 3427
rect 2569 3422 2694 3427
rect 2729 3422 2758 3427
rect 2849 3422 2950 3427
rect 321 3417 326 3422
rect 1849 3417 1926 3422
rect 3361 3417 3366 3427
rect 3489 3422 3542 3427
rect 3777 3422 3870 3427
rect 3881 3422 3910 3427
rect 4017 3422 4070 3427
rect 4137 3427 4142 3432
rect 4137 3422 4182 3427
rect 4505 3422 4646 3427
rect 321 3412 406 3417
rect 1121 3412 1262 3417
rect 1377 3412 1854 3417
rect 1921 3412 1950 3417
rect 2697 3412 2806 3417
rect 2825 3412 3342 3417
rect 3361 3412 3518 3417
rect 3561 3412 3998 3417
rect 4241 3412 4326 3417
rect 2033 3407 2118 3412
rect 2161 3407 2230 3412
rect 2329 3407 2678 3412
rect 425 3402 454 3407
rect 465 3402 878 3407
rect 1025 3402 1070 3407
rect 1641 3402 1686 3407
rect 1697 3402 1750 3407
rect 1865 3402 2038 3407
rect 2113 3402 2166 3407
rect 2225 3402 2334 3407
rect 2673 3402 2990 3407
rect 3457 3402 3542 3407
rect 3857 3402 3934 3407
rect 3945 3402 3990 3407
rect 4041 3402 4126 3407
rect 4313 3402 4382 3407
rect 4489 3402 4670 3407
rect 1425 3397 1574 3402
rect 1745 3397 1870 3402
rect 3049 3397 3262 3402
rect 3321 3397 3438 3402
rect 3561 3397 3702 3402
rect 4145 3397 4262 3402
rect 4489 3397 4494 3402
rect 193 3392 254 3397
rect 289 3392 390 3397
rect 897 3392 1006 3397
rect 1185 3392 1238 3397
rect 1401 3392 1430 3397
rect 1569 3392 1662 3397
rect 1889 3392 1974 3397
rect 2049 3392 2102 3397
rect 2177 3392 2214 3397
rect 2345 3392 2486 3397
rect 2505 3392 2910 3397
rect 3001 3392 3054 3397
rect 3257 3392 3326 3397
rect 3433 3392 3566 3397
rect 3697 3392 4150 3397
rect 4257 3392 4334 3397
rect 4465 3392 4494 3397
rect 4665 3397 4670 3402
rect 4665 3392 4694 3397
rect 569 3387 646 3392
rect 897 3387 902 3392
rect 233 3382 262 3387
rect 401 3382 574 3387
rect 641 3382 670 3387
rect 729 3382 902 3387
rect 1001 3387 1006 3392
rect 2233 3387 2326 3392
rect 2481 3387 2486 3392
rect 2905 3387 3006 3392
rect 1001 3382 2238 3387
rect 2321 3382 2406 3387
rect 2481 3382 2750 3387
rect 2785 3382 2830 3387
rect 2841 3382 2886 3387
rect 3065 3382 3102 3387
rect 3137 3382 3246 3387
rect 3337 3382 3686 3387
rect 3889 3382 3918 3387
rect 4065 3382 4246 3387
rect 4353 3382 4710 3387
rect 257 3377 262 3382
rect 329 3377 406 3382
rect 3913 3377 4070 3382
rect 4265 3377 4358 3382
rect 257 3372 334 3377
rect 585 3372 678 3377
rect 945 3372 1038 3377
rect 1209 3372 1246 3377
rect 1425 3372 1598 3377
rect 1809 3372 1838 3377
rect 465 3367 534 3372
rect 737 3367 822 3372
rect 1057 3367 1158 3372
rect 1833 3367 1838 3372
rect 1913 3372 3006 3377
rect 3249 3372 3318 3377
rect 3377 3372 3422 3377
rect 3513 3372 3574 3377
rect 3809 3372 3838 3377
rect 4089 3372 4270 3377
rect 1913 3367 1918 3372
rect 4393 3367 4510 3372
rect 353 3362 470 3367
rect 529 3362 558 3367
rect 609 3362 662 3367
rect 713 3362 742 3367
rect 817 3362 1062 3367
rect 1153 3362 1182 3367
rect 1457 3362 1614 3367
rect 1665 3362 1694 3367
rect 1833 3362 1918 3367
rect 1969 3362 2334 3367
rect 2433 3362 2462 3367
rect 2545 3362 2598 3367
rect 2705 3362 2894 3367
rect 3273 3362 3318 3367
rect 3481 3362 3558 3367
rect 3569 3362 3654 3367
rect 3905 3362 4062 3367
rect 4193 3362 4398 3367
rect 4505 3362 4662 3367
rect 2457 3357 2550 3362
rect 369 3352 398 3357
rect 481 3352 734 3357
rect 777 3352 806 3357
rect 1057 3352 1326 3357
rect 1937 3352 1966 3357
rect 2121 3352 2358 3357
rect 2569 3352 2622 3357
rect 2673 3352 2710 3357
rect 2809 3352 2862 3357
rect 2913 3352 3110 3357
rect 3169 3352 3302 3357
rect 3337 3352 3462 3357
rect 3481 3352 3678 3357
rect 3705 3352 4054 3357
rect 4257 3352 4582 3357
rect 393 3347 486 3352
rect 801 3347 806 3352
rect 945 3347 1062 3352
rect 2913 3347 2918 3352
rect 97 3342 334 3347
rect 505 3342 662 3347
rect 801 3342 950 3347
rect 1081 3342 1174 3347
rect 1257 3342 1302 3347
rect 1345 3342 1438 3347
rect 1505 3342 1582 3347
rect 1713 3342 2918 3347
rect 3105 3347 3110 3352
rect 3337 3347 3342 3352
rect 3105 3342 3342 3347
rect 3457 3347 3462 3352
rect 3457 3342 3694 3347
rect 3841 3342 3926 3347
rect 4009 3342 4038 3347
rect 4337 3342 4478 3347
rect 4497 3342 4542 3347
rect 1345 3337 1350 3342
rect 353 3332 486 3337
rect 969 3332 1054 3337
rect 1161 3332 1206 3337
rect 1281 3332 1350 3337
rect 1433 3337 1438 3342
rect 3689 3337 3846 3342
rect 3921 3337 4014 3342
rect 1433 3332 1702 3337
rect 2129 3332 2198 3337
rect 2209 3332 2398 3337
rect 2625 3332 2654 3337
rect 2793 3332 3414 3337
rect 3465 3332 3494 3337
rect 3617 3332 3670 3337
rect 3865 3332 3902 3337
rect 353 3327 358 3332
rect 481 3327 590 3332
rect 969 3327 974 3332
rect 313 3322 358 3327
rect 585 3322 614 3327
rect 609 3317 614 3322
rect 673 3322 822 3327
rect 945 3322 974 3327
rect 1049 3327 1054 3332
rect 1697 3327 1838 3332
rect 2129 3327 2134 3332
rect 2393 3327 2398 3332
rect 2521 3327 2630 3332
rect 1049 3322 1078 3327
rect 1201 3322 1310 3327
rect 1361 3322 1478 3327
rect 1513 3322 1574 3327
rect 1833 3322 2134 3327
rect 2201 3322 2254 3327
rect 2393 3322 2526 3327
rect 2737 3322 2774 3327
rect 2889 3322 2934 3327
rect 2993 3322 3198 3327
rect 673 3317 678 3322
rect 3193 3317 3198 3322
rect 3257 3322 3286 3327
rect 3793 3322 3910 3327
rect 4033 3322 4038 3342
rect 4289 3332 4486 3337
rect 4057 3322 4270 3327
rect 4401 3322 4518 3327
rect 4545 3322 4574 3327
rect 4609 3322 4638 3327
rect 3257 3317 3262 3322
rect 4057 3317 4062 3322
rect 145 3312 198 3317
rect 217 3312 246 3317
rect 257 3312 566 3317
rect 609 3312 678 3317
rect 921 3312 966 3317
rect 1025 3312 1070 3317
rect 1449 3312 1638 3317
rect 1777 3312 1814 3317
rect 2153 3312 2366 3317
rect 2545 3312 2598 3317
rect 2753 3312 2798 3317
rect 2841 3312 2862 3317
rect 2985 3312 3078 3317
rect 3121 3312 3174 3317
rect 3193 3312 3262 3317
rect 3401 3312 3470 3317
rect 3489 3312 3670 3317
rect 3689 3312 3726 3317
rect 3769 3312 3814 3317
rect 3913 3312 4062 3317
rect 4265 3317 4270 3322
rect 4265 3312 4350 3317
rect 4489 3312 4534 3317
rect 4561 3312 4582 3317
rect 4745 3312 4790 3317
rect 3489 3307 3494 3312
rect 233 3302 382 3307
rect 377 3297 382 3302
rect 457 3302 590 3307
rect 721 3302 950 3307
rect 457 3297 462 3302
rect 945 3297 950 3302
rect 1081 3302 1590 3307
rect 1801 3302 2566 3307
rect 2745 3302 2774 3307
rect 2833 3302 2910 3307
rect 2921 3302 3006 3307
rect 3441 3302 3494 3307
rect 3665 3307 3670 3312
rect 3665 3302 3870 3307
rect 4369 3302 4446 3307
rect 4585 3302 4622 3307
rect 1081 3297 1086 3302
rect 177 3292 222 3297
rect 217 3287 222 3292
rect 329 3292 358 3297
rect 377 3292 462 3297
rect 897 3292 926 3297
rect 945 3292 1086 3297
rect 1457 3292 1654 3297
rect 2201 3292 2310 3297
rect 2617 3292 2726 3297
rect 2969 3292 3014 3297
rect 3249 3292 3366 3297
rect 3385 3292 3486 3297
rect 3545 3292 3710 3297
rect 3881 3292 4278 3297
rect 329 3287 334 3292
rect 2481 3287 2622 3292
rect 2721 3287 2910 3292
rect 3249 3287 3254 3292
rect 217 3282 334 3287
rect 2401 3282 2486 3287
rect 2905 3282 3254 3287
rect 3361 3287 3366 3292
rect 3705 3287 3886 3292
rect 3361 3282 3390 3287
rect 3545 3282 3686 3287
rect 3385 3277 3550 3282
rect 537 3272 2430 3277
rect 2441 3272 2894 3277
rect 2993 3272 3022 3277
rect 3569 3272 4198 3277
rect 2889 3267 2998 3272
rect 249 3262 326 3267
rect 249 3257 254 3262
rect 225 3252 254 3257
rect 321 3257 326 3262
rect 385 3262 518 3267
rect 2273 3262 2422 3267
rect 2841 3262 2870 3267
rect 3057 3262 3118 3267
rect 3137 3262 3246 3267
rect 3265 3262 3358 3267
rect 3481 3262 3630 3267
rect 4209 3262 4326 3267
rect 385 3257 390 3262
rect 321 3252 390 3257
rect 513 3257 518 3262
rect 2417 3257 2846 3262
rect 3137 3257 3142 3262
rect 513 3252 710 3257
rect 1049 3252 1078 3257
rect 1305 3252 1462 3257
rect 1689 3252 1798 3257
rect 1865 3252 1894 3257
rect 2177 3252 2398 3257
rect 2913 3252 3142 3257
rect 3241 3257 3246 3262
rect 3625 3257 3630 3262
rect 3777 3257 3902 3262
rect 4209 3257 4214 3262
rect 3241 3252 3294 3257
rect 3369 3252 3606 3257
rect 3625 3252 3782 3257
rect 3897 3252 4214 3257
rect 1305 3247 1310 3252
rect 209 3242 310 3247
rect 401 3242 558 3247
rect 1121 3242 1262 3247
rect 1281 3242 1310 3247
rect 1457 3247 1462 3252
rect 3289 3247 3374 3252
rect 1457 3242 1486 3247
rect 1505 3242 1670 3247
rect 1721 3242 1774 3247
rect 1785 3242 1886 3247
rect 2089 3242 2158 3247
rect 2265 3242 2478 3247
rect 2529 3242 2558 3247
rect 2657 3242 2846 3247
rect 3089 3242 3270 3247
rect 3401 3242 3430 3247
rect 3537 3242 3566 3247
rect 3801 3242 3878 3247
rect 1121 3237 1126 3242
rect 145 3232 182 3237
rect 241 3232 270 3237
rect 545 3232 606 3237
rect 865 3232 974 3237
rect 1025 3232 1086 3237
rect 1097 3232 1126 3237
rect 1257 3237 1262 3242
rect 1505 3237 1510 3242
rect 1257 3232 1510 3237
rect 1665 3237 1670 3242
rect 2089 3237 2094 3242
rect 1665 3232 1694 3237
rect 1897 3232 2094 3237
rect 2153 3237 2158 3242
rect 2657 3237 2662 3242
rect 2153 3232 2254 3237
rect 2313 3232 2510 3237
rect 2569 3232 2662 3237
rect 2841 3237 2846 3242
rect 3425 3237 3542 3242
rect 3801 3237 3806 3242
rect 2841 3232 3390 3237
rect 3705 3232 3806 3237
rect 3873 3237 3878 3242
rect 4345 3242 4438 3247
rect 4345 3237 4350 3242
rect 3873 3232 3902 3237
rect 3921 3232 4030 3237
rect 4105 3232 4350 3237
rect 4433 3237 4438 3242
rect 4433 3232 4582 3237
rect 241 3227 246 3232
rect 865 3227 870 3232
rect 161 3222 246 3227
rect 265 3222 310 3227
rect 505 3222 582 3227
rect 593 3222 870 3227
rect 969 3227 974 3232
rect 1689 3227 1902 3232
rect 2249 3227 2318 3232
rect 2505 3227 2574 3232
rect 2697 3227 2790 3232
rect 3921 3227 3926 3232
rect 969 3222 1054 3227
rect 1065 3222 1174 3227
rect 2337 3222 2398 3227
rect 2409 3222 2486 3227
rect 2673 3222 2702 3227
rect 2785 3222 2830 3227
rect 3097 3222 3142 3227
rect 3465 3222 3510 3227
rect 3817 3222 3926 3227
rect 3937 3222 4118 3227
rect 4681 3222 4742 3227
rect 3161 3217 3446 3222
rect 1 3212 214 3217
rect 569 3212 646 3217
rect 881 3212 966 3217
rect 1001 3212 1046 3217
rect 1041 3207 1046 3212
rect 1177 3212 1230 3217
rect 1257 3212 1310 3217
rect 1329 3212 1894 3217
rect 1913 3212 1934 3217
rect 2105 3212 2262 3217
rect 2385 3212 2486 3217
rect 2505 3212 2622 3217
rect 2641 3212 3166 3217
rect 3441 3212 3542 3217
rect 3777 3212 3990 3217
rect 4233 3212 4422 3217
rect 1177 3207 1182 3212
rect 129 3202 182 3207
rect 345 3202 422 3207
rect 1041 3202 1182 3207
rect 345 3197 350 3202
rect 185 3192 214 3197
rect 249 3192 294 3197
rect 321 3192 350 3197
rect 417 3197 422 3202
rect 1329 3197 1334 3212
rect 2505 3207 2510 3212
rect 1897 3202 1982 3207
rect 2089 3202 2454 3207
rect 2473 3202 2510 3207
rect 2617 3207 2622 3212
rect 2617 3202 2838 3207
rect 3049 3202 3294 3207
rect 3321 3202 3438 3207
rect 3521 3202 3590 3207
rect 3617 3202 4094 3207
rect 4217 3202 4270 3207
rect 4441 3202 4574 3207
rect 1489 3197 1638 3202
rect 1801 3197 1878 3202
rect 2449 3197 2454 3202
rect 3433 3197 3526 3202
rect 417 3192 1022 3197
rect 1017 3187 1022 3192
rect 1201 3192 1334 3197
rect 1465 3192 1494 3197
rect 1633 3192 1806 3197
rect 1873 3192 2438 3197
rect 2449 3192 2558 3197
rect 2577 3192 2926 3197
rect 3121 3192 3206 3197
rect 3257 3192 3326 3197
rect 1201 3187 1206 3192
rect 3321 3187 3326 3192
rect 3545 3192 3574 3197
rect 3545 3187 3550 3192
rect 145 3182 326 3187
rect 1017 3182 1206 3187
rect 1417 3182 1558 3187
rect 1577 3182 1622 3187
rect 1689 3182 1710 3187
rect 1817 3182 1918 3187
rect 1929 3182 2110 3187
rect 2497 3182 2862 3187
rect 3073 3182 3158 3187
rect 321 3177 326 3182
rect 689 3177 798 3182
rect 865 3177 942 3182
rect 1329 3177 1398 3182
rect 2177 3177 2502 3182
rect 3153 3177 3158 3182
rect 3217 3182 3278 3187
rect 3321 3182 3550 3187
rect 3585 3187 3590 3202
rect 4441 3197 4446 3202
rect 3801 3192 3830 3197
rect 3889 3192 4014 3197
rect 4041 3192 4118 3197
rect 4225 3192 4278 3197
rect 4297 3192 4446 3197
rect 3801 3187 3806 3192
rect 3585 3182 3806 3187
rect 3825 3187 3830 3192
rect 4297 3187 4302 3192
rect 3825 3182 3950 3187
rect 3985 3182 4230 3187
rect 4273 3182 4302 3187
rect 4569 3187 4574 3202
rect 4633 3192 4702 3197
rect 4569 3182 4598 3187
rect 3217 3177 3222 3182
rect 113 3172 150 3177
rect 233 3172 302 3177
rect 321 3172 406 3177
rect 665 3172 694 3177
rect 793 3172 870 3177
rect 937 3172 998 3177
rect 1225 3172 1334 3177
rect 1393 3172 2182 3177
rect 2513 3172 2662 3177
rect 2881 3172 2974 3177
rect 3153 3172 3222 3177
rect 3921 3172 4054 3177
rect 4129 3172 4206 3177
rect 4241 3172 4694 3177
rect 2697 3167 2766 3172
rect 2817 3167 2886 3172
rect 2969 3167 2974 3172
rect 425 3162 574 3167
rect 721 3162 782 3167
rect 881 3162 926 3167
rect 1233 3162 1278 3167
rect 1345 3162 1438 3167
rect 1529 3162 1734 3167
rect 1849 3162 1950 3167
rect 2185 3162 2702 3167
rect 2761 3162 2822 3167
rect 2969 3162 3086 3167
rect 3241 3162 3302 3167
rect 3433 3162 3502 3167
rect 3521 3162 3566 3167
rect 3585 3162 3758 3167
rect 3849 3162 3902 3167
rect 3937 3162 3982 3167
rect 4081 3162 4110 3167
rect 4209 3162 4310 3167
rect 4465 3162 4494 3167
rect 425 3157 430 3162
rect 281 3152 334 3157
rect 345 3152 430 3157
rect 569 3157 574 3162
rect 1729 3157 1854 3162
rect 1945 3157 2190 3162
rect 3433 3157 3438 3162
rect 569 3152 598 3157
rect 641 3152 678 3157
rect 769 3152 870 3157
rect 865 3147 870 3152
rect 937 3152 1094 3157
rect 1313 3152 1454 3157
rect 1545 3152 1710 3157
rect 1873 3152 1926 3157
rect 2209 3152 2238 3157
rect 2425 3152 2462 3157
rect 2713 3152 2750 3157
rect 2833 3152 2966 3157
rect 3137 3152 3230 3157
rect 3281 3152 3310 3157
rect 3409 3152 3438 3157
rect 3497 3157 3502 3162
rect 3585 3157 3590 3162
rect 3497 3152 3590 3157
rect 3753 3157 3758 3162
rect 3977 3157 4086 3162
rect 3753 3152 3782 3157
rect 3817 3152 3886 3157
rect 3905 3152 3958 3157
rect 4113 3152 4214 3157
rect 4257 3152 4286 3157
rect 4377 3152 4758 3157
rect 937 3147 942 3152
rect 2257 3147 2406 3152
rect 2481 3147 2606 3152
rect 2985 3147 3118 3152
rect 161 3142 262 3147
rect 337 3142 438 3147
rect 465 3142 558 3147
rect 129 3132 174 3137
rect 465 3127 470 3142
rect 553 3137 558 3142
rect 625 3142 686 3147
rect 777 3142 814 3147
rect 865 3142 942 3147
rect 1233 3142 1326 3147
rect 1425 3142 1558 3147
rect 1577 3142 1654 3147
rect 1785 3142 1934 3147
rect 1953 3142 2110 3147
rect 2129 3142 2262 3147
rect 2401 3142 2486 3147
rect 2601 3142 2830 3147
rect 2881 3142 2990 3147
rect 3113 3142 3686 3147
rect 3929 3142 4038 3147
rect 4057 3142 4118 3147
rect 4153 3142 4262 3147
rect 4273 3142 4390 3147
rect 4401 3142 4494 3147
rect 4617 3142 4710 3147
rect 625 3137 630 3142
rect 1953 3137 1958 3142
rect 553 3132 630 3137
rect 1017 3132 1038 3137
rect 1105 3132 1230 3137
rect 1281 3132 1366 3137
rect 1537 3132 1566 3137
rect 1561 3127 1566 3132
rect 1665 3132 1958 3137
rect 2105 3137 2110 3142
rect 3721 3137 3910 3142
rect 4273 3137 4278 3142
rect 2105 3132 2590 3137
rect 2673 3132 3726 3137
rect 3905 3132 4278 3137
rect 1665 3127 1670 3132
rect 1977 3127 2046 3132
rect 2585 3127 2678 3132
rect 4297 3127 4582 3132
rect 217 3122 342 3127
rect 369 3122 470 3127
rect 649 3122 742 3127
rect 649 3117 654 3122
rect 249 3112 310 3117
rect 401 3112 510 3117
rect 569 3112 598 3117
rect 609 3112 654 3117
rect 737 3117 742 3122
rect 833 3122 902 3127
rect 1561 3122 1670 3127
rect 1777 3122 1982 3127
rect 2041 3122 2134 3127
rect 2233 3122 2342 3127
rect 2433 3122 2566 3127
rect 2697 3122 2790 3127
rect 2857 3122 3310 3127
rect 833 3117 838 3122
rect 737 3112 838 3117
rect 897 3117 902 3122
rect 2433 3117 2438 3122
rect 2561 3117 2566 3122
rect 3305 3117 3310 3122
rect 3417 3122 3662 3127
rect 3417 3117 3422 3122
rect 3657 3117 3662 3122
rect 3737 3122 3766 3127
rect 3801 3122 4302 3127
rect 4577 3122 4606 3127
rect 3737 3117 3742 3122
rect 897 3112 926 3117
rect 969 3112 1038 3117
rect 1977 3112 2030 3117
rect 2113 3112 2142 3117
rect 2185 3112 2438 3117
rect 2457 3112 2526 3117
rect 2561 3112 2646 3117
rect 2841 3112 2870 3117
rect 3081 3112 3166 3117
rect 3225 3112 3286 3117
rect 3305 3112 3422 3117
rect 3513 3112 3630 3117
rect 3657 3112 3742 3117
rect 3785 3112 4342 3117
rect 4385 3112 4670 3117
rect 969 3107 974 3112
rect 209 3102 246 3107
rect 457 3102 486 3107
rect 585 3102 614 3107
rect 657 3102 726 3107
rect 945 3102 974 3107
rect 1033 3107 1038 3112
rect 1809 3107 1958 3112
rect 2937 3107 3062 3112
rect 1033 3102 1214 3107
rect 1609 3102 1814 3107
rect 1953 3102 2942 3107
rect 3057 3102 3214 3107
rect 3441 3102 3638 3107
rect 3769 3102 3846 3107
rect 3857 3102 3886 3107
rect 4009 3102 4270 3107
rect 4321 3102 4574 3107
rect 481 3097 590 3102
rect 305 3092 390 3097
rect 385 3087 390 3092
rect 761 3092 790 3097
rect 825 3092 934 3097
rect 761 3087 766 3092
rect 385 3082 766 3087
rect 929 3087 934 3092
rect 993 3092 1022 3097
rect 1505 3092 1606 3097
rect 1825 3092 1854 3097
rect 1905 3092 2478 3097
rect 2497 3092 2582 3097
rect 2953 3092 3118 3097
rect 993 3087 998 3092
rect 3113 3087 3118 3092
rect 3225 3092 3262 3097
rect 3457 3092 3486 3097
rect 3225 3087 3230 3092
rect 3481 3087 3486 3092
rect 3593 3092 3758 3097
rect 3897 3092 3998 3097
rect 4241 3092 4382 3097
rect 4681 3092 4766 3097
rect 3593 3087 3598 3092
rect 3753 3087 3902 3092
rect 3993 3087 4246 3092
rect 4377 3087 4478 3092
rect 4681 3087 4686 3092
rect 929 3082 998 3087
rect 1257 3082 1494 3087
rect 1489 3077 1494 3082
rect 1617 3082 1814 3087
rect 2241 3082 3070 3087
rect 3113 3082 3230 3087
rect 3273 3082 3406 3087
rect 3481 3082 3598 3087
rect 4265 3082 4358 3087
rect 4473 3082 4686 3087
rect 4737 3082 4774 3087
rect 1617 3077 1622 3082
rect 1809 3077 2246 3082
rect 1489 3072 1622 3077
rect 1721 3072 1750 3077
rect 1745 3067 1750 3072
rect 2265 3072 2470 3077
rect 2905 3072 3046 3077
rect 2265 3067 2270 3072
rect 2465 3067 2638 3072
rect 809 3062 1054 3067
rect 1073 3062 1110 3067
rect 1745 3062 2270 3067
rect 2289 3062 2310 3067
rect 2345 3062 2446 3067
rect 2633 3062 2734 3067
rect 265 3052 302 3057
rect 393 3052 678 3057
rect 809 3047 814 3062
rect 1049 3047 1054 3062
rect 2729 3057 2734 3062
rect 2905 3057 2910 3072
rect 3065 3067 3070 3082
rect 3273 3067 3278 3082
rect 3617 3072 4254 3077
rect 4369 3072 4454 3077
rect 4249 3067 4374 3072
rect 2929 3062 2974 3067
rect 3065 3062 3278 3067
rect 1129 3052 1198 3057
rect 1129 3047 1134 3052
rect 785 3042 814 3047
rect 833 3042 926 3047
rect 1049 3042 1134 3047
rect 1193 3047 1198 3052
rect 1545 3052 1702 3057
rect 2521 3052 2614 3057
rect 2729 3052 2910 3057
rect 3489 3052 3526 3057
rect 3753 3052 3790 3057
rect 3833 3052 3886 3057
rect 3945 3052 4110 3057
rect 4177 3052 4622 3057
rect 1545 3047 1550 3052
rect 1193 3042 1550 3047
rect 1697 3047 1702 3052
rect 1697 3042 2094 3047
rect 2177 3042 2238 3047
rect 3121 3042 3222 3047
rect 833 3037 838 3042
rect 113 3032 190 3037
rect 665 3032 838 3037
rect 921 3037 926 3042
rect 2569 3037 2686 3042
rect 3121 3037 3126 3042
rect 921 3032 1182 3037
rect 1641 3032 1670 3037
rect 2225 3032 2374 3037
rect 2545 3032 2574 3037
rect 2681 3032 2710 3037
rect 3097 3032 3126 3037
rect 3217 3037 3222 3042
rect 3569 3042 3654 3047
rect 3865 3042 3926 3047
rect 4089 3042 4166 3047
rect 4313 3042 4342 3047
rect 3569 3037 3574 3042
rect 3217 3032 3246 3037
rect 3545 3032 3574 3037
rect 3649 3037 3654 3042
rect 3961 3037 4070 3042
rect 4161 3037 4318 3042
rect 3649 3032 3862 3037
rect 3937 3032 3966 3037
rect 4065 3032 4118 3037
rect 4345 3032 4430 3037
rect 4489 3032 4542 3037
rect 97 3022 134 3027
rect 241 3022 318 3027
rect 361 3022 406 3027
rect 793 3022 830 3027
rect 873 3022 910 3027
rect 1033 3022 1102 3027
rect 1561 3022 1686 3027
rect 1889 3022 2086 3027
rect 2153 3022 2198 3027
rect 2281 3022 2310 3027
rect 2601 3022 2646 3027
rect 2833 3022 2862 3027
rect 2889 3022 2910 3027
rect 3025 3022 3222 3027
rect 3657 3022 4182 3027
rect 4233 3022 4342 3027
rect 4409 3022 4454 3027
rect 4337 3017 4342 3022
rect 4449 3017 4454 3022
rect 4553 3022 4630 3027
rect 4553 3017 4558 3022
rect 137 3012 222 3017
rect 313 3012 390 3017
rect 945 3012 1286 3017
rect 1497 3012 1630 3017
rect 1865 3012 1886 3017
rect 2209 3012 2398 3017
rect 2673 3012 2694 3017
rect 2825 3012 2926 3017
rect 3009 3012 3038 3017
rect 3201 3012 3390 3017
rect 3569 3012 3702 3017
rect 3737 3012 4046 3017
rect 4161 3012 4190 3017
rect 4337 3012 4382 3017
rect 4449 3012 4558 3017
rect 1953 3007 2214 3012
rect 2673 3007 2678 3012
rect 3033 3007 3206 3012
rect 4041 3007 4166 3012
rect 185 3002 342 3007
rect 425 3002 926 3007
rect 1417 3002 1670 3007
rect 1929 3002 1958 3007
rect 2361 3002 2390 3007
rect 2417 3002 2518 3007
rect 2537 3002 2678 3007
rect 2737 3002 2870 3007
rect 3233 3002 3310 3007
rect 3985 3002 4022 3007
rect 4209 3002 4318 3007
rect 425 2997 430 3002
rect 945 2997 1118 3002
rect 2417 2997 2422 3002
rect 121 2992 150 2997
rect 273 2992 430 2997
rect 897 2992 950 2997
rect 1113 2992 1142 2997
rect 1201 2992 1398 2997
rect 1481 2992 1526 2997
rect 1769 2992 1838 2997
rect 1913 2992 2070 2997
rect 2081 2992 2230 2997
rect 2257 2992 2422 2997
rect 2513 2997 2518 3002
rect 2737 2997 2742 3002
rect 3817 2997 3966 3002
rect 4209 2997 4214 3002
rect 2513 2992 2742 2997
rect 3033 2992 3134 2997
rect 3177 2992 3286 2997
rect 3529 2992 3598 2997
rect 3681 2992 3782 2997
rect 3793 2992 3822 2997
rect 3961 2992 4214 2997
rect 4313 2997 4318 3002
rect 4313 2992 4366 2997
rect 4393 2992 4430 2997
rect 4593 2992 4630 2997
rect 4657 2992 4694 2997
rect 777 2987 878 2992
rect 1201 2987 1206 2992
rect 233 2982 302 2987
rect 449 2982 638 2987
rect 657 2982 782 2987
rect 873 2982 1166 2987
rect 1177 2982 1206 2987
rect 1393 2987 1398 2992
rect 1545 2987 1742 2992
rect 3793 2987 3798 2992
rect 1393 2982 1550 2987
rect 1737 2982 1782 2987
rect 1825 2982 2038 2987
rect 2073 2982 2862 2987
rect 3585 2982 3798 2987
rect 3833 2982 3942 2987
rect 4081 2982 4590 2987
rect 321 2977 454 2982
rect 633 2977 638 2982
rect 4001 2977 4086 2982
rect 4585 2977 4590 2982
rect 4649 2982 4702 2987
rect 4649 2977 4654 2982
rect 193 2972 326 2977
rect 633 2972 774 2977
rect 785 2972 894 2977
rect 473 2967 614 2972
rect 785 2967 790 2972
rect 169 2962 310 2967
rect 337 2962 478 2967
rect 609 2962 790 2967
rect 889 2967 894 2972
rect 977 2972 1710 2977
rect 977 2967 982 2972
rect 1705 2967 1710 2972
rect 1785 2972 1918 2977
rect 2017 2972 2078 2977
rect 2121 2972 2142 2977
rect 2169 2972 2198 2977
rect 2329 2972 2374 2977
rect 2393 2972 2830 2977
rect 3305 2972 3334 2977
rect 3609 2972 4006 2977
rect 4105 2972 4190 2977
rect 4209 2972 4310 2977
rect 1785 2967 1790 2972
rect 2217 2967 2310 2972
rect 4305 2967 4310 2972
rect 4377 2972 4406 2977
rect 4585 2972 4654 2977
rect 4377 2967 4382 2972
rect 889 2962 982 2967
rect 1033 2962 1062 2967
rect 1337 2962 1470 2967
rect 1705 2962 1790 2967
rect 1809 2962 2222 2967
rect 2305 2962 2358 2967
rect 2481 2962 3438 2967
rect 3609 2962 3782 2967
rect 4017 2962 4094 2967
rect 4185 2962 4214 2967
rect 4305 2962 4382 2967
rect 4425 2962 4566 2967
rect 1057 2957 1342 2962
rect 1465 2957 1654 2962
rect 185 2952 630 2957
rect 649 2952 694 2957
rect 801 2952 870 2957
rect 1361 2952 1446 2957
rect 689 2947 806 2952
rect 1649 2947 1654 2957
rect 1809 2947 1814 2962
rect 2353 2957 2486 2962
rect 3777 2957 3782 2962
rect 3905 2957 4022 2962
rect 4089 2957 4190 2962
rect 4425 2957 4430 2962
rect 1897 2952 1934 2957
rect 2033 2952 2334 2957
rect 2505 2952 2558 2957
rect 2609 2952 2846 2957
rect 3361 2952 3382 2957
rect 3465 2952 3606 2957
rect 3713 2952 3758 2957
rect 3777 2952 3910 2957
rect 4217 2952 4270 2957
rect 4401 2952 4430 2957
rect 4561 2947 4566 2962
rect 4681 2952 4718 2957
rect 401 2942 518 2947
rect 641 2942 670 2947
rect 1001 2942 1310 2947
rect 1489 2942 1630 2947
rect 1649 2942 1814 2947
rect 2001 2942 2286 2947
rect 513 2937 646 2942
rect 2281 2937 2286 2942
rect 2345 2942 2854 2947
rect 3377 2942 3502 2947
rect 3617 2942 3710 2947
rect 3929 2942 4006 2947
rect 4129 2942 4150 2947
rect 4233 2942 4390 2947
rect 4521 2942 4550 2947
rect 4561 2942 4694 2947
rect 2345 2937 2350 2942
rect 3929 2937 3934 2942
rect 369 2932 414 2937
rect 769 2932 814 2937
rect 1337 2932 1390 2937
rect 1553 2932 1582 2937
rect 1873 2932 2142 2937
rect 2193 2932 2262 2937
rect 2281 2932 2350 2937
rect 2473 2932 2502 2937
rect 2497 2927 2502 2932
rect 2577 2932 2774 2937
rect 3489 2932 3590 2937
rect 3777 2932 3886 2937
rect 3905 2932 3934 2937
rect 4001 2937 4006 2942
rect 4385 2937 4462 2942
rect 4521 2937 4526 2942
rect 4001 2932 4030 2937
rect 4225 2932 4254 2937
rect 4321 2932 4358 2937
rect 4457 2932 4526 2937
rect 4785 2932 4806 2937
rect 2577 2927 2582 2932
rect 3777 2927 3782 2932
rect 433 2922 478 2927
rect 561 2922 646 2927
rect 681 2922 726 2927
rect 1393 2922 1510 2927
rect 1833 2922 1862 2927
rect 1985 2922 2022 2927
rect 2113 2922 2206 2927
rect 2497 2922 2582 2927
rect 2601 2922 2926 2927
rect 3553 2922 3598 2927
rect 3633 2922 3782 2927
rect 3881 2927 3886 2932
rect 4121 2927 4206 2932
rect 3881 2922 4126 2927
rect 4201 2922 4238 2927
rect 4385 2922 4438 2927
rect 4761 2922 4782 2927
rect 561 2917 566 2922
rect 465 2912 566 2917
rect 641 2917 646 2922
rect 761 2917 886 2922
rect 1305 2917 1374 2922
rect 4257 2917 4350 2922
rect 641 2912 670 2917
rect 665 2907 670 2912
rect 737 2912 766 2917
rect 881 2912 1094 2917
rect 1145 2912 1310 2917
rect 1369 2912 1430 2917
rect 1521 2912 1974 2917
rect 2057 2912 2086 2917
rect 2137 2912 2406 2917
rect 2665 2912 2710 2917
rect 2865 2912 2918 2917
rect 3089 2912 3206 2917
rect 3329 2912 3590 2917
rect 3793 2912 3870 2917
rect 4137 2912 4262 2917
rect 4345 2912 4406 2917
rect 4425 2912 4470 2917
rect 4537 2912 4790 2917
rect 737 2907 742 2912
rect 1425 2907 1526 2912
rect 1969 2907 2062 2912
rect 3585 2907 3798 2912
rect 3865 2907 3966 2912
rect 4137 2907 4142 2912
rect 233 2902 270 2907
rect 305 2902 454 2907
rect 577 2902 630 2907
rect 665 2902 742 2907
rect 785 2902 870 2907
rect 1089 2902 1190 2907
rect 1321 2902 1406 2907
rect 2337 2902 2542 2907
rect 2633 2902 2662 2907
rect 449 2897 582 2902
rect 625 2887 630 2902
rect 785 2887 790 2902
rect 2657 2897 2662 2902
rect 2753 2902 2902 2907
rect 2929 2902 2974 2907
rect 3305 2902 3326 2907
rect 3505 2902 3566 2907
rect 3961 2902 4142 2907
rect 4209 2902 4334 2907
rect 2753 2897 2758 2902
rect 4329 2897 4334 2902
rect 4417 2902 4478 2907
rect 4417 2897 4422 2902
rect 889 2892 1070 2897
rect 1209 2892 1294 2897
rect 1401 2892 2198 2897
rect 2217 2892 2254 2897
rect 2657 2892 2758 2897
rect 3177 2892 3334 2897
rect 3353 2892 3486 2897
rect 889 2887 894 2892
rect 1065 2887 1214 2892
rect 1289 2887 1294 2892
rect 3353 2887 3358 2892
rect 297 2882 358 2887
rect 353 2877 358 2882
rect 505 2882 534 2887
rect 625 2882 790 2887
rect 809 2882 894 2887
rect 1289 2882 1318 2887
rect 1801 2882 1830 2887
rect 2841 2882 3038 2887
rect 3057 2882 3358 2887
rect 3481 2887 3486 2892
rect 3585 2892 3942 2897
rect 4329 2892 4422 2897
rect 3585 2887 3590 2892
rect 3481 2882 3590 2887
rect 3937 2887 3942 2892
rect 3937 2882 4046 2887
rect 505 2877 510 2882
rect 1337 2877 1486 2882
rect 2841 2877 2846 2882
rect 353 2872 510 2877
rect 865 2872 1342 2877
rect 1481 2872 2502 2877
rect 2777 2872 2846 2877
rect 3033 2877 3038 2882
rect 3609 2877 3838 2882
rect 3033 2872 3614 2877
rect 3833 2872 4286 2877
rect 2881 2867 3014 2872
rect 1049 2862 1470 2867
rect 1753 2862 1782 2867
rect 2857 2862 2886 2867
rect 3009 2862 3822 2867
rect 4081 2862 4110 2867
rect 4369 2862 4486 2867
rect 3817 2857 4086 2862
rect 4369 2857 4374 2862
rect 81 2852 310 2857
rect 625 2852 1214 2857
rect 1577 2852 1726 2857
rect 1745 2852 1790 2857
rect 1817 2852 1894 2857
rect 2625 2852 2702 2857
rect 2833 2852 3798 2857
rect 4345 2852 4374 2857
rect 4481 2857 4486 2862
rect 4481 2852 4510 2857
rect 1305 2847 1502 2852
rect 1577 2847 1582 2852
rect 1001 2842 1310 2847
rect 1497 2842 1582 2847
rect 1721 2847 1726 2852
rect 2625 2847 2630 2852
rect 1721 2842 1846 2847
rect 1905 2842 2630 2847
rect 2697 2847 2702 2852
rect 2697 2842 2822 2847
rect 1841 2837 1910 2842
rect 2817 2837 2822 2842
rect 2897 2842 2990 2847
rect 3177 2842 3718 2847
rect 3865 2842 4254 2847
rect 2897 2837 2902 2842
rect 2985 2837 3094 2842
rect 3177 2837 3182 2842
rect 521 2832 574 2837
rect 689 2832 726 2837
rect 993 2832 1038 2837
rect 1121 2832 1222 2837
rect 1033 2827 1126 2832
rect 1217 2827 1222 2832
rect 1321 2832 1406 2837
rect 1417 2832 1486 2837
rect 1321 2827 1326 2832
rect 1481 2827 1486 2832
rect 1593 2832 1822 2837
rect 2817 2832 2902 2837
rect 2937 2832 2966 2837
rect 3089 2832 3182 2837
rect 3201 2832 3254 2837
rect 3561 2832 3662 2837
rect 4313 2832 4374 2837
rect 4385 2832 4558 2837
rect 1593 2827 1598 2832
rect 3353 2827 3462 2832
rect 3921 2827 4134 2832
rect 353 2822 398 2827
rect 489 2822 534 2827
rect 577 2822 694 2827
rect 849 2822 902 2827
rect 201 2812 334 2817
rect 665 2812 878 2817
rect 201 2797 206 2812
rect 177 2792 206 2797
rect 329 2797 334 2812
rect 1009 2802 1014 2827
rect 1145 2822 1198 2827
rect 1217 2822 1326 2827
rect 1345 2822 1462 2827
rect 1481 2822 1598 2827
rect 1617 2822 1678 2827
rect 1801 2822 1846 2827
rect 2057 2822 2102 2827
rect 2313 2822 2422 2827
rect 2433 2822 2486 2827
rect 2641 2822 2686 2827
rect 2921 2822 2958 2827
rect 3025 2822 3070 2827
rect 3209 2822 3254 2827
rect 3329 2822 3358 2827
rect 3457 2822 3550 2827
rect 3617 2822 3646 2827
rect 3705 2822 3926 2827
rect 4129 2822 4350 2827
rect 4657 2822 4726 2827
rect 3545 2817 3622 2822
rect 4369 2817 4542 2822
rect 1129 2812 1174 2817
rect 2129 2812 2294 2817
rect 2401 2812 2494 2817
rect 2569 2812 2630 2817
rect 2705 2812 2790 2817
rect 2857 2812 2894 2817
rect 3057 2812 3198 2817
rect 3265 2812 3446 2817
rect 3809 2812 3838 2817
rect 3937 2812 4158 2817
rect 4257 2812 4374 2817
rect 4537 2812 4566 2817
rect 1777 2802 1806 2807
rect 2129 2797 2134 2812
rect 329 2792 446 2797
rect 753 2792 1782 2797
rect 1825 2792 1894 2797
rect 2105 2792 2134 2797
rect 2289 2797 2294 2812
rect 2625 2807 2710 2812
rect 3193 2807 3270 2812
rect 3833 2807 3942 2812
rect 4153 2807 4262 2812
rect 2361 2802 2502 2807
rect 2809 2802 2918 2807
rect 2945 2802 2998 2807
rect 3337 2802 3630 2807
rect 3961 2802 4014 2807
rect 4089 2802 4134 2807
rect 4281 2802 4534 2807
rect 2521 2797 2598 2802
rect 2289 2792 2526 2797
rect 2593 2792 2678 2797
rect 3161 2792 3262 2797
rect 3377 2792 3430 2797
rect 3601 2792 3846 2797
rect 4041 2792 4070 2797
rect 4145 2792 4270 2797
rect 4393 2792 4422 2797
rect 4473 2792 4590 2797
rect 1825 2787 1830 2792
rect 209 2782 294 2787
rect 305 2782 350 2787
rect 617 2782 758 2787
rect 1753 2782 1830 2787
rect 1889 2787 1894 2792
rect 2673 2787 2678 2792
rect 4065 2787 4150 2792
rect 4265 2787 4398 2792
rect 1889 2782 2014 2787
rect 2097 2782 2134 2787
rect 2185 2782 2486 2787
rect 2545 2782 2582 2787
rect 2673 2782 2750 2787
rect 2785 2782 2870 2787
rect 3281 2782 3326 2787
rect 4449 2782 4550 2787
rect 2785 2777 2790 2782
rect 385 2772 406 2777
rect 849 2772 1086 2777
rect 1137 2772 1174 2777
rect 1185 2772 1222 2777
rect 1401 2772 1470 2777
rect 1625 2772 1742 2777
rect 1809 2772 2086 2777
rect 2185 2772 2494 2777
rect 1737 2767 1814 2772
rect 2081 2767 2190 2772
rect 2489 2767 2494 2772
rect 2593 2772 2662 2777
rect 2593 2767 2598 2772
rect 649 2762 846 2767
rect 945 2762 974 2767
rect 1041 2762 1078 2767
rect 1273 2762 1302 2767
rect 2209 2762 2382 2767
rect 2425 2762 2470 2767
rect 2489 2762 2598 2767
rect 2657 2767 2662 2772
rect 2761 2772 2790 2777
rect 2865 2777 2870 2782
rect 2865 2772 3062 2777
rect 3081 2772 3190 2777
rect 3433 2772 4350 2777
rect 4433 2772 4646 2777
rect 2761 2767 2766 2772
rect 3081 2767 3086 2772
rect 2657 2762 2766 2767
rect 2801 2762 2854 2767
rect 3033 2762 3086 2767
rect 3185 2767 3190 2772
rect 3185 2762 3214 2767
rect 3921 2762 3950 2767
rect 4401 2762 4438 2767
rect 841 2757 950 2762
rect 1097 2757 1190 2762
rect 1553 2757 1678 2762
rect 1833 2757 1982 2762
rect 3665 2757 3926 2762
rect 4105 2757 4174 2762
rect 4433 2757 4438 2762
rect 4529 2762 4630 2767
rect 4529 2757 4534 2762
rect 233 2752 366 2757
rect 401 2752 670 2757
rect 793 2752 822 2757
rect 817 2747 822 2752
rect 985 2752 1102 2757
rect 1185 2752 1558 2757
rect 1673 2752 1838 2757
rect 1977 2752 2190 2757
rect 2233 2752 2310 2757
rect 2369 2752 2422 2757
rect 2905 2752 3502 2757
rect 3641 2752 3670 2757
rect 3953 2752 4110 2757
rect 4169 2752 4238 2757
rect 4433 2752 4534 2757
rect 4561 2752 4598 2757
rect 985 2747 990 2752
rect 129 2742 318 2747
rect 641 2742 678 2747
rect 817 2742 990 2747
rect 1049 2742 1174 2747
rect 1569 2742 1662 2747
rect 1849 2742 1878 2747
rect 1929 2742 2038 2747
rect 2401 2742 2446 2747
rect 2489 2742 2638 2747
rect 2657 2742 2806 2747
rect 3049 2742 3078 2747
rect 3169 2742 3198 2747
rect 3209 2742 3230 2747
rect 3449 2742 3598 2747
rect 3609 2742 3662 2747
rect 3721 2742 3838 2747
rect 3873 2742 3982 2747
rect 4041 2742 4062 2747
rect 4073 2742 4158 2747
rect 4289 2742 4414 2747
rect 4553 2742 4614 2747
rect 4657 2742 4718 2747
rect 1289 2737 1358 2742
rect 177 2732 222 2737
rect 1265 2732 1294 2737
rect 1353 2732 1462 2737
rect 1873 2727 1878 2742
rect 2489 2737 2494 2742
rect 1897 2732 1942 2737
rect 2129 2732 2494 2737
rect 2633 2737 2638 2742
rect 3321 2737 3430 2742
rect 4289 2737 4294 2742
rect 2633 2732 2686 2737
rect 2817 2732 3078 2737
rect 3297 2732 3326 2737
rect 3425 2732 3638 2737
rect 3769 2732 3894 2737
rect 3905 2732 3990 2737
rect 4041 2732 4294 2737
rect 2681 2727 2822 2732
rect 3073 2727 3078 2732
rect 3905 2727 3910 2732
rect 145 2722 350 2727
rect 689 2722 774 2727
rect 873 2722 926 2727
rect 961 2722 1070 2727
rect 1193 2722 1342 2727
rect 1449 2722 1686 2727
rect 1705 2722 1830 2727
rect 1873 2722 1982 2727
rect 2393 2722 2446 2727
rect 2625 2722 2662 2727
rect 3073 2722 3270 2727
rect 1705 2717 1710 2722
rect 89 2712 142 2717
rect 185 2712 246 2717
rect 281 2712 350 2717
rect 369 2712 478 2717
rect 497 2712 670 2717
rect 713 2712 774 2717
rect 785 2712 862 2717
rect 121 2702 150 2707
rect 265 2702 406 2707
rect 145 2697 270 2702
rect 497 2697 502 2712
rect 665 2702 670 2712
rect 785 2702 790 2712
rect 857 2707 862 2712
rect 937 2712 1238 2717
rect 1353 2712 1510 2717
rect 1601 2712 1710 2717
rect 1825 2717 1830 2722
rect 3361 2717 3366 2727
rect 3401 2722 3614 2727
rect 3745 2722 3774 2727
rect 3769 2717 3774 2722
rect 3857 2722 3910 2727
rect 3985 2727 3990 2732
rect 4577 2727 4582 2742
rect 4665 2732 4790 2737
rect 3985 2722 4094 2727
rect 4289 2722 4382 2727
rect 4417 2722 4558 2727
rect 4577 2722 4622 2727
rect 3857 2717 3862 2722
rect 1825 2712 1918 2717
rect 1993 2712 2286 2717
rect 2313 2712 2630 2717
rect 2641 2712 2686 2717
rect 2761 2712 2862 2717
rect 3233 2712 3366 2717
rect 3513 2712 3550 2717
rect 3769 2712 3862 2717
rect 3881 2712 3910 2717
rect 3953 2712 4046 2717
rect 4113 2712 4270 2717
rect 4665 2712 4734 2717
rect 937 2707 942 2712
rect 1233 2707 1358 2712
rect 1505 2707 1606 2712
rect 1913 2707 1998 2712
rect 2761 2707 2766 2712
rect 857 2702 942 2707
rect 993 2702 1086 2707
rect 1185 2702 1214 2707
rect 1417 2702 1486 2707
rect 1625 2702 1726 2707
rect 1849 2702 1894 2707
rect 2553 2702 2766 2707
rect 2857 2707 2862 2712
rect 3049 2707 3174 2712
rect 4113 2707 4118 2712
rect 4265 2707 4382 2712
rect 2857 2702 2886 2707
rect 2905 2702 3006 2707
rect 3025 2702 3054 2707
rect 3169 2702 3246 2707
rect 3465 2702 3526 2707
rect 3889 2702 4014 2707
rect 4089 2702 4118 2707
rect 4377 2702 4406 2707
rect 4553 2702 4646 2707
rect 665 2697 790 2702
rect 2049 2697 2118 2702
rect 2185 2697 2374 2702
rect 2905 2697 2910 2702
rect 289 2692 326 2697
rect 473 2692 502 2697
rect 961 2692 1406 2697
rect 1401 2687 1406 2692
rect 1497 2692 1614 2697
rect 1497 2687 1502 2692
rect 217 2682 798 2687
rect 881 2682 942 2687
rect 1033 2682 1062 2687
rect 1401 2682 1502 2687
rect 1609 2687 1614 2692
rect 1697 2692 1838 2697
rect 1697 2687 1702 2692
rect 1833 2687 1838 2692
rect 1905 2692 2054 2697
rect 2113 2692 2190 2697
rect 2369 2692 2542 2697
rect 2753 2692 2910 2697
rect 3001 2697 3006 2702
rect 3265 2697 3430 2702
rect 4137 2697 4214 2702
rect 3001 2692 3270 2697
rect 3425 2692 4142 2697
rect 4209 2692 4310 2697
rect 4361 2692 4470 2697
rect 1905 2687 1910 2692
rect 2537 2687 2758 2692
rect 1609 2682 1702 2687
rect 1721 2682 1806 2687
rect 1833 2682 1910 2687
rect 2065 2682 2102 2687
rect 2097 2677 2102 2682
rect 2201 2682 2358 2687
rect 2777 2682 3414 2687
rect 3489 2682 3574 2687
rect 3945 2682 4030 2687
rect 4145 2682 4198 2687
rect 2201 2677 2206 2682
rect 657 2672 694 2677
rect 745 2672 1118 2677
rect 1137 2672 1230 2677
rect 2017 2672 2078 2677
rect 2097 2672 2206 2677
rect 2225 2672 2254 2677
rect 2369 2672 2766 2677
rect 2849 2672 3302 2677
rect 3473 2672 3518 2677
rect 3785 2672 3910 2677
rect 3929 2672 4086 2677
rect 4249 2672 4510 2677
rect 2249 2667 2374 2672
rect 2761 2667 2854 2672
rect 3785 2667 3790 2672
rect 753 2662 1094 2667
rect 1249 2662 1702 2667
rect 1249 2657 1254 2662
rect 321 2652 646 2657
rect 969 2652 1254 2657
rect 1697 2657 1702 2662
rect 1849 2662 1998 2667
rect 2993 2662 3350 2667
rect 3593 2662 3742 2667
rect 3761 2662 3790 2667
rect 3905 2667 3910 2672
rect 3905 2662 3958 2667
rect 4177 2662 4246 2667
rect 1849 2657 1854 2662
rect 1993 2657 2094 2662
rect 2873 2657 2974 2662
rect 3593 2657 3598 2662
rect 1697 2652 1854 2657
rect 2089 2652 2118 2657
rect 2137 2652 2582 2657
rect 2761 2652 2878 2657
rect 2969 2652 3158 2657
rect 3249 2652 3486 2657
rect 3497 2652 3598 2657
rect 3737 2657 3742 2662
rect 3737 2652 4166 2657
rect 641 2647 646 2652
rect 841 2647 974 2652
rect 1345 2647 1558 2652
rect 2137 2647 2142 2652
rect 641 2642 846 2647
rect 993 2642 1022 2647
rect 1105 2642 1142 2647
rect 1321 2642 1350 2647
rect 1553 2642 1638 2647
rect 1945 2642 2142 2647
rect 2577 2647 2582 2652
rect 3153 2647 3254 2652
rect 4161 2647 4166 2652
rect 4249 2652 4350 2657
rect 4401 2652 4454 2657
rect 4249 2647 4254 2652
rect 2577 2642 2606 2647
rect 2625 2642 2742 2647
rect 2889 2642 3038 2647
rect 3521 2642 3870 2647
rect 4161 2642 4254 2647
rect 4473 2642 4614 2647
rect 321 2637 574 2642
rect 1161 2637 1278 2642
rect 2257 2637 2342 2642
rect 2625 2637 2630 2642
rect 297 2632 326 2637
rect 569 2632 598 2637
rect 865 2632 1166 2637
rect 1273 2632 1542 2637
rect 1649 2632 2086 2637
rect 2153 2632 2262 2637
rect 2337 2632 2630 2637
rect 2737 2637 2742 2642
rect 3057 2637 3134 2642
rect 3273 2637 3342 2642
rect 3945 2637 4094 2642
rect 4473 2637 4478 2642
rect 2737 2632 3062 2637
rect 3129 2632 3278 2637
rect 3337 2632 3590 2637
rect 1537 2627 1654 2632
rect 2081 2627 2158 2632
rect 3585 2627 3590 2632
rect 3705 2632 3950 2637
rect 4089 2632 4118 2637
rect 4273 2632 4342 2637
rect 4401 2632 4478 2637
rect 3705 2627 3710 2632
rect 4113 2627 4118 2632
rect 4401 2627 4406 2632
rect 81 2622 182 2627
rect 297 2622 342 2627
rect 361 2622 614 2627
rect 785 2622 894 2627
rect 929 2622 950 2627
rect 1073 2622 1118 2627
rect 1169 2622 1262 2627
rect 1345 2622 1398 2627
rect 1489 2622 1518 2627
rect 1889 2622 1934 2627
rect 2017 2622 2062 2627
rect 2273 2622 2326 2627
rect 2593 2622 2726 2627
rect 2937 2622 2998 2627
rect 3017 2622 3118 2627
rect 3289 2622 3326 2627
rect 3457 2622 3566 2627
rect 3585 2622 3710 2627
rect 3745 2622 3838 2627
rect 3961 2622 4094 2627
rect 4113 2622 4254 2627
rect 4353 2622 4406 2627
rect 4609 2627 4614 2642
rect 4609 2622 4638 2627
rect 4689 2622 4710 2627
rect 2377 2617 2558 2622
rect 345 2612 374 2617
rect 481 2612 510 2617
rect 369 2607 486 2612
rect 153 2592 190 2597
rect 425 2592 502 2597
rect 577 2592 582 2617
rect 945 2612 966 2617
rect 665 2602 862 2607
rect 665 2597 670 2602
rect 641 2592 670 2597
rect 857 2597 862 2602
rect 1025 2597 1030 2617
rect 1281 2612 1334 2617
rect 1617 2612 1686 2617
rect 1977 2612 2038 2617
rect 2081 2612 2182 2617
rect 2201 2612 2382 2617
rect 2553 2612 2582 2617
rect 1097 2607 1198 2612
rect 1617 2607 1622 2612
rect 1073 2602 1102 2607
rect 1193 2602 1622 2607
rect 1681 2607 1686 2612
rect 2081 2607 2086 2612
rect 1681 2602 1710 2607
rect 1729 2602 1870 2607
rect 1729 2597 1734 2602
rect 857 2592 886 2597
rect 1025 2592 1046 2597
rect 1105 2592 1182 2597
rect 1265 2592 1334 2597
rect 1633 2592 1734 2597
rect 1865 2597 1870 2602
rect 1985 2602 2086 2607
rect 2177 2607 2182 2612
rect 2593 2607 2598 2622
rect 2721 2617 2942 2622
rect 2993 2617 2998 2622
rect 3457 2617 3462 2622
rect 2961 2612 2982 2617
rect 2993 2612 3038 2617
rect 3129 2612 3254 2617
rect 3385 2612 3462 2617
rect 3473 2612 3502 2617
rect 3729 2612 3758 2617
rect 3857 2612 3982 2617
rect 4225 2612 4334 2617
rect 2177 2602 2294 2607
rect 1985 2597 1990 2602
rect 2289 2597 2294 2602
rect 2393 2602 2598 2607
rect 2617 2602 2702 2607
rect 2817 2602 2862 2607
rect 2961 2602 2966 2612
rect 3033 2607 3134 2612
rect 4329 2607 4334 2612
rect 4417 2612 4446 2617
rect 4489 2612 4646 2617
rect 4417 2607 4422 2612
rect 2977 2602 3014 2607
rect 4073 2602 4182 2607
rect 4329 2602 4422 2607
rect 4705 2602 4710 2622
rect 2393 2597 2398 2602
rect 1865 2592 1990 2597
rect 2033 2592 2230 2597
rect 2241 2592 2270 2597
rect 2289 2592 2398 2597
rect 2417 2592 2462 2597
rect 2545 2592 2670 2597
rect 2681 2592 2766 2597
rect 3057 2592 3214 2597
rect 3361 2592 3422 2597
rect 3529 2592 3574 2597
rect 3593 2592 3710 2597
rect 3985 2592 4038 2597
rect 4113 2592 4182 2597
rect 4625 2592 4694 2597
rect 425 2587 430 2592
rect 113 2582 294 2587
rect 313 2582 430 2587
rect 497 2587 502 2592
rect 1353 2587 1510 2592
rect 3593 2587 3598 2592
rect 497 2582 614 2587
rect 289 2567 294 2582
rect 609 2577 614 2582
rect 681 2582 1358 2587
rect 1505 2582 1806 2587
rect 1985 2582 2014 2587
rect 2217 2582 2254 2587
rect 2425 2582 2710 2587
rect 2745 2582 2846 2587
rect 2889 2582 2918 2587
rect 3401 2582 3598 2587
rect 3705 2587 3710 2592
rect 3705 2582 3974 2587
rect 4057 2582 4142 2587
rect 4273 2582 4310 2587
rect 681 2577 686 2582
rect 1825 2577 1926 2582
rect 2113 2577 2198 2582
rect 441 2572 486 2577
rect 609 2572 686 2577
rect 793 2572 830 2577
rect 881 2572 950 2577
rect 1017 2572 1494 2577
rect 1577 2572 1614 2577
rect 1705 2572 1830 2577
rect 1921 2572 2118 2577
rect 2193 2572 2294 2577
rect 2305 2572 2334 2577
rect 2577 2572 3230 2577
rect 3249 2572 3342 2577
rect 4065 2572 4134 2577
rect 4577 2572 4646 2577
rect 1489 2567 1582 2572
rect 2289 2567 2294 2572
rect 3249 2567 3254 2572
rect 3337 2567 3510 2572
rect 3761 2567 3894 2572
rect 289 2562 590 2567
rect 921 2562 1022 2567
rect 1065 2562 1318 2567
rect 1689 2562 1766 2567
rect 1825 2562 1910 2567
rect 2129 2562 2262 2567
rect 2289 2562 2310 2567
rect 2433 2562 2870 2567
rect 2889 2562 2926 2567
rect 3217 2562 3254 2567
rect 3505 2562 3726 2567
rect 3737 2562 3766 2567
rect 3889 2562 4054 2567
rect 1337 2557 1470 2562
rect 1601 2557 1670 2562
rect 1961 2557 2110 2562
rect 2945 2557 3182 2562
rect 4049 2557 4054 2562
rect 4145 2562 4230 2567
rect 4641 2562 4742 2567
rect 4145 2557 4150 2562
rect 161 2552 278 2557
rect 273 2537 278 2552
rect 481 2552 678 2557
rect 825 2552 1086 2557
rect 1097 2552 1118 2557
rect 1193 2552 1342 2557
rect 1465 2552 1606 2557
rect 1665 2552 1742 2557
rect 481 2537 486 2552
rect 1737 2547 1742 2552
rect 1849 2552 1966 2557
rect 2105 2552 2158 2557
rect 1849 2547 1854 2552
rect 2153 2547 2158 2552
rect 2265 2552 2422 2557
rect 2593 2552 2950 2557
rect 3177 2552 3206 2557
rect 2265 2547 2270 2552
rect 2417 2547 2598 2552
rect 3201 2547 3206 2552
rect 3265 2552 3494 2557
rect 3753 2552 3790 2557
rect 3833 2552 3878 2557
rect 4049 2552 4150 2557
rect 4329 2552 4366 2557
rect 3265 2547 3270 2552
rect 561 2542 614 2547
rect 665 2542 814 2547
rect 1065 2542 1134 2547
rect 1281 2542 1310 2547
rect 1361 2542 1454 2547
rect 1617 2542 1718 2547
rect 1737 2542 1854 2547
rect 1873 2542 1902 2547
rect 1977 2542 2134 2547
rect 2153 2542 2270 2547
rect 2881 2542 2926 2547
rect 2945 2542 3158 2547
rect 3201 2542 3270 2547
rect 3313 2542 3414 2547
rect 4241 2542 4342 2547
rect 4353 2542 4470 2547
rect 4553 2542 4654 2547
rect 4681 2542 4734 2547
rect 273 2532 486 2537
rect 809 2537 814 2542
rect 873 2537 1070 2542
rect 2617 2537 2838 2542
rect 2945 2537 2950 2542
rect 809 2532 878 2537
rect 1089 2532 1134 2537
rect 2289 2532 2366 2537
rect 2489 2532 2622 2537
rect 2833 2532 2950 2537
rect 3409 2537 3414 2542
rect 3409 2532 3726 2537
rect 3897 2532 4126 2537
rect 4409 2532 4446 2537
rect 4633 2532 4678 2537
rect 1945 2527 2030 2532
rect 2969 2527 3238 2532
rect 3297 2527 3366 2532
rect 4145 2527 4270 2532
rect 585 2522 718 2527
rect 713 2517 718 2522
rect 897 2522 1038 2527
rect 1097 2522 1126 2527
rect 1281 2522 1950 2527
rect 2025 2522 2478 2527
rect 2633 2522 2822 2527
rect 2905 2522 2974 2527
rect 3233 2522 3302 2527
rect 3361 2522 3390 2527
rect 4113 2522 4150 2527
rect 4265 2522 4310 2527
rect 897 2517 902 2522
rect 209 2512 254 2517
rect 505 2512 574 2517
rect 665 2512 694 2517
rect 713 2512 902 2517
rect 1049 2512 1078 2517
rect 1089 2512 1142 2517
rect 1161 2512 1262 2517
rect 1281 2512 1286 2522
rect 2473 2517 2638 2522
rect 4673 2517 4774 2522
rect 1961 2512 2014 2517
rect 2657 2512 2702 2517
rect 2969 2512 3006 2517
rect 3041 2512 3198 2517
rect 3313 2512 3342 2517
rect 3673 2512 3782 2517
rect 3817 2512 3910 2517
rect 4137 2512 4350 2517
rect 4601 2512 4638 2517
rect 4649 2512 4678 2517
rect 4769 2512 4798 2517
rect 1161 2507 1166 2512
rect 921 2502 1166 2507
rect 1257 2507 1262 2512
rect 1433 2507 1702 2512
rect 2297 2507 2366 2512
rect 3313 2507 3318 2512
rect 1257 2502 1438 2507
rect 1697 2502 1950 2507
rect 2025 2502 2302 2507
rect 2361 2502 2454 2507
rect 1945 2497 2030 2502
rect 2449 2497 2454 2502
rect 2537 2502 2646 2507
rect 2705 2502 2958 2507
rect 3193 2502 3318 2507
rect 4657 2502 4734 2507
rect 2537 2497 2542 2502
rect 2641 2497 2710 2502
rect 2953 2497 3198 2502
rect 201 2492 246 2497
rect 1009 2492 1038 2497
rect 1033 2487 1038 2492
rect 1137 2492 1334 2497
rect 1449 2492 1686 2497
rect 2313 2492 2350 2497
rect 2449 2492 2542 2497
rect 2561 2492 2590 2497
rect 1137 2487 1142 2492
rect 1329 2487 1454 2492
rect 2585 2487 2590 2492
rect 2729 2492 2758 2497
rect 3481 2492 3654 2497
rect 3873 2492 3918 2497
rect 2729 2487 2734 2492
rect 225 2482 294 2487
rect 401 2482 542 2487
rect 1033 2482 1142 2487
rect 1289 2482 1310 2487
rect 1473 2482 1518 2487
rect 1777 2482 2430 2487
rect 2585 2482 2734 2487
rect 3025 2482 3422 2487
rect 3433 2482 3462 2487
rect 1545 2477 1758 2482
rect 3481 2477 3486 2492
rect 3649 2487 3654 2492
rect 3649 2482 3854 2487
rect 4689 2482 4726 2487
rect 3849 2477 3854 2482
rect 665 2472 998 2477
rect 993 2467 998 2472
rect 1161 2472 1246 2477
rect 1161 2467 1166 2472
rect 1241 2467 1246 2472
rect 1409 2472 1550 2477
rect 1753 2472 1822 2477
rect 2409 2472 2430 2477
rect 2921 2472 3006 2477
rect 3425 2472 3486 2477
rect 3505 2472 3630 2477
rect 3849 2472 3902 2477
rect 3937 2472 4166 2477
rect 1409 2467 1414 2472
rect 1841 2467 2214 2472
rect 2273 2467 2390 2472
rect 2921 2467 2926 2472
rect 3001 2467 3406 2472
rect 3505 2467 3510 2472
rect 993 2462 1166 2467
rect 1185 2462 1222 2467
rect 1241 2462 1414 2467
rect 1433 2462 1462 2467
rect 1457 2457 1462 2462
rect 1561 2462 1846 2467
rect 2209 2462 2238 2467
rect 2249 2462 2278 2467
rect 2385 2462 2510 2467
rect 2609 2462 2878 2467
rect 2897 2462 2926 2467
rect 3401 2462 3510 2467
rect 3625 2467 3630 2472
rect 3937 2467 3942 2472
rect 3625 2462 3942 2467
rect 4161 2467 4166 2472
rect 4161 2462 4342 2467
rect 1561 2457 1566 2462
rect 2609 2457 2614 2462
rect 393 2452 630 2457
rect 393 2447 398 2452
rect 265 2442 398 2447
rect 265 2437 270 2442
rect 225 2432 270 2437
rect 625 2437 630 2452
rect 673 2452 918 2457
rect 1457 2452 1566 2457
rect 1585 2452 1654 2457
rect 673 2447 678 2452
rect 649 2442 678 2447
rect 913 2447 918 2452
rect 1649 2447 1654 2452
rect 1753 2452 2614 2457
rect 2873 2457 2878 2462
rect 2873 2452 3654 2457
rect 3665 2452 3702 2457
rect 4601 2452 4646 2457
rect 1753 2447 1758 2452
rect 3649 2447 3654 2452
rect 3721 2447 3838 2452
rect 913 2442 950 2447
rect 1649 2442 1758 2447
rect 1817 2442 2278 2447
rect 2369 2442 2446 2447
rect 2649 2442 2766 2447
rect 2801 2442 3270 2447
rect 3649 2442 3726 2447
rect 3833 2442 4150 2447
rect 4473 2442 4646 2447
rect 4657 2442 4678 2447
rect 2273 2437 2374 2442
rect 2649 2437 2654 2442
rect 625 2432 902 2437
rect 1057 2432 1182 2437
rect 1321 2432 1406 2437
rect 1449 2432 1630 2437
rect 1777 2432 1814 2437
rect 1825 2432 2254 2437
rect 2393 2432 2494 2437
rect 2625 2432 2654 2437
rect 2761 2437 2766 2442
rect 3473 2437 3630 2442
rect 2761 2432 2790 2437
rect 2817 2432 2854 2437
rect 2985 2432 3374 2437
rect 3449 2432 3478 2437
rect 3625 2432 3822 2437
rect 4345 2432 4614 2437
rect 4665 2432 4718 2437
rect 2849 2427 2990 2432
rect 137 2422 182 2427
rect 409 2422 454 2427
rect 481 2422 518 2427
rect 609 2422 694 2427
rect 689 2417 694 2422
rect 801 2422 846 2427
rect 1161 2422 1214 2427
rect 1801 2422 1918 2427
rect 2041 2422 2094 2427
rect 2273 2422 2334 2427
rect 2401 2422 2446 2427
rect 2569 2422 2646 2427
rect 2681 2422 2726 2427
rect 2785 2422 2830 2427
rect 3009 2422 3110 2427
rect 3121 2422 3174 2427
rect 3289 2422 3318 2427
rect 3385 2422 3462 2427
rect 3473 2422 3782 2427
rect 801 2417 806 2422
rect 1913 2417 2046 2422
rect 3473 2417 3478 2422
rect 3777 2417 3782 2422
rect 3929 2422 4070 2427
rect 4129 2422 4174 2427
rect 4257 2422 4342 2427
rect 4521 2422 4574 2427
rect 4585 2422 4622 2427
rect 4673 2422 4774 2427
rect 3929 2417 3934 2422
rect 281 2412 334 2417
rect 361 2412 630 2417
rect 689 2412 806 2417
rect 921 2412 1038 2417
rect 1281 2412 1390 2417
rect 2065 2412 2558 2417
rect 2841 2412 2966 2417
rect 921 2407 926 2412
rect 177 2402 478 2407
rect 825 2402 926 2407
rect 1033 2407 1038 2412
rect 2553 2407 2846 2412
rect 2961 2407 2966 2412
rect 3217 2412 3374 2417
rect 3433 2412 3478 2417
rect 3505 2412 3590 2417
rect 3689 2412 3718 2417
rect 3777 2412 3934 2417
rect 4265 2412 4294 2417
rect 4353 2412 4382 2417
rect 3217 2407 3222 2412
rect 3369 2407 3438 2412
rect 1033 2402 1278 2407
rect 1401 2402 2022 2407
rect 2249 2402 2302 2407
rect 2401 2402 2462 2407
rect 2897 2402 2942 2407
rect 2961 2402 3222 2407
rect 3241 2402 3278 2407
rect 3457 2402 3550 2407
rect 3633 2402 3670 2407
rect 4025 2402 4094 2407
rect 4313 2402 4718 2407
rect 1273 2397 1406 2402
rect 2041 2397 2230 2402
rect 161 2392 190 2397
rect 273 2392 302 2397
rect 313 2392 534 2397
rect 593 2392 670 2397
rect 1961 2392 2046 2397
rect 2225 2392 2494 2397
rect 2513 2392 2822 2397
rect 2865 2392 2918 2397
rect 3249 2392 3302 2397
rect 3345 2392 3526 2397
rect 3641 2392 3726 2397
rect 3953 2392 4038 2397
rect 4065 2392 4254 2397
rect 185 2387 278 2392
rect 593 2387 598 2392
rect 1145 2387 1254 2392
rect 1833 2387 1942 2392
rect 2513 2387 2518 2392
rect 305 2382 342 2387
rect 441 2382 598 2387
rect 689 2382 782 2387
rect 801 2382 878 2387
rect 905 2382 1150 2387
rect 1249 2382 1278 2387
rect 1377 2382 1542 2387
rect 1609 2382 1646 2387
rect 1761 2382 1838 2387
rect 1937 2382 2070 2387
rect 2081 2382 2286 2387
rect 2297 2382 2518 2387
rect 2817 2387 2822 2392
rect 4249 2387 4254 2392
rect 4353 2392 4406 2397
rect 4577 2392 4598 2397
rect 4705 2392 4726 2397
rect 4353 2387 4358 2392
rect 2817 2382 2846 2387
rect 3617 2382 3646 2387
rect 3689 2382 3734 2387
rect 4249 2382 4358 2387
rect 4401 2387 4406 2392
rect 4401 2382 4470 2387
rect 4585 2382 4630 2387
rect 4689 2382 4758 2387
rect 689 2377 694 2382
rect 81 2372 150 2377
rect 145 2367 150 2372
rect 209 2372 366 2377
rect 505 2372 550 2377
rect 609 2372 694 2377
rect 777 2377 782 2382
rect 2537 2377 2798 2382
rect 777 2372 870 2377
rect 1161 2372 1262 2377
rect 1529 2372 1686 2377
rect 1785 2372 1870 2377
rect 1897 2372 1958 2377
rect 2257 2372 2542 2377
rect 2793 2372 2870 2377
rect 2937 2372 3150 2377
rect 209 2367 214 2372
rect 1953 2367 2262 2372
rect 145 2362 214 2367
rect 233 2362 398 2367
rect 609 2362 638 2367
rect 1121 2362 1390 2367
rect 1417 2362 1502 2367
rect 1521 2362 1830 2367
rect 1913 2362 1934 2367
rect 2281 2362 2790 2367
rect 2937 2362 2942 2372
rect 1417 2357 1422 2362
rect 657 2352 854 2357
rect 937 2352 982 2357
rect 1081 2352 1142 2357
rect 1153 2352 1214 2357
rect 1361 2352 1422 2357
rect 1497 2357 1502 2362
rect 2809 2357 2942 2362
rect 3145 2357 3150 2372
rect 3425 2372 3566 2377
rect 3425 2367 3430 2372
rect 3561 2367 3798 2372
rect 3265 2362 3430 2367
rect 3793 2362 3846 2367
rect 4441 2362 4510 2367
rect 4441 2357 4446 2362
rect 1497 2352 1742 2357
rect 1873 2352 1966 2357
rect 2017 2352 2294 2357
rect 2393 2352 2422 2357
rect 2513 2352 2558 2357
rect 2673 2352 2814 2357
rect 2961 2352 3126 2357
rect 3145 2352 3174 2357
rect 3441 2352 3494 2357
rect 3521 2352 3550 2357
rect 353 2347 430 2352
rect 2553 2347 2678 2352
rect 2961 2347 2966 2352
rect 329 2342 358 2347
rect 425 2342 630 2347
rect 673 2342 702 2347
rect 825 2342 854 2347
rect 1041 2342 1062 2347
rect 1129 2342 1174 2347
rect 1433 2342 1550 2347
rect 1745 2342 1982 2347
rect 2329 2342 2534 2347
rect 2697 2342 2966 2347
rect 3121 2347 3126 2352
rect 3545 2347 3550 2352
rect 3625 2352 3814 2357
rect 4233 2352 4446 2357
rect 4505 2357 4510 2362
rect 4505 2352 4598 2357
rect 3625 2347 3630 2352
rect 3121 2342 3222 2347
rect 3465 2342 3502 2347
rect 3545 2342 3630 2347
rect 4017 2342 4118 2347
rect 4433 2342 4494 2347
rect 4609 2342 4694 2347
rect 697 2337 830 2342
rect 2033 2337 2190 2342
rect 257 2332 414 2337
rect 929 2332 1478 2337
rect 1473 2327 1478 2332
rect 1561 2332 1734 2337
rect 1793 2332 2038 2337
rect 2185 2332 2318 2337
rect 2545 2332 2726 2337
rect 2865 2332 3326 2337
rect 3649 2332 3758 2337
rect 1561 2327 1566 2332
rect 1729 2327 1798 2332
rect 2313 2327 2550 2332
rect 2721 2327 2870 2332
rect 3649 2327 3654 2332
rect 393 2322 534 2327
rect 753 2322 910 2327
rect 1193 2322 1230 2327
rect 1385 2322 1454 2327
rect 1473 2322 1566 2327
rect 1817 2322 1942 2327
rect 2049 2322 2174 2327
rect 2649 2322 2702 2327
rect 2889 2322 2934 2327
rect 3057 2322 3110 2327
rect 3153 2322 3270 2327
rect 217 2317 326 2322
rect 657 2317 758 2322
rect 905 2317 910 2322
rect 3265 2317 3270 2322
rect 3337 2322 3654 2327
rect 3753 2327 3758 2332
rect 3833 2332 3918 2337
rect 4617 2332 4766 2337
rect 3833 2327 3838 2332
rect 3753 2322 3838 2327
rect 3913 2327 3918 2332
rect 3913 2322 3990 2327
rect 4161 2322 4222 2327
rect 4641 2322 4670 2327
rect 3337 2317 3342 2322
rect 161 2312 222 2317
rect 321 2312 350 2317
rect 441 2312 486 2317
rect 633 2312 662 2317
rect 905 2312 1014 2317
rect 1081 2312 1182 2317
rect 1249 2312 1366 2317
rect 1649 2312 3158 2317
rect 3201 2312 3246 2317
rect 3265 2312 3342 2317
rect 3393 2312 3446 2317
rect 3657 2312 3742 2317
rect 3889 2312 3966 2317
rect 4097 2312 4126 2317
rect 4233 2312 4310 2317
rect 4409 2312 4566 2317
rect 4601 2312 4638 2317
rect 1249 2307 1254 2312
rect 1361 2307 1526 2312
rect 4121 2307 4238 2312
rect 209 2302 286 2307
rect 281 2287 286 2302
rect 481 2302 510 2307
rect 561 2302 702 2307
rect 481 2287 486 2302
rect 697 2297 702 2302
rect 769 2302 1254 2307
rect 1521 2302 1550 2307
rect 1785 2302 1838 2307
rect 2025 2302 2070 2307
rect 2681 2302 2726 2307
rect 2945 2302 2998 2307
rect 3033 2302 3174 2307
rect 3465 2302 3518 2307
rect 3529 2302 3574 2307
rect 3825 2302 3950 2307
rect 3985 2302 4070 2307
rect 769 2297 774 2302
rect 1569 2297 1766 2302
rect 1857 2297 2006 2302
rect 2089 2297 2350 2302
rect 3985 2297 3990 2302
rect 697 2292 774 2297
rect 1001 2292 1030 2297
rect 1233 2292 1574 2297
rect 1761 2292 1862 2297
rect 2001 2292 2094 2297
rect 2345 2292 2670 2297
rect 2737 2292 2934 2297
rect 3041 2292 3118 2297
rect 3185 2292 3454 2297
rect 3529 2292 3646 2297
rect 1025 2287 1238 2292
rect 2665 2287 2742 2292
rect 2929 2287 3046 2292
rect 3113 2287 3190 2292
rect 3449 2287 3534 2292
rect 3641 2287 3646 2292
rect 3753 2292 3814 2297
rect 3913 2292 3990 2297
rect 4065 2297 4070 2302
rect 4065 2292 4086 2297
rect 3753 2287 3758 2292
rect 3809 2287 3918 2292
rect 4081 2287 4086 2292
rect 4153 2292 4286 2297
rect 4361 2292 4462 2297
rect 4153 2287 4158 2292
rect 281 2282 486 2287
rect 793 2282 822 2287
rect 897 2282 990 2287
rect 1497 2282 1526 2287
rect 1545 2282 2334 2287
rect 3065 2282 3094 2287
rect 3385 2282 3414 2287
rect 985 2277 990 2282
rect 1257 2277 1390 2282
rect 1497 2277 1502 2282
rect 3409 2277 3414 2282
rect 3553 2282 3582 2287
rect 3641 2282 3758 2287
rect 3937 2282 4030 2287
rect 4081 2282 4158 2287
rect 4177 2282 4254 2287
rect 3553 2277 3558 2282
rect 985 2272 1262 2277
rect 1385 2272 1502 2277
rect 1577 2272 1774 2277
rect 1937 2272 2998 2277
rect 3017 2272 3190 2277
rect 3209 2272 3310 2277
rect 3409 2272 3558 2277
rect 3889 2272 3982 2277
rect 1769 2267 1942 2272
rect 2993 2267 2998 2272
rect 1281 2262 1366 2267
rect 1721 2262 1750 2267
rect 1961 2262 2214 2267
rect 2993 2262 3054 2267
rect 4569 2262 4718 2267
rect 1585 2257 1702 2262
rect 2233 2257 2406 2262
rect 4569 2257 4574 2262
rect 225 2252 254 2257
rect 945 2252 1142 2257
rect 1161 2252 1590 2257
rect 1697 2252 2238 2257
rect 2401 2252 3278 2257
rect 4001 2252 4246 2257
rect 4505 2252 4574 2257
rect 4713 2257 4718 2262
rect 4713 2252 4742 2257
rect 289 2242 462 2247
rect 481 2242 598 2247
rect 889 2242 926 2247
rect 481 2237 486 2242
rect 177 2232 246 2237
rect 457 2232 486 2237
rect 593 2237 598 2242
rect 945 2237 950 2252
rect 1137 2242 1142 2252
rect 4001 2247 4006 2252
rect 1289 2242 1310 2247
rect 1601 2242 1694 2247
rect 1929 2242 2110 2247
rect 2161 2242 2326 2247
rect 2353 2242 2390 2247
rect 3417 2242 3486 2247
rect 3593 2242 3638 2247
rect 3657 2242 3878 2247
rect 3897 2242 3926 2247
rect 3961 2242 4006 2247
rect 4241 2247 4246 2252
rect 4241 2242 4382 2247
rect 1137 2237 1230 2242
rect 1329 2237 1526 2242
rect 3025 2237 3190 2242
rect 3657 2237 3662 2242
rect 593 2232 622 2237
rect 801 2232 830 2237
rect 897 2232 950 2237
rect 1225 2232 1334 2237
rect 1521 2232 1830 2237
rect 2025 2232 2118 2237
rect 2249 2232 2374 2237
rect 1825 2227 1830 2232
rect 1945 2227 2030 2232
rect 2113 2227 2254 2232
rect 2369 2227 2374 2232
rect 2601 2232 3030 2237
rect 3185 2232 3214 2237
rect 2601 2227 2606 2232
rect 3209 2227 3214 2232
rect 3289 2232 3662 2237
rect 3873 2237 3878 2242
rect 3873 2232 4142 2237
rect 3289 2227 3294 2232
rect 4137 2227 4142 2232
rect 4201 2232 4230 2237
rect 4585 2232 4614 2237
rect 4665 2232 4734 2237
rect 4201 2227 4206 2232
rect 129 2222 174 2227
rect 201 2222 246 2227
rect 417 2222 494 2227
rect 553 2222 598 2227
rect 689 2222 1046 2227
rect 1153 2222 1214 2227
rect 1321 2222 1438 2227
rect 1481 2222 1510 2227
rect 1505 2217 1510 2222
rect 1649 2222 1710 2227
rect 1777 2222 1806 2227
rect 1825 2222 1950 2227
rect 2049 2222 2094 2227
rect 2273 2222 2350 2227
rect 2369 2222 2606 2227
rect 3041 2222 3070 2227
rect 1649 2217 1654 2222
rect 3065 2217 3070 2222
rect 3129 2222 3190 2227
rect 3209 2222 3294 2227
rect 3457 2222 3526 2227
rect 3537 2222 3590 2227
rect 3681 2222 3854 2227
rect 3921 2222 4030 2227
rect 4137 2222 4206 2227
rect 4393 2222 4574 2227
rect 4601 2222 4702 2227
rect 3129 2217 3134 2222
rect 3681 2217 3686 2222
rect 393 2212 454 2217
rect 481 2212 574 2217
rect 641 2212 758 2217
rect 913 2212 942 2217
rect 1201 2212 1230 2217
rect 1505 2212 1654 2217
rect 1969 2212 2006 2217
rect 2113 2212 2182 2217
rect 2625 2212 2790 2217
rect 2865 2212 2894 2217
rect 3065 2212 3134 2217
rect 3417 2212 3686 2217
rect 3849 2217 3854 2222
rect 3849 2212 3958 2217
rect 4337 2212 4358 2217
rect 913 2202 918 2212
rect 2113 2207 2118 2212
rect 4377 2207 4518 2212
rect 1065 2202 1110 2207
rect 1145 2202 1198 2207
rect 2081 2202 2118 2207
rect 2233 2202 2342 2207
rect 2921 2202 2982 2207
rect 3153 2202 3182 2207
rect 3345 2202 3502 2207
rect 3529 2202 3558 2207
rect 3569 2202 3806 2207
rect 3865 2202 3966 2207
rect 4025 2202 4118 2207
rect 4305 2202 4382 2207
rect 4513 2202 4598 2207
rect 4641 2202 4670 2207
rect 2233 2197 2238 2202
rect 217 2192 294 2197
rect 617 2192 646 2197
rect 689 2192 798 2197
rect 857 2192 1030 2197
rect 1065 2192 1214 2197
rect 1401 2192 1582 2197
rect 1681 2192 1782 2197
rect 1809 2192 1846 2197
rect 1977 2192 2070 2197
rect 2209 2192 2238 2197
rect 2337 2197 2342 2202
rect 3569 2197 3574 2202
rect 2337 2192 2462 2197
rect 2881 2192 3014 2197
rect 3049 2192 3350 2197
rect 2065 2187 2150 2192
rect 3345 2187 3350 2192
rect 3449 2192 3478 2197
rect 3489 2192 3574 2197
rect 3649 2192 3734 2197
rect 3873 2192 3918 2197
rect 3937 2192 3942 2202
rect 4225 2192 4294 2197
rect 4369 2192 4398 2197
rect 4417 2192 4502 2197
rect 3449 2187 3454 2192
rect 4289 2187 4374 2192
rect 185 2182 214 2187
rect 777 2182 862 2187
rect 1041 2182 1070 2187
rect 1065 2177 1070 2182
rect 1177 2182 1334 2187
rect 1865 2182 1958 2187
rect 2145 2182 2422 2187
rect 2537 2182 2694 2187
rect 3345 2182 3454 2187
rect 3545 2182 3990 2187
rect 4417 2182 4718 2187
rect 1177 2177 1182 2182
rect 1561 2177 1694 2182
rect 1865 2177 1870 2182
rect 1065 2172 1182 2177
rect 1201 2172 1278 2177
rect 1433 2172 1566 2177
rect 1689 2172 1870 2177
rect 1953 2177 1958 2182
rect 2537 2177 2542 2182
rect 1953 2172 2494 2177
rect 2513 2172 2542 2177
rect 2689 2177 2694 2182
rect 2689 2172 2902 2177
rect 2969 2172 3086 2177
rect 3689 2172 3726 2177
rect 3801 2172 4438 2177
rect 513 2162 550 2167
rect 593 2162 614 2167
rect 1281 2162 1382 2167
rect 1577 2162 1678 2167
rect 2161 2162 2366 2167
rect 2561 2162 2662 2167
rect 2841 2162 2958 2167
rect 3081 2162 3326 2167
rect 3497 2162 3590 2167
rect 3825 2162 3854 2167
rect 3897 2162 3998 2167
rect 4697 2162 4758 2167
rect 2393 2157 2566 2162
rect 2657 2157 2662 2162
rect 2953 2157 3086 2162
rect 3497 2157 3502 2162
rect 505 2152 558 2157
rect 633 2152 678 2157
rect 945 2152 982 2157
rect 1041 2152 1182 2157
rect 1209 2152 1278 2157
rect 1729 2152 1758 2157
rect 449 2142 678 2147
rect 849 2142 950 2147
rect 1041 2137 1046 2152
rect 529 2127 534 2137
rect 737 2132 838 2137
rect 961 2132 1046 2137
rect 1177 2137 1182 2152
rect 1753 2147 1758 2152
rect 1873 2152 2398 2157
rect 2657 2152 2758 2157
rect 3105 2152 3134 2157
rect 3345 2152 3454 2157
rect 3473 2152 3502 2157
rect 3585 2157 3590 2162
rect 4409 2157 4494 2162
rect 3585 2152 3814 2157
rect 1873 2147 1878 2152
rect 2753 2147 2758 2152
rect 3217 2147 3350 2152
rect 3449 2147 3454 2152
rect 3809 2147 3814 2152
rect 3897 2152 3926 2157
rect 4089 2152 4198 2157
rect 4385 2152 4414 2157
rect 4489 2152 4654 2157
rect 3897 2147 3902 2152
rect 4089 2147 4094 2152
rect 1257 2142 1286 2147
rect 1393 2142 1598 2147
rect 1393 2137 1398 2142
rect 1177 2132 1398 2137
rect 1593 2137 1598 2142
rect 1697 2142 1726 2147
rect 1753 2142 1878 2147
rect 2057 2142 2086 2147
rect 2409 2142 2662 2147
rect 2753 2142 3222 2147
rect 3449 2142 3550 2147
rect 3561 2142 3598 2147
rect 3809 2142 3902 2147
rect 4001 2142 4038 2147
rect 4065 2142 4094 2147
rect 4193 2147 4198 2152
rect 4193 2142 4262 2147
rect 4441 2142 4478 2147
rect 4585 2142 4630 2147
rect 1697 2137 1702 2142
rect 2081 2137 2414 2142
rect 1593 2132 1702 2137
rect 1897 2132 1942 2137
rect 2433 2132 2510 2137
rect 2617 2132 2678 2137
rect 2713 2132 2742 2137
rect 833 2127 966 2132
rect 2737 2127 2742 2132
rect 2865 2132 2910 2137
rect 2993 2132 3062 2137
rect 3233 2132 3302 2137
rect 3321 2132 3366 2137
rect 3617 2132 3702 2137
rect 4057 2132 4182 2137
rect 4673 2132 4726 2137
rect 2865 2127 2870 2132
rect 3113 2127 3190 2132
rect 3617 2127 3622 2132
rect 249 2122 294 2127
rect 529 2122 574 2127
rect 609 2122 734 2127
rect 1057 2122 1238 2127
rect 1945 2122 2062 2127
rect 2145 2122 2582 2127
rect 2737 2122 2870 2127
rect 2889 2122 3118 2127
rect 3185 2122 3222 2127
rect 3313 2122 3342 2127
rect 3369 2122 3622 2127
rect 3697 2127 3702 2132
rect 3697 2122 3886 2127
rect 3217 2117 3318 2122
rect 425 2112 550 2117
rect 753 2112 830 2117
rect 569 2107 758 2112
rect 825 2107 830 2112
rect 945 2112 1038 2117
rect 945 2107 950 2112
rect 433 2102 574 2107
rect 825 2102 950 2107
rect 1033 2107 1038 2112
rect 1441 2112 1574 2117
rect 1921 2112 2046 2117
rect 2361 2112 2390 2117
rect 2465 2112 2510 2117
rect 2561 2112 2646 2117
rect 2969 2112 2990 2117
rect 3001 2112 3038 2117
rect 3129 2112 3174 2117
rect 3577 2112 3686 2117
rect 4057 2112 4254 2117
rect 4329 2112 4366 2117
rect 4457 2112 4542 2117
rect 1033 2102 1102 2107
rect 1121 2102 1366 2107
rect 1385 2102 1422 2107
rect 1121 2097 1126 2102
rect 441 2092 814 2097
rect 809 2087 814 2092
rect 961 2092 1126 2097
rect 1361 2097 1366 2102
rect 1441 2097 1446 2112
rect 1361 2092 1446 2097
rect 1569 2097 1574 2112
rect 1681 2102 1838 2107
rect 1929 2102 2350 2107
rect 2657 2102 2774 2107
rect 3001 2102 3030 2107
rect 3225 2102 3262 2107
rect 4041 2102 4070 2107
rect 1681 2097 1686 2102
rect 1569 2092 1686 2097
rect 1833 2097 1838 2102
rect 2345 2097 2454 2102
rect 2545 2097 2662 2102
rect 1833 2092 1862 2097
rect 2049 2092 2078 2097
rect 2161 2092 2190 2097
rect 2449 2092 2550 2097
rect 3049 2092 3206 2097
rect 961 2087 966 2092
rect 2073 2087 2166 2092
rect 3049 2087 3054 2092
rect 361 2082 430 2087
rect 761 2082 790 2087
rect 809 2082 966 2087
rect 985 2082 1110 2087
rect 1129 2082 1558 2087
rect 1721 2082 1814 2087
rect 425 2077 430 2082
rect 649 2077 766 2082
rect 1105 2077 1110 2082
rect 1721 2077 1726 2082
rect 425 2072 654 2077
rect 1105 2072 1134 2077
rect 1281 2072 1310 2077
rect 1577 2072 1678 2077
rect 1697 2072 1726 2077
rect 1809 2077 1814 2082
rect 1881 2082 2030 2087
rect 2569 2082 2638 2087
rect 2657 2082 2934 2087
rect 2953 2082 3054 2087
rect 3201 2087 3206 2092
rect 3281 2092 3350 2097
rect 3281 2087 3286 2092
rect 3201 2082 3286 2087
rect 3345 2087 3350 2092
rect 3393 2092 3510 2097
rect 3393 2087 3398 2092
rect 3345 2082 3398 2087
rect 3505 2087 3510 2092
rect 4065 2087 4070 2102
rect 4353 2102 4382 2107
rect 4353 2087 4358 2102
rect 3505 2082 3534 2087
rect 3945 2082 3982 2087
rect 4065 2082 4358 2087
rect 1881 2077 1886 2082
rect 1809 2072 1886 2077
rect 2025 2077 2030 2082
rect 2657 2077 2662 2082
rect 2025 2072 2662 2077
rect 2929 2077 2934 2082
rect 3073 2077 3182 2082
rect 2929 2072 3078 2077
rect 3177 2072 3222 2077
rect 4025 2072 4046 2077
rect 1129 2067 1286 2072
rect 1417 2067 1582 2072
rect 1673 2067 1678 2072
rect 3241 2067 3518 2072
rect 241 2062 342 2067
rect 241 2057 246 2062
rect 217 2052 246 2057
rect 337 2057 342 2062
rect 673 2062 1086 2067
rect 1393 2062 1422 2067
rect 1673 2062 2030 2067
rect 2217 2062 2246 2067
rect 2505 2062 3246 2067
rect 3513 2062 3654 2067
rect 673 2057 678 2062
rect 337 2052 678 2057
rect 1081 2057 1086 2062
rect 2025 2057 2222 2062
rect 1081 2052 1734 2057
rect 2593 2052 2662 2057
rect 2961 2052 3502 2057
rect 3681 2052 3838 2057
rect 833 2047 942 2052
rect 1793 2047 2006 2052
rect 2465 2047 2574 2052
rect 689 2042 838 2047
rect 937 2042 1078 2047
rect 1345 2042 1798 2047
rect 2001 2042 2470 2047
rect 2569 2042 2950 2047
rect 3025 2042 3286 2047
rect 1073 2037 1078 2042
rect 1233 2037 1350 2042
rect 2945 2037 3030 2042
rect 3313 2037 3430 2042
rect 3681 2037 3686 2052
rect 177 2032 374 2037
rect 521 2032 1054 2037
rect 1073 2032 1238 2037
rect 1369 2032 1462 2037
rect 1545 2032 1630 2037
rect 1809 2032 1990 2037
rect 2481 2032 2694 2037
rect 3289 2032 3318 2037
rect 3425 2032 3454 2037
rect 3513 2032 3534 2037
rect 3657 2032 3686 2037
rect 3833 2037 3838 2052
rect 3881 2052 3950 2057
rect 4153 2052 4214 2057
rect 3881 2047 3886 2052
rect 3857 2042 3886 2047
rect 3945 2047 3950 2052
rect 3945 2042 4038 2047
rect 3833 2032 3918 2037
rect 4601 2032 4694 2037
rect 1457 2027 1550 2032
rect 1625 2027 1814 2032
rect 2121 2027 2310 2032
rect 3049 2027 3270 2032
rect 65 2022 142 2027
rect 161 2022 454 2027
rect 537 2022 982 2027
rect 993 2022 1014 2027
rect 1257 2022 1438 2027
rect 1569 2022 1606 2027
rect 1833 2022 1926 2027
rect 2025 2022 2126 2027
rect 2305 2022 2398 2027
rect 2465 2022 2606 2027
rect 2649 2022 2750 2027
rect 2897 2022 2958 2027
rect 2969 2022 3054 2027
rect 3265 2022 3350 2027
rect 3401 2022 3582 2027
rect 3665 2022 3750 2027
rect 3873 2022 3934 2027
rect 4033 2022 4070 2027
rect 4281 2022 4374 2027
rect 4625 2022 4750 2027
rect 65 2017 70 2022
rect 0 2012 70 2017
rect 137 2017 142 2022
rect 137 2012 222 2017
rect 233 2012 278 2017
rect 321 2012 382 2017
rect 489 2012 518 2017
rect 561 2012 614 2017
rect 705 2012 878 2017
rect 377 2007 494 2012
rect 609 2007 710 2012
rect 873 2007 878 2012
rect 1025 2012 1246 2017
rect 1449 2012 1558 2017
rect 1617 2012 1822 2017
rect 1025 2007 1030 2012
rect 1241 2007 1454 2012
rect 1553 2007 1622 2012
rect 1817 2007 1822 2012
rect 1913 2012 1942 2017
rect 1985 2012 2014 2017
rect 2137 2012 2366 2017
rect 2569 2012 2598 2017
rect 2769 2012 2878 2017
rect 2937 2012 2982 2017
rect 3065 2012 3470 2017
rect 3593 2012 3622 2017
rect 3657 2012 3694 2017
rect 3905 2012 4070 2017
rect 1913 2007 1918 2012
rect 2009 2007 2142 2012
rect 2361 2007 2454 2012
rect 2569 2007 2574 2012
rect 2769 2007 2774 2012
rect 209 2002 310 2007
rect 553 2002 590 2007
rect 729 2002 838 2007
rect 873 2002 1030 2007
rect 1817 2002 1918 2007
rect 2449 2002 2574 2007
rect 2729 2002 2774 2007
rect 2873 2007 2878 2012
rect 3465 2007 3598 2012
rect 3729 2007 3870 2012
rect 2873 2002 2902 2007
rect 2993 2002 3334 2007
rect 3649 2002 3670 2007
rect 3705 2002 3734 2007
rect 3865 2002 4078 2007
rect 2161 1997 2342 2002
rect 2897 1997 2998 2002
rect 3329 1997 3334 2002
rect 81 1992 190 1997
rect 241 1992 462 1997
rect 545 1992 718 1997
rect 825 1992 854 1997
rect 1297 1992 1414 1997
rect 1585 1992 1622 1997
rect 2049 1992 2166 1997
rect 2337 1992 2366 1997
rect 2617 1992 2710 1997
rect 3025 1992 3110 1997
rect 3137 1992 3310 1997
rect 3329 1992 3358 1997
rect 713 1987 830 1992
rect 1297 1987 1302 1992
rect 97 1982 174 1987
rect 273 1982 342 1987
rect 873 1982 1254 1987
rect 1273 1982 1302 1987
rect 1409 1987 1414 1992
rect 2617 1987 2622 1992
rect 2705 1987 2862 1992
rect 3353 1987 3358 1992
rect 3513 1992 3542 1997
rect 3617 1992 3646 1997
rect 3513 1987 3518 1992
rect 1409 1982 1438 1987
rect 1457 1982 1566 1987
rect 873 1977 878 1982
rect 281 1972 422 1977
rect 577 1972 622 1977
rect 617 1967 622 1972
rect 761 1972 878 1977
rect 1249 1977 1254 1982
rect 1457 1977 1462 1982
rect 1249 1972 1462 1977
rect 1561 1977 1566 1982
rect 1705 1982 2030 1987
rect 2177 1982 2486 1987
rect 2545 1982 2622 1987
rect 2857 1982 2974 1987
rect 3105 1982 3326 1987
rect 3353 1982 3518 1987
rect 1705 1977 1710 1982
rect 1561 1972 1606 1977
rect 1649 1972 1710 1977
rect 2025 1977 2030 1982
rect 3641 1977 3646 1992
rect 3761 1992 3854 1997
rect 3921 1992 3950 1997
rect 3761 1977 3766 1992
rect 3945 1987 3950 1992
rect 4025 1992 4054 1997
rect 4065 1992 4166 1997
rect 4209 1992 4238 1997
rect 4361 1992 4398 1997
rect 4025 1987 4030 1992
rect 3945 1982 4030 1987
rect 2025 1972 2846 1977
rect 761 1967 766 1972
rect 2841 1967 2846 1972
rect 2945 1972 3046 1977
rect 3145 1972 3174 1977
rect 2945 1967 2950 1972
rect 3169 1967 3174 1972
rect 3289 1972 3318 1977
rect 3641 1972 3766 1977
rect 3833 1972 3910 1977
rect 3289 1967 3294 1972
rect 3833 1967 3838 1972
rect 337 1962 358 1967
rect 617 1962 766 1967
rect 833 1962 1342 1967
rect 1337 1957 1342 1962
rect 1473 1962 1598 1967
rect 1745 1962 1830 1967
rect 1897 1962 2046 1967
rect 2241 1962 2822 1967
rect 2841 1962 2950 1967
rect 2969 1962 3054 1967
rect 3169 1962 3294 1967
rect 3809 1962 3838 1967
rect 3905 1967 3910 1972
rect 3905 1962 3934 1967
rect 3953 1962 4038 1967
rect 1473 1957 1478 1962
rect 1745 1957 1750 1962
rect 497 1952 598 1957
rect 1337 1952 1478 1957
rect 1721 1952 1750 1957
rect 1825 1957 1830 1962
rect 3953 1957 3958 1962
rect 1825 1952 1982 1957
rect 2209 1952 2270 1957
rect 3785 1952 3958 1957
rect 4033 1957 4038 1962
rect 4033 1952 4062 1957
rect 977 1947 1294 1952
rect 1521 1947 1702 1952
rect 2289 1947 2782 1952
rect 121 1942 270 1947
rect 377 1942 478 1947
rect 785 1942 982 1947
rect 1289 1942 1318 1947
rect 1497 1942 1526 1947
rect 1697 1942 1814 1947
rect 2009 1942 2054 1947
rect 2073 1942 2166 1947
rect 2185 1942 2294 1947
rect 2777 1942 2926 1947
rect 2945 1942 3278 1947
rect 3697 1942 3726 1947
rect 3777 1942 3806 1947
rect 3817 1942 3966 1947
rect 4025 1942 4326 1947
rect 4385 1942 4510 1947
rect 377 1937 382 1942
rect 137 1932 166 1937
rect 161 1927 166 1932
rect 281 1932 382 1937
rect 473 1937 478 1942
rect 1313 1937 1318 1942
rect 1833 1937 1902 1942
rect 2073 1937 2078 1942
rect 473 1932 582 1937
rect 721 1932 750 1937
rect 993 1932 1270 1937
rect 1313 1932 1838 1937
rect 1897 1932 2078 1937
rect 2161 1937 2166 1942
rect 2945 1937 2950 1942
rect 2161 1932 2766 1937
rect 2921 1932 2950 1937
rect 3593 1932 3654 1937
rect 3745 1932 3798 1937
rect 3833 1932 3878 1937
rect 281 1927 286 1932
rect 745 1927 998 1932
rect 2761 1927 2926 1932
rect 161 1922 286 1927
rect 1673 1922 1886 1927
rect 1993 1922 2206 1927
rect 2361 1922 2526 1927
rect 2569 1922 2742 1927
rect 3009 1922 3198 1927
rect 3305 1922 3478 1927
rect 3497 1922 3590 1927
rect 1017 1917 1590 1922
rect 2201 1917 2366 1922
rect 3473 1917 3478 1922
rect 361 1912 406 1917
rect 457 1912 518 1917
rect 577 1912 646 1917
rect 689 1912 1022 1917
rect 1585 1912 1726 1917
rect 1801 1912 1846 1917
rect 1945 1912 2054 1917
rect 2385 1912 2470 1917
rect 2481 1912 2734 1917
rect 2817 1912 2998 1917
rect 3201 1912 3318 1917
rect 3473 1912 3718 1917
rect 4121 1912 4174 1917
rect 4505 1912 4534 1917
rect 2073 1907 2182 1912
rect 353 1902 406 1907
rect 529 1902 558 1907
rect 553 1897 558 1902
rect 641 1902 670 1907
rect 1033 1902 1574 1907
rect 1737 1902 2078 1907
rect 2177 1902 2374 1907
rect 2457 1902 2806 1907
rect 3009 1902 3126 1907
rect 3209 1902 3238 1907
rect 641 1897 646 1902
rect 1569 1897 1742 1902
rect 2369 1897 2462 1902
rect 2801 1897 3014 1902
rect 3233 1897 3238 1902
rect 3305 1902 3598 1907
rect 3305 1897 3310 1902
rect 3593 1897 3598 1902
rect 3729 1902 3798 1907
rect 3729 1897 3734 1902
rect 265 1892 342 1897
rect 441 1892 470 1897
rect 553 1892 646 1897
rect 721 1892 1326 1897
rect 1521 1892 1550 1897
rect 1825 1892 2166 1897
rect 3081 1892 3150 1897
rect 3233 1892 3310 1897
rect 3329 1892 3358 1897
rect 337 1887 446 1892
rect 1377 1887 1502 1892
rect 2481 1887 2742 1892
rect 3353 1887 3358 1892
rect 3497 1892 3526 1897
rect 3545 1892 3574 1897
rect 3593 1892 3734 1897
rect 3809 1892 4110 1897
rect 3497 1887 3502 1892
rect 721 1882 742 1887
rect 985 1882 1014 1887
rect 1009 1877 1014 1882
rect 1097 1882 1150 1887
rect 1337 1882 1382 1887
rect 1497 1882 1814 1887
rect 2089 1882 2486 1887
rect 2737 1882 3134 1887
rect 3353 1882 3502 1887
rect 1097 1877 1102 1882
rect 1145 1877 1342 1882
rect 1809 1877 2094 1882
rect 3569 1877 3574 1892
rect 3809 1877 3814 1892
rect 4105 1887 4110 1892
rect 4185 1892 4742 1897
rect 4185 1887 4190 1892
rect 4105 1882 4190 1887
rect 393 1872 566 1877
rect 585 1872 846 1877
rect 1009 1872 1102 1877
rect 1393 1872 1558 1877
rect 2497 1872 2726 1877
rect 3033 1872 3078 1877
rect 3569 1872 3814 1877
rect 841 1867 846 1872
rect 1393 1867 1398 1872
rect 1577 1867 1774 1872
rect 2113 1867 2270 1872
rect 2313 1867 2502 1872
rect 841 1862 974 1867
rect 969 1857 974 1862
rect 1121 1862 1398 1867
rect 1457 1862 1582 1867
rect 1769 1862 2118 1867
rect 2265 1862 2318 1867
rect 2521 1862 2878 1867
rect 1121 1857 1126 1862
rect 433 1852 462 1857
rect 785 1852 822 1857
rect 969 1852 1126 1857
rect 1417 1852 1758 1857
rect 2129 1852 2550 1857
rect 2585 1852 2614 1857
rect 2897 1852 3014 1857
rect 3433 1852 3526 1857
rect 1753 1847 1846 1852
rect 2129 1847 2134 1852
rect 2633 1847 2902 1852
rect 3009 1847 3014 1852
rect 745 1842 782 1847
rect 1169 1842 1294 1847
rect 1337 1842 1734 1847
rect 1841 1842 2134 1847
rect 2257 1842 2446 1847
rect 2529 1842 2638 1847
rect 3009 1842 3422 1847
rect 2441 1837 2534 1842
rect 3417 1837 3422 1842
rect 3537 1842 3750 1847
rect 4521 1842 4598 1847
rect 3537 1837 3542 1842
rect 1145 1832 1198 1837
rect 1441 1832 1822 1837
rect 2377 1832 2422 1837
rect 2553 1832 3006 1837
rect 3417 1832 3542 1837
rect 3713 1832 3814 1837
rect 4209 1832 4246 1837
rect 4617 1832 4646 1837
rect 201 1822 246 1827
rect 449 1822 526 1827
rect 649 1822 1430 1827
rect 1425 1817 1430 1822
rect 1601 1822 1702 1827
rect 1713 1822 1742 1827
rect 1857 1822 1902 1827
rect 1945 1822 1974 1827
rect 2049 1822 2134 1827
rect 2233 1822 2366 1827
rect 1601 1817 1606 1822
rect 249 1812 294 1817
rect 305 1812 382 1817
rect 1425 1812 1606 1817
rect 1697 1817 1702 1822
rect 2361 1817 2366 1822
rect 2433 1822 2638 1827
rect 2433 1817 2438 1822
rect 2633 1817 2638 1822
rect 2705 1822 2734 1827
rect 2857 1822 2902 1827
rect 2969 1822 3070 1827
rect 3745 1822 3798 1827
rect 3825 1822 3894 1827
rect 3929 1822 4006 1827
rect 4073 1822 4182 1827
rect 4225 1822 4262 1827
rect 4345 1822 4438 1827
rect 4457 1822 4630 1827
rect 4681 1822 4718 1827
rect 4761 1822 4790 1827
rect 2705 1817 2710 1822
rect 3929 1817 3934 1822
rect 1697 1812 1886 1817
rect 1985 1812 2062 1817
rect 2361 1812 2438 1817
rect 2529 1812 2566 1817
rect 2633 1812 2710 1817
rect 3153 1812 3262 1817
rect 3873 1812 3934 1817
rect 4001 1817 4006 1822
rect 4345 1817 4350 1822
rect 4001 1812 4030 1817
rect 4321 1812 4350 1817
rect 4433 1817 4438 1822
rect 4433 1812 4614 1817
rect 289 1807 294 1812
rect 1153 1807 1358 1812
rect 1881 1807 1990 1812
rect 2121 1807 2238 1812
rect 3753 1807 3846 1812
rect 233 1802 262 1807
rect 289 1802 542 1807
rect 673 1802 726 1807
rect 977 1802 1110 1807
rect 1129 1802 1158 1807
rect 1353 1802 1382 1807
rect 977 1797 982 1802
rect 81 1792 158 1797
rect 241 1792 366 1797
rect 593 1792 670 1797
rect 793 1792 814 1797
rect 833 1792 934 1797
rect 953 1792 982 1797
rect 1105 1797 1110 1802
rect 1377 1797 1382 1802
rect 1625 1802 1654 1807
rect 1785 1802 1862 1807
rect 1625 1797 1630 1802
rect 1857 1797 1862 1802
rect 2097 1802 2126 1807
rect 2233 1802 2262 1807
rect 2273 1802 2302 1807
rect 2569 1802 2614 1807
rect 2753 1802 2886 1807
rect 3585 1802 3758 1807
rect 3841 1802 3902 1807
rect 4049 1802 4118 1807
rect 4177 1802 4646 1807
rect 2097 1797 2102 1802
rect 4049 1797 4054 1802
rect 1105 1792 1174 1797
rect 1185 1792 1358 1797
rect 1377 1792 1630 1797
rect 1777 1792 1838 1797
rect 1857 1792 2102 1797
rect 2121 1792 2470 1797
rect 3385 1792 3502 1797
rect 3769 1792 3830 1797
rect 3945 1792 4054 1797
rect 4113 1797 4118 1802
rect 4641 1797 4646 1802
rect 4113 1792 4198 1797
rect 4457 1792 4566 1797
rect 4641 1792 4686 1797
rect 361 1787 366 1792
rect 441 1787 582 1792
rect 833 1787 838 1792
rect 129 1782 262 1787
rect 361 1782 446 1787
rect 577 1782 838 1787
rect 929 1787 934 1792
rect 929 1782 1350 1787
rect 2193 1782 2286 1787
rect 2905 1782 2974 1787
rect 3785 1782 4270 1787
rect 4425 1782 4686 1787
rect 2905 1777 2910 1782
rect 257 1772 334 1777
rect 465 1772 494 1777
rect 489 1767 494 1772
rect 617 1772 1022 1777
rect 1281 1772 1310 1777
rect 1769 1772 1886 1777
rect 2129 1772 2262 1777
rect 2625 1772 2670 1777
rect 2809 1772 2910 1777
rect 2969 1777 2974 1782
rect 2969 1772 3038 1777
rect 3337 1772 3398 1777
rect 3753 1772 3950 1777
rect 4049 1772 4078 1777
rect 4097 1772 4134 1777
rect 4313 1772 4406 1777
rect 4625 1772 4734 1777
rect 617 1767 622 1772
rect 1057 1767 1206 1772
rect 1769 1767 1774 1772
rect 489 1762 622 1767
rect 641 1762 934 1767
rect 929 1757 934 1762
rect 1033 1762 1062 1767
rect 1201 1762 1462 1767
rect 1497 1762 1710 1767
rect 1745 1762 1774 1767
rect 1881 1767 1886 1772
rect 4313 1767 4318 1772
rect 4401 1767 4606 1772
rect 1881 1762 1910 1767
rect 2065 1762 2406 1767
rect 3417 1762 3582 1767
rect 3777 1762 4318 1767
rect 4601 1762 4702 1767
rect 1033 1757 1038 1762
rect 649 1752 894 1757
rect 929 1752 1038 1757
rect 1081 1752 1246 1757
rect 1265 1752 1326 1757
rect 1497 1747 1502 1762
rect 1705 1747 1710 1762
rect 3417 1757 3422 1762
rect 1729 1752 1974 1757
rect 2145 1752 2510 1757
rect 2865 1752 3206 1757
rect 3257 1752 3422 1757
rect 3577 1757 3582 1762
rect 3577 1752 3606 1757
rect 3737 1752 4134 1757
rect 4329 1752 4606 1757
rect 209 1742 278 1747
rect 353 1742 414 1747
rect 705 1742 830 1747
rect 873 1742 910 1747
rect 1105 1742 1174 1747
rect 1193 1742 1262 1747
rect 1393 1742 1422 1747
rect 1433 1742 1502 1747
rect 1561 1742 1638 1747
rect 1705 1742 1750 1747
rect 1817 1742 2014 1747
rect 2025 1742 2254 1747
rect 2281 1742 2374 1747
rect 2625 1742 2742 1747
rect 3401 1742 3542 1747
rect 3625 1742 3670 1747
rect 3785 1742 4166 1747
rect 4393 1742 4502 1747
rect 1561 1737 1566 1742
rect 201 1732 334 1737
rect 449 1732 478 1737
rect 521 1732 622 1737
rect 329 1727 454 1732
rect 521 1727 526 1732
rect 233 1722 262 1727
rect 273 1722 310 1727
rect 481 1722 526 1727
rect 617 1727 622 1732
rect 617 1722 646 1727
rect 321 1712 366 1717
rect 553 1712 582 1717
rect 657 1712 662 1737
rect 769 1732 790 1737
rect 881 1732 950 1737
rect 1073 1732 1102 1737
rect 1177 1732 1222 1737
rect 1329 1732 1382 1737
rect 945 1727 950 1732
rect 1377 1727 1382 1732
rect 1449 1732 1566 1737
rect 1633 1737 1638 1742
rect 1633 1732 2150 1737
rect 1449 1727 1454 1732
rect 2225 1727 2230 1742
rect 2625 1737 2630 1742
rect 2265 1732 2294 1737
rect 2433 1727 2438 1737
rect 2601 1732 2630 1737
rect 2737 1737 2742 1742
rect 2849 1737 2942 1742
rect 3049 1737 3230 1742
rect 3265 1737 3382 1742
rect 3537 1737 3630 1742
rect 4497 1737 4502 1742
rect 4617 1742 4678 1747
rect 4617 1737 4622 1742
rect 2737 1732 2854 1737
rect 2937 1732 3054 1737
rect 3225 1732 3270 1737
rect 3377 1732 3486 1737
rect 3649 1732 3750 1737
rect 3865 1732 3966 1737
rect 4001 1732 4046 1737
rect 4153 1732 4206 1737
rect 4497 1732 4622 1737
rect 4001 1727 4006 1732
rect 745 1722 862 1727
rect 945 1722 966 1727
rect 1033 1722 1206 1727
rect 1377 1722 1454 1727
rect 1473 1722 1494 1727
rect 1577 1722 1622 1727
rect 2225 1722 2438 1727
rect 2529 1722 2678 1727
rect 2865 1722 2926 1727
rect 3065 1722 3214 1727
rect 3281 1722 3414 1727
rect 3601 1722 3638 1727
rect 1641 1717 1974 1722
rect 689 1712 838 1717
rect 1065 1712 1270 1717
rect 1585 1712 1646 1717
rect 1969 1712 2030 1717
rect 2057 1712 2214 1717
rect 2273 1712 2302 1717
rect 2441 1712 2486 1717
rect 2537 1712 2726 1717
rect 2929 1712 3070 1717
rect 3081 1712 3150 1717
rect 3177 1712 3246 1717
rect 3425 1712 3526 1717
rect 1409 1707 1478 1712
rect 2209 1707 2278 1712
rect 3633 1707 3638 1722
rect 3761 1722 3846 1727
rect 3761 1707 3766 1722
rect 3841 1717 3846 1722
rect 3953 1722 4182 1727
rect 4737 1722 4766 1727
rect 3953 1717 3958 1722
rect 3841 1712 3958 1717
rect 4137 1712 4270 1717
rect 4329 1712 4374 1717
rect 4441 1712 4486 1717
rect 4553 1712 4590 1717
rect 4625 1712 4734 1717
rect 4017 1707 4118 1712
rect 425 1702 742 1707
rect 753 1702 886 1707
rect 905 1702 1046 1707
rect 1225 1702 1414 1707
rect 1473 1702 2078 1707
rect 2625 1702 2646 1707
rect 3137 1702 3438 1707
rect 3633 1702 3766 1707
rect 3993 1702 4022 1707
rect 4113 1702 4502 1707
rect 4593 1702 4774 1707
rect 737 1697 742 1702
rect 905 1697 910 1702
rect 1041 1697 1206 1702
rect 369 1692 398 1697
rect 393 1687 398 1692
rect 529 1692 558 1697
rect 737 1692 766 1697
rect 849 1692 910 1697
rect 1201 1692 1462 1697
rect 1873 1692 2022 1697
rect 2249 1692 2678 1697
rect 2745 1692 2910 1697
rect 3073 1692 3214 1697
rect 3977 1692 4438 1697
rect 529 1687 534 1692
rect 761 1687 854 1692
rect 929 1687 1022 1692
rect 1457 1687 1462 1692
rect 1673 1687 1878 1692
rect 257 1682 334 1687
rect 393 1682 534 1687
rect 873 1682 934 1687
rect 1017 1682 1326 1687
rect 1369 1682 1390 1687
rect 1457 1682 1678 1687
rect 1897 1682 1934 1687
rect 2097 1682 2166 1687
rect 2745 1682 2750 1692
rect 2905 1687 2910 1692
rect 2905 1682 3054 1687
rect 3233 1682 3550 1687
rect 4049 1682 4078 1687
rect 4177 1682 4230 1687
rect 4369 1682 4710 1687
rect 1953 1677 2102 1682
rect 2161 1677 2166 1682
rect 2609 1677 2750 1682
rect 3049 1677 3238 1682
rect 3545 1677 3550 1682
rect 4073 1677 4182 1682
rect 4225 1677 4374 1682
rect 217 1672 246 1677
rect 561 1672 1438 1677
rect 1697 1672 1830 1677
rect 1849 1672 1958 1677
rect 2161 1672 2238 1677
rect 1697 1667 1702 1672
rect 217 1662 278 1667
rect 1457 1662 1654 1667
rect 1673 1662 1702 1667
rect 1825 1667 1830 1672
rect 2233 1667 2238 1672
rect 2345 1672 2614 1677
rect 3545 1672 3574 1677
rect 2345 1667 2350 1672
rect 1825 1662 2046 1667
rect 2233 1662 2350 1667
rect 2369 1662 2398 1667
rect 977 1657 1398 1662
rect 1457 1657 1462 1662
rect 201 1652 230 1657
rect 353 1652 438 1657
rect 681 1652 982 1657
rect 1393 1652 1462 1657
rect 1649 1657 1654 1662
rect 2393 1657 2398 1662
rect 2625 1662 3518 1667
rect 3761 1662 3798 1667
rect 3817 1662 3942 1667
rect 2625 1657 2630 1662
rect 3817 1657 3822 1662
rect 1649 1652 1814 1657
rect 1881 1652 2150 1657
rect 2393 1652 2630 1657
rect 2649 1652 2678 1657
rect 3073 1652 3158 1657
rect 353 1647 358 1652
rect 329 1642 358 1647
rect 433 1647 438 1652
rect 1809 1647 1886 1652
rect 2673 1647 2814 1652
rect 2913 1647 3078 1652
rect 3153 1647 3158 1652
rect 3513 1652 3630 1657
rect 3785 1652 3822 1657
rect 3937 1657 3942 1662
rect 4057 1662 4214 1667
rect 4057 1657 4062 1662
rect 3937 1652 4062 1657
rect 4209 1657 4214 1662
rect 4257 1662 4374 1667
rect 4257 1657 4262 1662
rect 4209 1652 4262 1657
rect 4369 1657 4374 1662
rect 4369 1652 4566 1657
rect 3513 1647 3518 1652
rect 433 1642 670 1647
rect 665 1637 670 1642
rect 993 1642 1382 1647
rect 1449 1642 1678 1647
rect 1689 1642 1742 1647
rect 1905 1642 1934 1647
rect 993 1637 998 1642
rect 1929 1637 1934 1642
rect 1993 1642 2030 1647
rect 2809 1642 2918 1647
rect 3097 1642 3134 1647
rect 3153 1642 3518 1647
rect 3769 1642 4582 1647
rect 4681 1642 4758 1647
rect 1993 1637 1998 1642
rect 177 1632 390 1637
rect 665 1632 998 1637
rect 1017 1632 1246 1637
rect 1353 1632 1398 1637
rect 1633 1632 1790 1637
rect 1929 1632 1998 1637
rect 2713 1632 2790 1637
rect 2937 1632 3118 1637
rect 3537 1632 3606 1637
rect 3705 1632 4206 1637
rect 4201 1627 4206 1632
rect 4289 1632 4622 1637
rect 4657 1632 4694 1637
rect 4289 1627 4294 1632
rect 129 1622 182 1627
rect 265 1622 310 1627
rect 377 1622 422 1627
rect 489 1622 534 1627
rect 569 1622 590 1627
rect 761 1622 830 1627
rect 985 1622 1030 1627
rect 1089 1622 1134 1627
rect 1345 1622 1478 1627
rect 1577 1622 1702 1627
rect 2049 1622 2166 1627
rect 2441 1622 2534 1627
rect 2657 1622 2710 1627
rect 3169 1622 3222 1627
rect 3329 1622 3390 1627
rect 3545 1622 4134 1627
rect 4201 1622 4294 1627
rect 4369 1622 4454 1627
rect 2049 1617 2054 1622
rect 353 1612 398 1617
rect 873 1612 942 1617
rect 201 1602 246 1607
rect 521 1602 590 1607
rect 177 1592 198 1597
rect 297 1592 430 1597
rect 457 1592 518 1597
rect 809 1592 862 1597
rect 889 1592 942 1597
rect 1153 1592 1158 1617
rect 1329 1612 1446 1617
rect 2017 1612 2054 1617
rect 2161 1617 2166 1622
rect 2161 1612 2430 1617
rect 1465 1607 1590 1612
rect 2425 1607 2430 1612
rect 2545 1612 2646 1617
rect 2545 1607 2550 1612
rect 1257 1602 1286 1607
rect 1321 1602 1470 1607
rect 1585 1602 1646 1607
rect 1657 1602 1750 1607
rect 2425 1602 2550 1607
rect 2641 1607 2646 1612
rect 2721 1612 2926 1617
rect 2721 1607 2726 1612
rect 2641 1602 2726 1607
rect 2921 1607 2926 1612
rect 2985 1612 3158 1617
rect 3249 1612 3278 1617
rect 3713 1612 3798 1617
rect 4041 1612 4102 1617
rect 4137 1612 4182 1617
rect 4609 1612 4670 1617
rect 2985 1607 2990 1612
rect 3153 1607 3254 1612
rect 3913 1607 4022 1612
rect 2921 1602 2990 1607
rect 3425 1602 3478 1607
rect 3553 1602 3574 1607
rect 3673 1602 3750 1607
rect 3569 1597 3574 1602
rect 3745 1597 3750 1602
rect 3841 1602 3918 1607
rect 4017 1602 4366 1607
rect 3841 1597 3846 1602
rect 4361 1597 4366 1602
rect 4449 1602 4534 1607
rect 4449 1597 4454 1602
rect 1417 1592 1486 1597
rect 1513 1592 1574 1597
rect 1681 1592 1710 1597
rect 1785 1592 1902 1597
rect 1921 1592 2150 1597
rect 3009 1592 3278 1597
rect 3449 1592 3558 1597
rect 3569 1592 3590 1597
rect 3681 1592 3726 1597
rect 3745 1592 3846 1597
rect 3865 1592 3974 1597
rect 4009 1592 4054 1597
rect 4073 1592 4094 1597
rect 4169 1592 4246 1597
rect 4289 1592 4342 1597
rect 4361 1592 4454 1597
rect 4473 1592 4542 1597
rect 4593 1592 4638 1597
rect 1785 1587 1790 1592
rect 401 1582 478 1587
rect 817 1582 870 1587
rect 1105 1582 1206 1587
rect 1641 1582 1790 1587
rect 1897 1587 1902 1592
rect 1897 1582 1942 1587
rect 1937 1577 1942 1582
rect 2081 1582 2654 1587
rect 2721 1582 2758 1587
rect 3017 1582 3102 1587
rect 3217 1582 3254 1587
rect 3297 1582 3398 1587
rect 3521 1582 3574 1587
rect 2081 1577 2086 1582
rect 3297 1577 3302 1582
rect 441 1572 478 1577
rect 561 1572 654 1577
rect 673 1572 694 1577
rect 1249 1572 1358 1577
rect 1617 1572 1838 1577
rect 1937 1572 2086 1577
rect 3057 1572 3110 1577
rect 3193 1572 3302 1577
rect 3393 1577 3398 1582
rect 3393 1572 3446 1577
rect 3529 1572 3614 1577
rect 3913 1572 4222 1577
rect 561 1567 566 1572
rect 289 1562 366 1567
rect 409 1562 566 1567
rect 649 1567 654 1572
rect 833 1567 910 1572
rect 2281 1567 2534 1572
rect 3913 1567 3918 1572
rect 649 1562 838 1567
rect 905 1562 934 1567
rect 1233 1562 1270 1567
rect 1441 1562 1518 1567
rect 1633 1562 1678 1567
rect 289 1557 294 1562
rect 185 1552 294 1557
rect 361 1557 366 1562
rect 1441 1557 1446 1562
rect 361 1552 390 1557
rect 673 1552 702 1557
rect 697 1547 702 1552
rect 849 1552 894 1557
rect 985 1552 1326 1557
rect 1345 1552 1446 1557
rect 1513 1557 1518 1562
rect 1673 1557 1678 1562
rect 1753 1562 1918 1567
rect 2105 1562 2238 1567
rect 2257 1562 2286 1567
rect 2529 1562 2558 1567
rect 2577 1562 2950 1567
rect 3209 1562 3462 1567
rect 3689 1562 3854 1567
rect 3873 1562 3918 1567
rect 4217 1567 4222 1572
rect 4217 1562 4246 1567
rect 4697 1562 4726 1567
rect 1753 1557 1758 1562
rect 2105 1557 2110 1562
rect 1513 1552 1654 1557
rect 1673 1552 1758 1557
rect 1825 1552 1854 1557
rect 1969 1552 2110 1557
rect 2233 1557 2238 1562
rect 2577 1557 2582 1562
rect 2233 1552 2582 1557
rect 2945 1557 2950 1562
rect 3033 1557 3190 1562
rect 2945 1552 3038 1557
rect 3185 1552 3262 1557
rect 3401 1552 3494 1557
rect 849 1547 854 1552
rect 1345 1547 1350 1552
rect 305 1542 454 1547
rect 577 1542 614 1547
rect 697 1542 854 1547
rect 1233 1542 1262 1547
rect 1289 1542 1350 1547
rect 1401 1542 1494 1547
rect 129 1532 174 1537
rect 305 1532 326 1537
rect 561 1532 606 1537
rect 873 1532 918 1537
rect 305 1527 310 1532
rect 257 1522 310 1527
rect 337 1522 366 1527
rect 913 1522 918 1532
rect 1049 1532 1206 1537
rect 1225 1532 1246 1537
rect 1377 1532 1414 1537
rect 1481 1532 1526 1537
rect 1049 1527 1054 1532
rect 977 1522 1054 1527
rect 1201 1527 1206 1532
rect 1377 1527 1382 1532
rect 1649 1527 1654 1552
rect 3689 1547 3694 1562
rect 2121 1542 2454 1547
rect 2449 1537 2454 1542
rect 2545 1542 2686 1547
rect 2729 1542 2782 1547
rect 2809 1542 2870 1547
rect 3049 1542 3102 1547
rect 3145 1542 3342 1547
rect 3665 1542 3694 1547
rect 3849 1547 3854 1562
rect 4009 1557 4198 1562
rect 3929 1552 4014 1557
rect 4193 1552 4334 1557
rect 4353 1552 4454 1557
rect 4585 1552 4798 1557
rect 4353 1547 4358 1552
rect 3849 1542 3918 1547
rect 4025 1542 4150 1547
rect 4193 1542 4358 1547
rect 4449 1547 4454 1552
rect 4449 1542 4478 1547
rect 4545 1542 4598 1547
rect 4609 1542 4638 1547
rect 4665 1542 4694 1547
rect 2545 1537 2550 1542
rect 3913 1537 4030 1542
rect 2017 1532 2142 1537
rect 2449 1532 2550 1537
rect 2737 1532 2934 1537
rect 3041 1532 3102 1537
rect 3201 1532 3230 1537
rect 3249 1532 3270 1537
rect 3697 1532 3734 1537
rect 3809 1532 3886 1537
rect 4049 1532 4086 1537
rect 4113 1532 4158 1537
rect 4233 1532 4262 1537
rect 3097 1527 3206 1532
rect 1201 1522 1254 1527
rect 1281 1522 1310 1527
rect 1377 1522 1406 1527
rect 1417 1522 1438 1527
rect 1569 1522 1598 1527
rect 1649 1522 1694 1527
rect 1929 1522 1958 1527
rect 2153 1522 2318 1527
rect 2745 1522 2798 1527
rect 2913 1522 3078 1527
rect 257 1517 262 1522
rect 977 1517 982 1522
rect 3249 1517 3254 1532
rect 4257 1527 4262 1532
rect 4345 1532 4454 1537
rect 4513 1532 4574 1537
rect 4665 1532 4718 1537
rect 4345 1527 4350 1532
rect 209 1512 262 1517
rect 273 1512 318 1517
rect 353 1512 710 1517
rect 721 1512 822 1517
rect 873 1512 982 1517
rect 1065 1512 1254 1517
rect 273 1502 342 1507
rect 705 1497 710 1512
rect 1249 1507 1254 1512
rect 1321 1512 1366 1517
rect 1729 1512 1758 1517
rect 1873 1512 1918 1517
rect 2041 1512 2070 1517
rect 1321 1507 1326 1512
rect 849 1502 878 1507
rect 969 1502 1086 1507
rect 1209 1502 1230 1507
rect 1249 1502 1326 1507
rect 1361 1507 1366 1512
rect 1601 1507 1734 1512
rect 2065 1507 2070 1512
rect 2329 1512 2598 1517
rect 2753 1512 3214 1517
rect 3249 1512 3262 1517
rect 2329 1507 2334 1512
rect 1361 1502 1606 1507
rect 2065 1502 2334 1507
rect 2881 1502 2918 1507
rect 3017 1502 3046 1507
rect 3257 1502 3262 1512
rect 3313 1507 3318 1527
rect 3329 1522 3486 1527
rect 3601 1522 3678 1527
rect 3713 1522 4070 1527
rect 4097 1522 4134 1527
rect 4257 1522 4350 1527
rect 4649 1522 4678 1527
rect 3601 1517 3606 1522
rect 3553 1512 3606 1517
rect 3673 1517 3678 1522
rect 3673 1512 3846 1517
rect 4025 1512 4054 1517
rect 4665 1512 4726 1517
rect 4769 1512 4790 1517
rect 3281 1502 3318 1507
rect 3457 1502 3910 1507
rect 4369 1502 4406 1507
rect 849 1497 854 1502
rect 705 1492 854 1497
rect 1649 1492 1718 1497
rect 1649 1487 1654 1492
rect 153 1482 238 1487
rect 513 1482 534 1487
rect 1145 1482 1182 1487
rect 1625 1482 1654 1487
rect 1713 1487 1718 1492
rect 1905 1492 1982 1497
rect 2529 1492 2558 1497
rect 3689 1492 4358 1497
rect 4417 1492 4486 1497
rect 1905 1487 1910 1492
rect 1713 1482 1910 1487
rect 1977 1487 1982 1492
rect 4353 1487 4422 1492
rect 1977 1482 2006 1487
rect 2209 1482 2382 1487
rect 3065 1482 3238 1487
rect 3065 1477 3070 1482
rect 481 1472 638 1477
rect 1377 1472 1702 1477
rect 1697 1467 1702 1472
rect 1921 1472 2182 1477
rect 2337 1472 3070 1477
rect 3233 1477 3238 1482
rect 3337 1482 3670 1487
rect 3337 1477 3342 1482
rect 3665 1477 3750 1482
rect 3801 1477 3894 1482
rect 3233 1472 3342 1477
rect 3745 1472 3806 1477
rect 3889 1472 4046 1477
rect 1921 1467 1926 1472
rect 4041 1467 4046 1472
rect 4353 1472 4382 1477
rect 4353 1467 4358 1472
rect 417 1462 494 1467
rect 657 1462 790 1467
rect 1697 1462 1926 1467
rect 2961 1462 2990 1467
rect 657 1457 662 1462
rect 313 1452 430 1457
rect 537 1452 662 1457
rect 537 1447 542 1452
rect 113 1442 150 1447
rect 433 1442 542 1447
rect 785 1447 790 1462
rect 2985 1457 2990 1462
rect 3057 1462 3734 1467
rect 3817 1462 3878 1467
rect 4041 1462 4358 1467
rect 3057 1457 3062 1462
rect 3729 1457 3822 1462
rect 1209 1452 1278 1457
rect 1945 1452 2038 1457
rect 2201 1452 2270 1457
rect 2985 1452 3062 1457
rect 3217 1452 3254 1457
rect 3361 1452 3574 1457
rect 1209 1447 1214 1452
rect 785 1442 854 1447
rect 1185 1442 1214 1447
rect 1273 1447 1278 1452
rect 2201 1447 2206 1452
rect 1273 1442 1454 1447
rect 1857 1442 2206 1447
rect 2265 1447 2270 1452
rect 3105 1447 3198 1452
rect 3593 1447 3710 1452
rect 2265 1442 2918 1447
rect 3081 1442 3110 1447
rect 3193 1442 3382 1447
rect 3409 1442 3598 1447
rect 3705 1442 4022 1447
rect 161 1432 310 1437
rect 553 1432 774 1437
rect 873 1432 966 1437
rect 1089 1432 1262 1437
rect 1769 1432 1982 1437
rect 2193 1432 2254 1437
rect 2993 1432 3062 1437
rect 3089 1432 3222 1437
rect 873 1427 878 1432
rect 129 1422 174 1427
rect 465 1422 518 1427
rect 537 1422 598 1427
rect 809 1422 878 1427
rect 961 1427 966 1432
rect 2657 1427 2766 1432
rect 2993 1427 2998 1432
rect 961 1422 1134 1427
rect 1161 1422 1246 1427
rect 1401 1422 1462 1427
rect 1505 1422 1550 1427
rect 1833 1422 1878 1427
rect 1961 1422 1998 1427
rect 2089 1422 2118 1427
rect 2633 1422 2662 1427
rect 2761 1422 2814 1427
rect 2113 1417 2118 1422
rect 2809 1417 2814 1422
rect 2905 1422 2998 1427
rect 3009 1422 3054 1427
rect 3129 1422 3166 1427
rect 3241 1422 3334 1427
rect 2905 1417 2910 1422
rect 3241 1417 3246 1422
rect 569 1412 606 1417
rect 649 1412 686 1417
rect 817 1412 870 1417
rect 1177 1412 1198 1417
rect 1241 1412 1302 1417
rect 1705 1407 1710 1417
rect 1857 1412 1902 1417
rect 2113 1412 2166 1417
rect 2521 1412 2590 1417
rect 2657 1412 2782 1417
rect 2809 1412 2910 1417
rect 2929 1412 3086 1417
rect 3169 1412 3246 1417
rect 3329 1417 3334 1422
rect 3441 1417 3446 1437
rect 3529 1432 3590 1437
rect 3609 1432 3694 1437
rect 4521 1432 4590 1437
rect 3841 1422 3934 1427
rect 4057 1422 4126 1427
rect 4137 1422 4238 1427
rect 4257 1422 4438 1427
rect 4497 1422 4694 1427
rect 3465 1417 3630 1422
rect 3841 1417 3846 1422
rect 3329 1412 3358 1417
rect 3441 1412 3470 1417
rect 3625 1412 3654 1417
rect 3721 1412 3758 1417
rect 3817 1412 3846 1417
rect 3929 1417 3934 1422
rect 4257 1417 4262 1422
rect 3929 1412 4078 1417
rect 4113 1412 4262 1417
rect 4433 1417 4438 1422
rect 4433 1412 4558 1417
rect 4761 1412 4790 1417
rect 145 1402 166 1407
rect 689 1402 950 1407
rect 1089 1402 1294 1407
rect 1705 1402 1734 1407
rect 2201 1402 2254 1407
rect 3041 1402 3134 1407
rect 3209 1402 3398 1407
rect 3409 1402 3710 1407
rect 3857 1402 3974 1407
rect 4121 1402 4166 1407
rect 4281 1402 4358 1407
rect 3705 1397 3862 1402
rect 497 1392 646 1397
rect 697 1392 838 1397
rect 1153 1392 1198 1397
rect 1393 1392 1518 1397
rect 1577 1392 1670 1397
rect 1809 1392 1846 1397
rect 2417 1392 2790 1397
rect 2993 1392 3118 1397
rect 3289 1392 3390 1397
rect 3513 1392 3566 1397
rect 3657 1392 3686 1397
rect 4001 1392 4422 1397
rect 4489 1392 4526 1397
rect 4665 1392 4694 1397
rect 1217 1387 1350 1392
rect 441 1382 470 1387
rect 593 1382 622 1387
rect 641 1382 670 1387
rect 865 1382 894 1387
rect 945 1382 982 1387
rect 993 1382 1222 1387
rect 1345 1382 1454 1387
rect 3065 1382 3238 1387
rect 3273 1382 3310 1387
rect 3401 1382 3510 1387
rect 3529 1382 3566 1387
rect 3745 1382 3990 1387
rect 465 1377 598 1382
rect 665 1377 670 1382
rect 729 1377 870 1382
rect 3305 1377 3406 1382
rect 3985 1377 3990 1382
rect 4081 1382 4166 1387
rect 4081 1377 4086 1382
rect 4161 1377 4166 1382
rect 4321 1382 4486 1387
rect 4649 1382 4686 1387
rect 4321 1377 4326 1382
rect 89 1372 126 1377
rect 665 1372 734 1377
rect 929 1372 958 1377
rect 225 1362 262 1367
rect 513 1362 574 1367
rect 753 1362 798 1367
rect 953 1357 958 1372
rect 1137 1372 1334 1377
rect 1137 1357 1142 1372
rect 1329 1367 1334 1372
rect 1441 1372 1670 1377
rect 2649 1372 2678 1377
rect 2729 1372 2758 1377
rect 3193 1372 3286 1377
rect 3481 1372 3670 1377
rect 3985 1372 4086 1377
rect 4105 1372 4142 1377
rect 4161 1372 4326 1377
rect 4345 1372 4502 1377
rect 1441 1367 1446 1372
rect 1217 1362 1270 1367
rect 1329 1362 1446 1367
rect 2377 1362 2550 1367
rect 2673 1362 2718 1367
rect 2809 1362 2910 1367
rect 3225 1362 3390 1367
rect 3545 1362 3694 1367
rect 3865 1362 3934 1367
rect 3929 1357 3934 1362
rect 4369 1362 4438 1367
rect 4457 1362 4510 1367
rect 4369 1357 4374 1362
rect 321 1352 782 1357
rect 953 1352 1142 1357
rect 1201 1352 1246 1357
rect 1265 1352 1310 1357
rect 1465 1352 1542 1357
rect 1681 1352 1894 1357
rect 2393 1352 2422 1357
rect 2529 1352 2750 1357
rect 2889 1352 3006 1357
rect 3177 1352 3206 1357
rect 3377 1352 3422 1357
rect 3489 1352 3566 1357
rect 3561 1347 3566 1352
rect 3705 1352 3838 1357
rect 3929 1352 4374 1357
rect 3705 1347 3710 1352
rect 553 1342 606 1347
rect 673 1342 694 1347
rect 761 1342 806 1347
rect 1161 1342 1238 1347
rect 1257 1342 1318 1347
rect 1337 1342 1414 1347
rect 1497 1342 1598 1347
rect 1721 1342 1750 1347
rect 2185 1342 2214 1347
rect 2401 1342 2542 1347
rect 2897 1342 2934 1347
rect 2977 1342 3022 1347
rect 3049 1342 3126 1347
rect 3169 1342 3270 1347
rect 3521 1342 3542 1347
rect 3561 1342 3710 1347
rect 3873 1342 3910 1347
rect 4393 1342 4478 1347
rect 4657 1342 4774 1347
rect 1337 1337 1342 1342
rect 169 1332 334 1337
rect 673 1332 702 1337
rect 1281 1332 1342 1337
rect 1409 1337 1414 1342
rect 1409 1332 1678 1337
rect 1769 1332 1838 1337
rect 2177 1332 2198 1337
rect 1769 1327 1774 1332
rect 1649 1322 1774 1327
rect 1833 1327 1838 1332
rect 1833 1322 2006 1327
rect 137 1312 182 1317
rect 337 1312 446 1317
rect 545 1312 582 1317
rect 609 1312 646 1317
rect 1185 1312 1278 1317
rect 1289 1312 1398 1317
rect 1465 1312 1638 1317
rect 1737 1312 1766 1317
rect 1777 1312 1822 1317
rect 2193 1312 2198 1332
rect 2209 1312 2214 1342
rect 3785 1332 3862 1337
rect 4481 1332 4566 1337
rect 3121 1327 3278 1332
rect 2465 1322 2486 1327
rect 3097 1322 3126 1327
rect 3273 1322 3494 1327
rect 3881 1322 3910 1327
rect 4073 1322 4174 1327
rect 4257 1322 4438 1327
rect 4497 1322 4526 1327
rect 4537 1322 4566 1327
rect 2481 1307 2486 1322
rect 2617 1312 2694 1317
rect 3121 1312 3182 1317
rect 3241 1312 3262 1317
rect 3569 1312 3694 1317
rect 3817 1312 3862 1317
rect 4113 1312 4150 1317
rect 4265 1312 4286 1317
rect 4673 1312 4742 1317
rect 265 1302 326 1307
rect 321 1287 326 1302
rect 529 1302 614 1307
rect 633 1302 694 1307
rect 1721 1302 1750 1307
rect 529 1287 534 1302
rect 609 1297 614 1302
rect 1201 1297 1462 1302
rect 1745 1297 1750 1302
rect 2001 1302 2030 1307
rect 2353 1302 2438 1307
rect 2457 1302 2486 1307
rect 2697 1302 2758 1307
rect 2793 1302 2846 1307
rect 3169 1302 3214 1307
rect 3697 1302 3790 1307
rect 3913 1302 3998 1307
rect 4041 1302 4070 1307
rect 4129 1302 4294 1307
rect 2001 1297 2006 1302
rect 609 1292 782 1297
rect 921 1292 990 1297
rect 1017 1292 1206 1297
rect 1457 1292 1566 1297
rect 1745 1292 2006 1297
rect 2585 1292 2670 1297
rect 921 1287 926 1292
rect 321 1282 534 1287
rect 649 1282 742 1287
rect 777 1282 926 1287
rect 985 1287 990 1292
rect 985 1282 1006 1287
rect 937 1272 974 1277
rect 1001 1267 1006 1282
rect 1217 1282 1270 1287
rect 1217 1267 1222 1282
rect 1265 1277 1270 1282
rect 1433 1282 1462 1287
rect 1433 1277 1438 1282
rect 1265 1272 1294 1277
rect 1409 1272 1438 1277
rect 2265 1272 2310 1277
rect 4553 1272 4638 1277
rect 1289 1267 1414 1272
rect 1001 1262 1222 1267
rect 3969 1262 4182 1267
rect 3969 1257 3974 1262
rect 1305 1252 1534 1257
rect 2305 1252 2534 1257
rect 3785 1252 3974 1257
rect 4177 1257 4182 1262
rect 4289 1262 4374 1267
rect 4289 1257 4294 1262
rect 4177 1252 4294 1257
rect 4369 1257 4374 1262
rect 4369 1252 4750 1257
rect 1241 1242 1286 1247
rect 1305 1237 1310 1252
rect 1529 1237 1534 1252
rect 1553 1242 1638 1247
rect 2321 1242 2350 1247
rect 2617 1242 2646 1247
rect 265 1232 302 1237
rect 817 1232 894 1237
rect 1265 1232 1310 1237
rect 1329 1232 1510 1237
rect 1529 1232 1654 1237
rect 2545 1232 2638 1237
rect 2865 1232 2910 1237
rect 3009 1232 3070 1237
rect 3985 1232 4166 1237
rect 1329 1227 1334 1232
rect 185 1222 374 1227
rect 537 1222 582 1227
rect 649 1222 702 1227
rect 729 1222 766 1227
rect 881 1222 934 1227
rect 1129 1222 1214 1227
rect 1225 1222 1334 1227
rect 1505 1227 1510 1232
rect 4161 1227 4166 1232
rect 4305 1232 4358 1237
rect 4609 1232 4686 1237
rect 4305 1227 4310 1232
rect 4609 1227 4614 1232
rect 1505 1222 1630 1227
rect 1657 1222 1758 1227
rect 2449 1222 2494 1227
rect 2513 1222 2582 1227
rect 2633 1222 2742 1227
rect 2801 1222 2854 1227
rect 3553 1222 3630 1227
rect 3729 1222 3958 1227
rect 4161 1222 4310 1227
rect 4329 1222 4614 1227
rect 1393 1217 1486 1222
rect 3729 1217 3734 1222
rect 105 1212 358 1217
rect 665 1212 822 1217
rect 953 1212 1022 1217
rect 1257 1212 1286 1217
rect 1297 1212 1398 1217
rect 1481 1212 1718 1217
rect 2217 1212 2246 1217
rect 2553 1212 2590 1217
rect 2721 1212 2830 1217
rect 3673 1212 3734 1217
rect 3953 1217 3958 1222
rect 3953 1212 4142 1217
rect 4481 1212 4550 1217
rect 953 1207 958 1212
rect 737 1202 958 1207
rect 1017 1207 1022 1212
rect 1297 1207 1302 1212
rect 1017 1202 1054 1207
rect 1121 1202 1302 1207
rect 1345 1202 1494 1207
rect 1617 1202 1646 1207
rect 249 1197 334 1202
rect 1641 1197 1646 1202
rect 1729 1202 1806 1207
rect 2353 1202 2486 1207
rect 2497 1202 2526 1207
rect 2873 1202 2998 1207
rect 3633 1202 3662 1207
rect 3745 1202 3854 1207
rect 4473 1202 4526 1207
rect 1729 1197 1734 1202
rect 3657 1197 3750 1202
rect 3969 1197 4118 1202
rect 225 1192 254 1197
rect 329 1192 414 1197
rect 801 1192 862 1197
rect 969 1192 1006 1197
rect 1233 1192 1262 1197
rect 1273 1192 1390 1197
rect 1457 1192 1486 1197
rect 1481 1187 1486 1192
rect 1569 1192 1598 1197
rect 1641 1192 1734 1197
rect 1865 1192 1966 1197
rect 2217 1192 2334 1197
rect 2801 1192 2870 1197
rect 1569 1187 1574 1192
rect 2865 1187 2870 1192
rect 3009 1192 3102 1197
rect 3889 1192 3974 1197
rect 4113 1192 4142 1197
rect 4233 1192 4422 1197
rect 4441 1192 4470 1197
rect 4537 1192 4590 1197
rect 3009 1187 3014 1192
rect 193 1182 318 1187
rect 433 1182 550 1187
rect 569 1182 702 1187
rect 1217 1182 1278 1187
rect 1393 1182 1454 1187
rect 1481 1182 1574 1187
rect 2193 1182 2214 1187
rect 2865 1182 3014 1187
rect 3521 1182 3734 1187
rect 3985 1182 4086 1187
rect 4401 1182 4550 1187
rect 433 1177 438 1182
rect 297 1172 438 1177
rect 545 1177 550 1182
rect 3729 1177 3734 1182
rect 3881 1177 3990 1182
rect 4105 1177 4182 1182
rect 4401 1177 4406 1182
rect 545 1172 958 1177
rect 953 1167 958 1172
rect 1017 1172 1094 1177
rect 1249 1172 1358 1177
rect 1601 1172 1854 1177
rect 1017 1167 1022 1172
rect 233 1162 262 1167
rect 449 1162 678 1167
rect 697 1162 758 1167
rect 953 1162 1022 1167
rect 1849 1167 1854 1172
rect 1953 1172 2070 1177
rect 2497 1172 2590 1177
rect 2609 1172 2670 1177
rect 3601 1172 3710 1177
rect 3729 1172 3886 1177
rect 4065 1172 4110 1177
rect 4177 1172 4406 1177
rect 4417 1172 4710 1177
rect 1953 1167 1958 1172
rect 2497 1167 2502 1172
rect 1849 1162 1958 1167
rect 2089 1162 2230 1167
rect 2393 1162 2502 1167
rect 2585 1167 2590 1172
rect 2585 1162 2646 1167
rect 2849 1162 3006 1167
rect 3345 1162 3470 1167
rect 3905 1162 4038 1167
rect 4081 1162 4166 1167
rect 4537 1162 4582 1167
rect 257 1157 454 1162
rect 673 1157 678 1162
rect 673 1152 870 1157
rect 1073 1152 1158 1157
rect 1473 1152 1502 1157
rect 1625 1152 1774 1157
rect 2985 1152 3022 1157
rect 3081 1152 3150 1157
rect 3217 1152 3334 1157
rect 1073 1147 1078 1152
rect 257 1142 358 1147
rect 457 1142 486 1147
rect 481 1137 486 1142
rect 649 1142 918 1147
rect 1049 1142 1078 1147
rect 1153 1147 1158 1152
rect 3345 1147 3350 1162
rect 3465 1157 3470 1162
rect 3465 1152 3494 1157
rect 4193 1152 4278 1157
rect 4297 1152 4334 1157
rect 4353 1152 4486 1157
rect 4577 1152 4654 1157
rect 4193 1147 4198 1152
rect 1153 1142 1182 1147
rect 1305 1142 1358 1147
rect 1689 1142 1734 1147
rect 1977 1142 2054 1147
rect 2513 1142 2590 1147
rect 649 1137 654 1142
rect 2585 1137 2590 1142
rect 2657 1142 2742 1147
rect 2865 1142 3350 1147
rect 3377 1142 3478 1147
rect 3857 1142 3910 1147
rect 3969 1142 4022 1147
rect 4177 1142 4198 1147
rect 4273 1147 4278 1152
rect 4353 1147 4358 1152
rect 4273 1142 4358 1147
rect 4481 1147 4486 1152
rect 4481 1142 4590 1147
rect 2657 1137 2662 1142
rect 4177 1137 4182 1142
rect 481 1132 654 1137
rect 673 1132 702 1137
rect 697 1127 702 1132
rect 769 1132 878 1137
rect 1001 1132 1070 1137
rect 1121 1132 1158 1137
rect 1169 1132 1190 1137
rect 1545 1132 1638 1137
rect 1665 1132 1750 1137
rect 2097 1132 2206 1137
rect 2585 1132 2662 1137
rect 2881 1132 2910 1137
rect 3081 1132 3214 1137
rect 3321 1132 3390 1137
rect 3505 1132 4182 1137
rect 4217 1132 4470 1137
rect 769 1127 774 1132
rect 1121 1127 1126 1132
rect 193 1122 214 1127
rect 697 1122 774 1127
rect 793 1122 838 1127
rect 897 1122 950 1127
rect 1097 1122 1126 1127
rect 1145 1122 1166 1127
rect 1185 1117 1190 1132
rect 2905 1127 2910 1132
rect 3001 1127 3086 1132
rect 4465 1127 4470 1132
rect 4561 1132 4774 1137
rect 4561 1127 4566 1132
rect 1617 1122 1646 1127
rect 1801 1122 1918 1127
rect 1953 1122 2006 1127
rect 2193 1122 2254 1127
rect 2433 1122 2454 1127
rect 2905 1122 3006 1127
rect 3105 1122 3342 1127
rect 3505 1122 3550 1127
rect 3809 1122 3902 1127
rect 3969 1122 4102 1127
rect 4321 1122 4342 1127
rect 4465 1122 4566 1127
rect 4585 1122 4606 1127
rect 1681 1117 1774 1122
rect 97 1112 214 1117
rect 265 1112 310 1117
rect 865 1112 894 1117
rect 889 1107 894 1112
rect 969 1112 1126 1117
rect 1153 1112 1190 1117
rect 1609 1112 1686 1117
rect 1769 1112 1790 1117
rect 1881 1112 1966 1117
rect 2057 1112 2102 1117
rect 969 1107 974 1112
rect 1785 1107 1886 1112
rect 177 1102 230 1107
rect 281 1102 654 1107
rect 745 1102 790 1107
rect 825 1102 854 1107
rect 889 1102 974 1107
rect 1017 1102 1070 1107
rect 1081 1102 1182 1107
rect 1537 1102 1598 1107
rect 1697 1102 1758 1107
rect 1905 1102 1998 1107
rect 2177 1102 2222 1107
rect 2449 1102 2454 1122
rect 2529 1112 2566 1117
rect 2753 1112 2886 1117
rect 3065 1112 3110 1117
rect 3105 1107 3110 1112
rect 3177 1112 3206 1117
rect 3217 1112 3310 1117
rect 3369 1112 3486 1117
rect 3817 1112 3870 1117
rect 3945 1112 3990 1117
rect 4225 1112 4286 1117
rect 4361 1112 4446 1117
rect 3177 1107 3182 1112
rect 2473 1102 2502 1107
rect 3025 1102 3086 1107
rect 3105 1102 3182 1107
rect 3225 1102 3278 1107
rect 3561 1102 3670 1107
rect 4073 1102 4302 1107
rect 4345 1102 4374 1107
rect 4369 1097 4374 1102
rect 4457 1102 4694 1107
rect 4457 1097 4462 1102
rect 777 1092 846 1097
rect 1049 1092 1118 1097
rect 1209 1092 1518 1097
rect 1713 1092 1958 1097
rect 1969 1092 2014 1097
rect 2185 1092 2510 1097
rect 4369 1092 4462 1097
rect 681 1082 710 1087
rect 993 1082 1030 1087
rect 1209 1077 1214 1092
rect 1513 1087 1518 1092
rect 1953 1087 1958 1092
rect 1513 1082 1670 1087
rect 1953 1082 2038 1087
rect 2169 1082 2214 1087
rect 2497 1082 2614 1087
rect 3633 1082 3974 1087
rect 953 1072 1214 1077
rect 1665 1077 1670 1082
rect 1665 1072 1694 1077
rect 1713 1072 1934 1077
rect 2057 1072 2142 1077
rect 4057 1072 4166 1077
rect 1537 1067 1646 1072
rect 1713 1067 1718 1072
rect 1929 1067 2062 1072
rect 2137 1067 2142 1072
rect 3769 1067 4014 1072
rect 4057 1067 4062 1072
rect 705 1062 1094 1067
rect 1225 1062 1542 1067
rect 1641 1062 1718 1067
rect 2137 1062 2166 1067
rect 2233 1062 2358 1067
rect 3745 1062 3774 1067
rect 4009 1062 4062 1067
rect 4161 1067 4166 1072
rect 4161 1062 4190 1067
rect 1089 1057 1230 1062
rect 1801 1057 1910 1062
rect 2233 1057 2238 1062
rect 297 1052 358 1057
rect 473 1052 630 1057
rect 1553 1052 1582 1057
rect 1601 1052 1806 1057
rect 1905 1052 2022 1057
rect 2057 1052 2150 1057
rect 2209 1052 2238 1057
rect 2353 1057 2358 1062
rect 2353 1052 2382 1057
rect 2729 1052 2838 1057
rect 2857 1052 2878 1057
rect 3513 1052 3662 1057
rect 3681 1052 4254 1057
rect 4369 1052 4622 1057
rect 273 1037 430 1042
rect 473 1037 478 1052
rect 249 1032 278 1037
rect 425 1032 478 1037
rect 625 1037 630 1052
rect 937 1047 1070 1052
rect 1601 1047 1606 1052
rect 2729 1047 2734 1052
rect 769 1042 894 1047
rect 913 1042 942 1047
rect 1065 1042 1606 1047
rect 1617 1042 2030 1047
rect 2105 1042 2150 1047
rect 2161 1042 2358 1047
rect 2601 1042 2646 1047
rect 2681 1042 2734 1047
rect 2833 1047 2838 1052
rect 3513 1047 3518 1052
rect 2833 1042 2870 1047
rect 3377 1042 3470 1047
rect 3489 1042 3518 1047
rect 3657 1047 3662 1052
rect 3657 1042 3782 1047
rect 3793 1042 4310 1047
rect 769 1037 774 1042
rect 625 1032 774 1037
rect 889 1037 894 1042
rect 889 1032 1270 1037
rect 169 1022 230 1027
rect 241 1022 390 1027
rect 425 1022 614 1027
rect 785 1022 830 1027
rect 849 1022 918 1027
rect 1009 1022 1062 1027
rect 1145 1022 1190 1027
rect 633 1017 702 1022
rect 849 1017 854 1022
rect 1265 1017 1270 1032
rect 1617 1017 1622 1042
rect 3377 1037 3382 1042
rect 1641 1032 1974 1037
rect 1969 1027 1974 1032
rect 2113 1032 2142 1037
rect 2177 1032 2270 1037
rect 2761 1032 2854 1037
rect 2865 1032 2902 1037
rect 3025 1032 3054 1037
rect 3073 1032 3182 1037
rect 3257 1032 3382 1037
rect 3465 1037 3470 1042
rect 4369 1037 4374 1052
rect 4617 1047 4622 1052
rect 4617 1042 4678 1047
rect 3465 1032 3646 1037
rect 3665 1032 4374 1037
rect 4393 1032 4422 1037
rect 2113 1027 2118 1032
rect 3073 1027 3078 1032
rect 1673 1022 1878 1027
rect 1889 1022 1950 1027
rect 1969 1022 2118 1027
rect 2273 1022 2318 1027
rect 2561 1022 2606 1027
rect 2745 1022 2774 1027
rect 1873 1017 1878 1022
rect 2769 1017 2774 1022
rect 2873 1022 3078 1027
rect 3089 1022 3118 1027
rect 3297 1022 3326 1027
rect 3393 1022 3542 1027
rect 3657 1022 3742 1027
rect 3761 1022 3798 1027
rect 3961 1022 4030 1027
rect 4185 1022 4326 1027
rect 4369 1022 4414 1027
rect 4441 1022 4566 1027
rect 4625 1022 4662 1027
rect 2873 1017 2878 1022
rect 3321 1017 3398 1022
rect 393 1012 478 1017
rect 609 1012 638 1017
rect 697 1012 854 1017
rect 873 1012 894 1017
rect 937 1012 998 1017
rect 1073 1012 1134 1017
rect 1217 1012 1246 1017
rect 1265 1012 1622 1017
rect 1713 1012 1774 1017
rect 1873 1012 1934 1017
rect 2769 1012 2878 1017
rect 3105 1012 3174 1017
rect 993 1007 1078 1012
rect 1129 1007 1222 1012
rect 3729 1007 3734 1017
rect 3753 1012 3830 1017
rect 4385 1012 4406 1017
rect 4497 1012 4518 1017
rect 4553 1012 4654 1017
rect 4401 1007 4406 1012
rect 193 1002 246 1007
rect 345 1002 422 1007
rect 657 1002 686 1007
rect 769 1002 894 1007
rect 2361 1002 2438 1007
rect 2449 1002 2486 1007
rect 2625 997 2630 1007
rect 3105 1002 3230 1007
rect 3345 1002 3462 1007
rect 3729 1002 3750 1007
rect 3793 1002 3854 1007
rect 4057 1002 4110 1007
rect 4289 1002 4358 1007
rect 4377 1002 4406 1007
rect 4505 1002 4566 1007
rect 4289 997 4294 1002
rect 201 992 278 997
rect 473 992 502 997
rect 593 992 630 997
rect 729 992 886 997
rect 961 992 998 997
rect 1081 992 1190 997
rect 1913 992 1998 997
rect 2193 992 2222 997
rect 2353 992 2406 997
rect 2497 992 2574 997
rect 2625 992 2726 997
rect 2897 992 2998 997
rect 3057 992 3182 997
rect 3209 992 3374 997
rect 217 982 414 987
rect 449 982 590 987
rect 697 982 814 987
rect 833 982 902 987
rect 1113 982 1678 987
rect 2193 982 2342 987
rect 65 972 94 977
rect 177 972 214 977
rect 257 972 286 977
rect 185 962 238 967
rect 281 957 286 972
rect 633 972 1134 977
rect 2225 972 2254 977
rect 633 957 638 972
rect 1241 967 1454 972
rect 2337 967 2342 982
rect 2497 967 2502 992
rect 2625 987 2630 992
rect 2897 987 2902 992
rect 2521 982 2630 987
rect 2689 982 2734 987
rect 2873 982 2902 987
rect 2993 987 2998 992
rect 3369 987 3374 992
rect 3457 992 3574 997
rect 3737 992 3790 997
rect 3929 992 4046 997
rect 4145 992 4198 997
rect 4249 992 4294 997
rect 4353 997 4358 1002
rect 4353 992 4398 997
rect 4449 992 4502 997
rect 4641 992 4798 997
rect 3457 987 3462 992
rect 2993 982 3022 987
rect 3065 982 3102 987
rect 3369 982 3462 987
rect 3609 982 3678 987
rect 3729 982 3822 987
rect 4305 982 4446 987
rect 4457 982 4510 987
rect 4609 982 4646 987
rect 3937 977 4286 982
rect 2577 972 2646 977
rect 2841 972 2870 977
rect 2865 967 2870 972
rect 2953 972 2990 977
rect 3241 972 3350 977
rect 3721 972 3774 977
rect 3849 972 3942 977
rect 4281 972 4486 977
rect 4737 972 4758 977
rect 2953 967 2958 972
rect 4505 967 4638 972
rect 921 962 966 967
rect 1217 962 1246 967
rect 1449 962 1478 967
rect 681 957 758 962
rect 817 957 902 962
rect 1473 957 1478 962
rect 1617 962 1654 967
rect 1961 962 2014 967
rect 2049 962 2086 967
rect 2225 962 2302 967
rect 2337 962 2502 967
rect 2649 962 2678 967
rect 2865 962 2958 967
rect 2977 962 3710 967
rect 3857 962 3886 967
rect 1617 957 1622 962
rect 3881 957 3886 962
rect 3953 962 4326 967
rect 4393 962 4510 967
rect 4633 962 4662 967
rect 3953 957 3958 962
rect 281 952 638 957
rect 657 952 686 957
rect 753 952 822 957
rect 897 952 1014 957
rect 1281 952 1438 957
rect 1473 952 1622 957
rect 1641 952 1702 957
rect 2097 952 2134 957
rect 3161 952 3238 957
rect 3881 952 3958 957
rect 4041 952 4222 957
rect 4217 947 4222 952
rect 4305 952 4398 957
rect 4457 952 4598 957
rect 4305 947 4310 952
rect 713 942 742 947
rect 737 937 742 942
rect 833 942 862 947
rect 873 942 934 947
rect 1297 942 1366 947
rect 1417 942 1454 947
rect 3137 942 3158 947
rect 3217 942 3262 947
rect 3321 942 3510 947
rect 3697 942 3758 947
rect 3977 942 4030 947
rect 4057 942 4102 947
rect 4145 942 4198 947
rect 4217 942 4310 947
rect 4329 942 4462 947
rect 4545 942 4574 947
rect 833 937 838 942
rect 169 932 222 937
rect 737 932 838 937
rect 1385 932 1446 937
rect 1729 932 1878 937
rect 89 922 294 927
rect 1161 922 1198 927
rect 1345 922 1670 927
rect 137 912 182 917
rect 193 912 222 917
rect 337 912 382 917
rect 553 912 598 917
rect 689 912 758 917
rect 777 912 822 917
rect 913 912 982 917
rect 1105 912 1238 917
rect 1401 912 1438 917
rect 1665 912 1670 922
rect 1729 917 1734 932
rect 1705 912 1734 917
rect 1873 917 1878 932
rect 2569 932 2654 937
rect 2753 932 2854 937
rect 3081 932 3126 937
rect 2569 927 2574 932
rect 2273 922 2310 927
rect 2329 922 2446 927
rect 2545 922 2574 927
rect 2649 927 2654 932
rect 3137 927 3142 942
rect 3161 932 3342 937
rect 3593 932 3686 937
rect 3777 932 3958 937
rect 3777 927 3782 932
rect 2649 922 2734 927
rect 3137 922 3158 927
rect 3217 922 3310 927
rect 3329 922 3390 927
rect 3409 922 3478 927
rect 3713 922 3782 927
rect 3953 927 3958 932
rect 3953 922 3998 927
rect 4017 922 4134 927
rect 4153 922 4262 927
rect 4273 922 4366 927
rect 4409 922 4438 927
rect 4537 922 4590 927
rect 2329 917 2334 922
rect 1873 912 1902 917
rect 2009 912 2086 917
rect 2161 912 2334 917
rect 2441 917 2446 922
rect 3409 917 3414 922
rect 2441 912 2470 917
rect 2505 912 2614 917
rect 3065 912 3150 917
rect 3265 912 3414 917
rect 3473 917 3478 922
rect 4017 917 4022 922
rect 3473 912 3502 917
rect 3521 912 3638 917
rect 3657 912 4022 917
rect 4129 917 4134 922
rect 4129 912 4406 917
rect 4425 912 4454 917
rect 4505 912 4566 917
rect 4769 912 4790 917
rect 689 907 694 912
rect 185 902 214 907
rect 209 887 214 902
rect 393 902 614 907
rect 665 902 694 907
rect 753 907 758 912
rect 2009 907 2014 912
rect 753 902 806 907
rect 825 902 870 907
rect 1097 902 1190 907
rect 1209 902 1342 907
rect 1369 902 1454 907
rect 1713 902 2014 907
rect 2081 907 2086 912
rect 3521 907 3526 912
rect 2081 902 2110 907
rect 2305 902 2326 907
rect 2481 902 2638 907
rect 3073 902 3118 907
rect 3289 902 3526 907
rect 3633 907 3638 912
rect 4401 907 4406 912
rect 3633 902 3806 907
rect 3993 902 4166 907
rect 4177 902 4214 907
rect 4281 902 4390 907
rect 4401 902 4614 907
rect 393 887 398 902
rect 209 882 398 887
rect 609 887 614 902
rect 1713 897 1718 902
rect 2345 897 2462 902
rect 3825 897 3974 902
rect 4385 897 4390 902
rect 713 892 790 897
rect 905 892 1118 897
rect 1145 892 1246 897
rect 1329 892 1718 897
rect 2185 892 2350 897
rect 2457 892 2590 897
rect 3369 892 3830 897
rect 3969 892 4094 897
rect 4193 892 4358 897
rect 4385 892 4518 897
rect 4553 892 4678 897
rect 713 887 718 892
rect 785 887 910 892
rect 3209 887 3302 892
rect 4353 887 4358 892
rect 609 882 718 887
rect 737 882 766 887
rect 761 877 766 882
rect 1137 882 1166 887
rect 2025 882 2182 887
rect 2281 882 2526 887
rect 2849 882 3062 887
rect 1137 877 1142 882
rect 1321 877 1454 882
rect 3057 877 3062 882
rect 3129 882 3214 887
rect 3297 882 3326 887
rect 3361 882 3398 887
rect 3489 882 4126 887
rect 4353 882 4382 887
rect 4489 882 4598 887
rect 3129 877 3134 882
rect 4377 877 4494 882
rect 761 872 1142 877
rect 1297 872 1326 877
rect 1449 872 1478 877
rect 1497 872 1678 877
rect 1697 872 1974 877
rect 2417 872 2478 877
rect 3057 872 3134 877
rect 3225 872 3302 877
rect 1497 867 1502 872
rect 1185 862 1278 867
rect 1313 862 1502 867
rect 1673 867 1678 872
rect 3297 867 3302 872
rect 3393 872 3478 877
rect 3393 867 3398 872
rect 1673 862 1726 867
rect 3297 862 3398 867
rect 3473 867 3478 872
rect 3561 872 3654 877
rect 3753 872 4078 877
rect 3561 867 3566 872
rect 3649 867 3758 872
rect 3473 862 3566 867
rect 3777 862 3950 867
rect 4089 862 4494 867
rect 1185 857 1190 862
rect 745 852 1190 857
rect 1273 857 1278 862
rect 1537 857 1654 862
rect 1745 857 1958 862
rect 3945 857 4094 862
rect 1273 852 1302 857
rect 1409 852 1542 857
rect 1649 852 1750 857
rect 1953 852 2238 857
rect 3585 852 3646 857
rect 3673 852 3758 857
rect 1297 847 1414 852
rect 3673 847 3678 852
rect 481 842 566 847
rect 481 837 486 842
rect 233 832 270 837
rect 433 832 486 837
rect 561 837 566 842
rect 609 842 726 847
rect 1433 842 1462 847
rect 1553 842 1942 847
rect 2745 842 2854 847
rect 3257 842 3278 847
rect 3417 842 3574 847
rect 609 837 614 842
rect 561 832 614 837
rect 721 837 726 842
rect 1457 837 1558 842
rect 3569 837 3574 842
rect 3657 842 3678 847
rect 3753 847 3758 852
rect 3857 847 3926 852
rect 3753 842 3862 847
rect 3921 842 4014 847
rect 4185 842 4262 847
rect 3657 837 3662 842
rect 4185 837 4190 842
rect 721 832 806 837
rect 801 827 806 832
rect 905 832 1294 837
rect 905 827 910 832
rect 1289 827 1294 832
rect 1409 832 1438 837
rect 1577 832 1646 837
rect 1665 832 1854 837
rect 1953 832 2078 837
rect 2329 832 2374 837
rect 2433 832 2494 837
rect 2625 832 2742 837
rect 3185 832 3278 837
rect 3569 832 3662 837
rect 3689 832 3742 837
rect 3873 832 3910 837
rect 4081 832 4190 837
rect 4257 837 4262 842
rect 4305 842 4414 847
rect 4513 842 4598 847
rect 4305 837 4310 842
rect 4513 837 4518 842
rect 4257 832 4310 837
rect 4329 832 4518 837
rect 4593 837 4598 842
rect 4593 832 4638 837
rect 1409 827 1414 832
rect 1849 827 1958 832
rect 2833 827 2918 832
rect 129 822 174 827
rect 201 822 246 827
rect 497 822 542 827
rect 553 822 606 827
rect 649 822 750 827
rect 801 822 910 827
rect 1081 822 1126 827
rect 1289 822 1414 827
rect 1545 822 1590 827
rect 1785 822 1830 827
rect 2009 822 2038 827
rect 2577 822 2630 827
rect 2697 822 2750 827
rect 2809 822 2838 827
rect 2913 822 2982 827
rect 3057 822 3118 827
rect 3193 822 3358 827
rect 3377 822 3470 827
rect 3689 822 3734 827
rect 3889 822 3966 827
rect 4025 822 4102 827
rect 4201 822 4254 827
rect 4345 822 4422 827
rect 4529 822 4566 827
rect 3377 817 3382 822
rect 233 812 254 817
rect 369 812 422 817
rect 417 807 422 812
rect 505 812 646 817
rect 657 812 1030 817
rect 1065 812 1134 817
rect 1737 812 1806 817
rect 1929 812 2022 817
rect 2305 812 2382 817
rect 2857 812 2902 817
rect 3049 812 3382 817
rect 3465 817 3470 822
rect 3465 812 3494 817
rect 3529 812 3550 817
rect 3713 812 4070 817
rect 505 807 510 812
rect 1025 807 1030 812
rect 3649 807 3718 812
rect 4065 807 4070 812
rect 4169 812 4198 817
rect 4249 812 4310 817
rect 4537 812 4582 817
rect 4169 807 4174 812
rect 257 802 326 807
rect 417 802 510 807
rect 529 802 798 807
rect 809 802 1014 807
rect 1025 802 1270 807
rect 1905 802 1982 807
rect 2209 802 2294 807
rect 2393 802 2510 807
rect 3217 802 3654 807
rect 3945 802 4046 807
rect 4065 802 4174 807
rect 4449 802 4654 807
rect 2289 797 2398 802
rect 161 792 230 797
rect 633 792 726 797
rect 777 792 846 797
rect 889 792 918 797
rect 1041 792 1070 797
rect 1257 792 1286 797
rect 1497 792 1534 797
rect 2945 792 3030 797
rect 3201 792 3318 797
rect 3329 792 3390 797
rect 3513 792 3534 797
rect 3665 792 3694 797
rect 3785 792 3870 797
rect 3897 792 3926 797
rect 4305 792 4358 797
rect 4441 792 4486 797
rect 4617 792 4646 797
rect 913 787 1046 792
rect 681 782 806 787
rect 833 782 862 787
rect 1233 782 1286 787
rect 1625 782 1654 787
rect 2193 782 2326 787
rect 2321 777 2326 782
rect 2521 782 2558 787
rect 2729 782 2838 787
rect 2849 782 2934 787
rect 2521 777 2526 782
rect 273 772 454 777
rect 745 772 782 777
rect 881 772 1014 777
rect 1273 772 1334 777
rect 1505 772 1542 777
rect 2321 772 2526 777
rect 2929 777 2934 782
rect 3017 782 3054 787
rect 3089 782 3182 787
rect 3297 782 3358 787
rect 3817 782 3838 787
rect 3857 782 3910 787
rect 4297 782 4326 787
rect 4337 782 4406 787
rect 4473 782 4542 787
rect 4617 782 4678 787
rect 3017 777 3022 782
rect 3089 777 3094 782
rect 2929 772 3022 777
rect 3065 772 3094 777
rect 3177 777 3182 782
rect 3177 772 3246 777
rect 273 757 278 772
rect 449 757 454 772
rect 881 767 886 772
rect 473 762 638 767
rect 785 762 886 767
rect 1009 767 1014 772
rect 1009 762 1038 767
rect 1121 762 1214 767
rect 1241 762 1262 767
rect 3041 762 3230 767
rect 3305 762 3422 767
rect 4281 762 4334 767
rect 1121 757 1126 762
rect 249 752 278 757
rect 313 752 430 757
rect 449 752 734 757
rect 313 747 318 752
rect 241 742 318 747
rect 425 747 430 752
rect 729 747 734 752
rect 801 752 1014 757
rect 1097 752 1126 757
rect 1209 757 1214 762
rect 1209 752 1382 757
rect 1625 752 1742 757
rect 1841 752 1894 757
rect 3041 752 3126 757
rect 801 747 806 752
rect 425 742 454 747
rect 545 742 590 747
rect 729 742 806 747
rect 825 742 870 747
rect 1049 742 1078 747
rect 1137 742 1246 747
rect 1073 737 1142 742
rect 1241 737 1246 742
rect 1393 742 1694 747
rect 1729 742 1902 747
rect 2097 742 2174 747
rect 2225 742 2278 747
rect 2417 742 2470 747
rect 2545 742 2606 747
rect 2761 742 2830 747
rect 2993 742 3350 747
rect 3737 742 3790 747
rect 4257 742 4302 747
rect 4465 742 4518 747
rect 4569 742 4686 747
rect 1393 737 1398 742
rect 2761 737 2766 742
rect 169 732 262 737
rect 329 732 526 737
rect 577 732 662 737
rect 905 732 942 737
rect 1241 732 1398 737
rect 1649 732 1710 737
rect 2345 732 2438 737
rect 2577 732 2622 737
rect 2705 732 2766 737
rect 2825 737 2830 742
rect 2825 732 2854 737
rect 3697 732 3894 737
rect 4081 732 4190 737
rect 3145 727 3286 732
rect 4209 727 4214 737
rect 4225 732 4270 737
rect 4633 732 4670 737
rect 841 722 878 727
rect 1185 722 1222 727
rect 1985 722 2078 727
rect 2145 722 2278 727
rect 2849 722 2894 727
rect 2969 722 3014 727
rect 3121 722 3150 727
rect 3281 722 3310 727
rect 3777 722 3846 727
rect 4193 722 4214 727
rect 4289 722 4366 727
rect 4417 722 4486 727
rect 4601 722 4678 727
rect 1985 717 1990 722
rect 137 712 182 717
rect 345 712 390 717
rect 441 712 470 717
rect 521 712 814 717
rect 857 712 910 717
rect 1049 712 1078 717
rect 1289 712 1334 717
rect 1609 712 1646 717
rect 1681 712 1710 717
rect 1753 712 1774 717
rect 1881 712 1942 717
rect 1961 712 1990 717
rect 2073 717 2078 722
rect 3121 717 3126 722
rect 2073 712 2174 717
rect 2249 712 2294 717
rect 2401 712 2486 717
rect 2585 712 2694 717
rect 2689 707 2694 712
rect 2777 712 2806 717
rect 2865 712 3126 717
rect 3145 712 3190 717
rect 3241 712 3286 717
rect 3409 712 3518 717
rect 3649 712 3894 717
rect 4185 712 4598 717
rect 4705 712 4758 717
rect 2777 707 2782 712
rect 377 702 462 707
rect 457 687 462 702
rect 649 702 678 707
rect 825 702 862 707
rect 2689 702 2782 707
rect 2977 702 3022 707
rect 3593 702 3678 707
rect 3745 702 3910 707
rect 4169 702 4198 707
rect 649 687 654 702
rect 4193 697 4198 702
rect 4273 702 4526 707
rect 4273 697 4278 702
rect 833 692 862 697
rect 217 682 310 687
rect 457 682 654 687
rect 857 687 862 692
rect 921 692 1726 697
rect 921 687 926 692
rect 857 682 926 687
rect 1721 687 1726 692
rect 1785 692 1990 697
rect 1785 687 1790 692
rect 1721 682 1790 687
rect 1913 682 1966 687
rect 1985 677 1990 692
rect 2185 692 2302 697
rect 2609 692 2630 697
rect 2873 692 2902 697
rect 2185 677 2190 692
rect 2897 687 2902 692
rect 3233 692 3262 697
rect 3577 692 3766 697
rect 3825 692 3918 697
rect 4193 692 4278 697
rect 3233 687 3238 692
rect 2897 682 3238 687
rect 3681 682 3814 687
rect 3809 677 3814 682
rect 3929 682 3982 687
rect 3929 677 3934 682
rect 1985 672 2190 677
rect 3265 672 3454 677
rect 3809 672 3934 677
rect 1169 662 1278 667
rect 1169 657 1174 662
rect 257 652 406 657
rect 1057 652 1174 657
rect 1273 657 1278 662
rect 1433 662 1702 667
rect 1273 652 1302 657
rect 257 637 262 652
rect 233 632 262 637
rect 401 637 406 652
rect 1433 647 1438 662
rect 1697 647 1702 662
rect 3153 652 3246 657
rect 3153 647 3158 652
rect 1185 642 1270 647
rect 1377 642 1438 647
rect 1561 642 1638 647
rect 1697 642 1726 647
rect 2529 642 2662 647
rect 3041 642 3158 647
rect 3241 647 3246 652
rect 3985 652 4102 657
rect 3985 647 3990 652
rect 3241 642 3358 647
rect 3961 642 3990 647
rect 4097 647 4102 652
rect 4097 642 4190 647
rect 1561 637 1566 642
rect 401 632 430 637
rect 481 632 638 637
rect 849 632 894 637
rect 481 627 486 632
rect 201 622 238 627
rect 289 622 366 627
rect 417 622 486 627
rect 633 627 638 632
rect 1233 627 1238 637
rect 1417 632 1566 637
rect 1633 637 1638 642
rect 1633 632 1814 637
rect 2737 632 2870 637
rect 3097 632 3182 637
rect 3273 632 3454 637
rect 3673 632 3846 637
rect 3905 632 4214 637
rect 633 622 662 627
rect 673 622 718 627
rect 881 622 958 627
rect 1153 622 1262 627
rect 1353 622 1406 627
rect 1577 622 1622 627
rect 1689 622 1718 627
rect 1753 622 1822 627
rect 2265 622 2310 627
rect 2521 622 2566 627
rect 3137 622 3286 627
rect 3521 622 3590 627
rect 3609 622 3654 627
rect 3521 617 3526 622
rect 193 612 318 617
rect 345 612 398 617
rect 625 612 766 617
rect 1073 612 1102 617
rect 1201 612 1238 617
rect 1345 612 1398 617
rect 1425 612 1542 617
rect 1561 612 1638 617
rect 1745 612 1806 617
rect 2033 612 2054 617
rect 2513 612 2622 617
rect 3009 612 3182 617
rect 3497 612 3526 617
rect 3585 617 3590 622
rect 3673 617 3678 632
rect 3585 612 3678 617
rect 3841 617 3846 632
rect 3889 622 4070 627
rect 4065 617 4070 622
rect 4185 622 4286 627
rect 4537 622 4606 627
rect 4185 617 4190 622
rect 3841 612 3870 617
rect 3985 612 4030 617
rect 4065 612 4190 617
rect 4585 612 4742 617
rect 417 607 558 612
rect 1425 607 1430 612
rect 233 602 422 607
rect 553 602 790 607
rect 1057 602 1430 607
rect 1537 607 1542 612
rect 1537 602 1694 607
rect 161 592 206 597
rect 337 592 414 597
rect 433 592 574 597
rect 601 592 654 597
rect 1113 592 1350 597
rect 1369 592 1574 597
rect 1729 592 1766 597
rect 1825 592 2014 597
rect 2033 592 2038 612
rect 3865 607 3990 612
rect 3409 602 3566 607
rect 3577 602 3830 607
rect 4681 602 4750 607
rect 2049 592 2078 597
rect 2417 592 2534 597
rect 3129 592 3166 597
rect 3633 592 3710 597
rect 3881 592 3926 597
rect 4105 592 4150 597
rect 4185 592 4342 597
rect 4553 592 4710 597
rect 1825 587 1830 592
rect 537 582 694 587
rect 713 582 942 587
rect 961 582 1014 587
rect 1057 582 1150 587
rect 1169 582 1238 587
rect 449 577 518 582
rect 713 577 718 582
rect 233 572 454 577
rect 513 572 718 577
rect 937 577 942 582
rect 1233 577 1238 582
rect 1337 582 1422 587
rect 1449 582 1478 587
rect 1505 582 1694 587
rect 1801 582 1830 587
rect 2009 587 2014 592
rect 2009 582 2222 587
rect 3113 582 3142 587
rect 3585 582 3662 587
rect 3913 582 3990 587
rect 4033 582 4118 587
rect 4649 582 4694 587
rect 1337 577 1342 582
rect 1689 577 1806 582
rect 937 572 1022 577
rect 1233 572 1342 577
rect 1361 572 1494 577
rect 1041 567 1190 572
rect 1489 567 1494 572
rect 1561 572 1590 577
rect 1953 572 2030 577
rect 2769 572 2854 577
rect 3481 572 3574 577
rect 1561 567 1566 572
rect 2769 567 2774 572
rect 465 562 518 567
rect 633 562 1046 567
rect 1185 562 1214 567
rect 1385 562 1462 567
rect 1489 562 1566 567
rect 1721 562 2038 567
rect 2073 562 2126 567
rect 2745 562 2774 567
rect 2849 567 2854 572
rect 3569 567 3574 572
rect 3665 572 3902 577
rect 4129 572 4222 577
rect 4537 572 4558 577
rect 3665 567 3670 572
rect 3897 567 3998 572
rect 4129 567 4134 572
rect 2849 562 2878 567
rect 3201 562 3286 567
rect 3305 562 3430 567
rect 3569 562 3670 567
rect 3993 562 4134 567
rect 513 557 638 562
rect 3201 557 3206 562
rect 121 552 198 557
rect 369 552 494 557
rect 657 552 758 557
rect 769 552 894 557
rect 993 552 1030 557
rect 1065 552 1294 557
rect 1401 552 1470 557
rect 1945 552 2182 557
rect 2905 552 2982 557
rect 3041 552 3206 557
rect 3281 557 3286 562
rect 3281 552 3334 557
rect 3689 552 3974 557
rect 4537 552 4630 557
rect 121 547 126 552
rect 97 542 126 547
rect 193 547 198 552
rect 193 542 222 547
rect 345 542 494 547
rect 617 542 734 547
rect 753 537 758 552
rect 889 547 998 552
rect 4537 547 4542 552
rect 809 542 870 547
rect 1017 542 1046 547
rect 1105 542 1174 547
rect 1201 542 1262 547
rect 1321 542 1478 547
rect 1497 542 1662 547
rect 1681 542 1974 547
rect 2009 542 2102 547
rect 2361 542 2590 547
rect 2673 542 2886 547
rect 3177 542 3310 547
rect 3425 542 3494 547
rect 3625 542 3710 547
rect 3881 542 4038 547
rect 4161 542 4262 547
rect 4289 542 4318 547
rect 4329 542 4414 547
rect 4513 542 4542 547
rect 4625 547 4630 552
rect 4625 542 4654 547
rect 4665 542 4726 547
rect 1105 537 1110 542
rect 1497 537 1502 542
rect 129 532 174 537
rect 209 532 518 537
rect 585 532 670 537
rect 753 532 1110 537
rect 1129 532 1166 537
rect 1337 532 1502 537
rect 1657 537 1662 542
rect 1657 532 1702 537
rect 2081 532 2134 537
rect 3289 532 3390 537
rect 3449 532 3870 537
rect 4049 532 4766 537
rect 1185 527 1318 532
rect 1833 527 1958 532
rect 3865 527 3870 532
rect 3985 527 4054 532
rect 161 522 254 527
rect 393 522 446 527
rect 505 522 982 527
rect 1041 522 1190 527
rect 1313 522 1430 527
rect 1513 522 1694 527
rect 1809 522 1838 527
rect 1953 522 1982 527
rect 2025 522 2046 527
rect 2969 522 3070 527
rect 3865 522 3990 527
rect 4113 522 4182 527
rect 4265 522 4702 527
rect 1425 517 1518 522
rect 4177 517 4270 522
rect 193 512 214 517
rect 241 512 278 517
rect 273 507 278 512
rect 409 512 502 517
rect 641 512 686 517
rect 705 512 734 517
rect 745 512 950 517
rect 409 507 414 512
rect 81 502 254 507
rect 273 502 414 507
rect 433 502 462 507
rect 513 502 630 507
rect 625 497 630 502
rect 705 497 710 512
rect 945 507 950 512
rect 1113 512 1182 517
rect 1241 512 1294 517
rect 1305 512 1406 517
rect 1113 507 1118 512
rect 1401 507 1406 512
rect 1609 512 1638 517
rect 1673 512 1894 517
rect 1905 512 1950 517
rect 2089 512 2134 517
rect 2441 512 2694 517
rect 2857 512 2902 517
rect 3105 512 3206 517
rect 3665 512 3702 517
rect 3721 512 3790 517
rect 4009 512 4054 517
rect 4289 512 4406 517
rect 1609 507 1614 512
rect 1889 507 1894 512
rect 4401 507 4406 512
rect 4521 512 4574 517
rect 4521 507 4526 512
rect 753 502 830 507
rect 841 502 918 507
rect 945 502 1118 507
rect 1281 502 1342 507
rect 1401 502 1614 507
rect 1681 502 1718 507
rect 1889 502 1910 507
rect 3449 502 3542 507
rect 3889 502 4174 507
rect 4169 497 4174 502
rect 4241 502 4270 507
rect 4401 502 4526 507
rect 4569 507 4574 512
rect 4657 512 4686 517
rect 4657 507 4662 512
rect 4569 502 4662 507
rect 4241 497 4246 502
rect 201 492 230 497
rect 497 492 526 497
rect 625 492 710 497
rect 729 492 782 497
rect 857 492 926 497
rect 521 477 526 492
rect 729 477 734 492
rect 921 487 926 492
rect 1137 492 1382 497
rect 3545 492 3734 497
rect 4073 492 4134 497
rect 4169 492 4246 497
rect 1137 487 1142 492
rect 809 482 902 487
rect 921 482 1142 487
rect 1401 482 1662 487
rect 1769 482 1814 487
rect 4121 482 4150 487
rect 4641 482 4790 487
rect 1289 477 1406 482
rect 1657 477 1662 482
rect 521 472 734 477
rect 1265 472 1294 477
rect 1657 472 1710 477
rect 3561 472 3734 477
rect 1161 462 1470 467
rect 1465 457 1470 462
rect 1569 462 1622 467
rect 1569 457 1574 462
rect 625 452 774 457
rect 817 452 934 457
rect 1081 452 1358 457
rect 1465 452 1574 457
rect 481 442 582 447
rect 481 437 486 442
rect 457 432 486 437
rect 577 437 582 442
rect 625 437 630 452
rect 577 432 630 437
rect 769 437 774 452
rect 1617 447 1622 462
rect 1777 462 1806 467
rect 3849 462 3926 467
rect 1777 447 1782 462
rect 3505 457 3590 462
rect 3849 457 3854 462
rect 2057 452 2150 457
rect 3481 452 3510 457
rect 3585 452 3854 457
rect 3921 457 3926 462
rect 3921 452 4518 457
rect 2057 447 2062 452
rect 1217 442 1270 447
rect 1617 442 1782 447
rect 1993 442 2022 447
rect 2033 442 2062 447
rect 2145 447 2150 452
rect 2145 442 2334 447
rect 2801 442 2854 447
rect 2945 442 3014 447
rect 3393 442 3574 447
rect 2945 437 2950 442
rect 769 432 862 437
rect 857 427 862 432
rect 945 432 966 437
rect 1257 432 1438 437
rect 1937 432 2030 437
rect 2833 432 2950 437
rect 3009 437 3014 442
rect 3009 432 3046 437
rect 3097 432 3262 437
rect 3473 432 3550 437
rect 945 427 950 432
rect 185 422 366 427
rect 385 422 454 427
rect 489 422 534 427
rect 729 422 766 427
rect 793 422 838 427
rect 857 422 950 427
rect 961 427 966 432
rect 3569 427 3574 442
rect 3865 442 3910 447
rect 3865 427 3870 442
rect 4457 432 4566 437
rect 961 422 1166 427
rect 1249 422 1318 427
rect 1337 422 1382 427
rect 1401 422 1494 427
rect 1529 422 1574 427
rect 1681 422 1790 427
rect 1801 422 1998 427
rect 2009 422 2038 427
rect 2089 422 2134 427
rect 2641 422 2766 427
rect 2897 422 2998 427
rect 3081 422 3142 427
rect 3209 422 3318 427
rect 3569 422 3870 427
rect 4169 422 4454 427
rect 385 417 390 422
rect 2641 417 2646 422
rect 177 412 198 417
rect 297 412 326 417
rect 361 412 390 417
rect 433 412 582 417
rect 633 412 726 417
rect 801 412 838 417
rect 1057 412 1086 417
rect 1305 412 1334 417
rect 1329 407 1334 412
rect 1457 412 1550 417
rect 2457 412 2646 417
rect 2761 417 2766 422
rect 4449 417 4454 422
rect 4561 422 4686 427
rect 4729 422 4750 427
rect 4561 417 4566 422
rect 2761 412 2926 417
rect 3329 412 3454 417
rect 4225 412 4254 417
rect 4449 412 4566 417
rect 1457 407 1462 412
rect 4137 407 4206 412
rect 4273 407 4374 412
rect 4609 407 4614 417
rect 529 402 558 407
rect 1041 402 1070 407
rect 1065 397 1070 402
rect 1129 402 1222 407
rect 1329 402 1462 407
rect 2761 402 2830 407
rect 1129 397 1134 402
rect 2825 397 2830 402
rect 2913 402 2966 407
rect 3377 402 3446 407
rect 3889 402 4006 407
rect 4025 402 4142 407
rect 4201 402 4278 407
rect 4369 402 4430 407
rect 4609 402 4686 407
rect 2913 397 2918 402
rect 3889 397 3894 402
rect 81 392 302 397
rect 873 392 990 397
rect 1065 392 1134 397
rect 1153 392 1270 397
rect 1689 392 1734 397
rect 2137 392 2182 397
rect 2313 392 2374 397
rect 2577 392 2806 397
rect 2825 392 2918 397
rect 3337 392 3366 397
rect 3457 392 3518 397
rect 3609 392 3710 397
rect 3729 392 3894 397
rect 4001 397 4006 402
rect 4001 392 4030 397
rect 4153 392 4230 397
rect 4273 392 4358 397
rect 4433 392 4502 397
rect 4561 392 4606 397
rect 4673 392 4734 397
rect 249 382 510 387
rect 1161 382 1206 387
rect 1721 382 2102 387
rect 2305 382 2342 387
rect 2577 382 2646 387
rect 3545 382 3630 387
rect 3681 382 3726 387
rect 3905 382 4070 387
rect 4329 382 4382 387
rect 4393 382 4454 387
rect 4473 382 4726 387
rect 3745 377 3910 382
rect 529 372 750 377
rect 529 357 534 372
rect 745 357 750 372
rect 1521 372 1598 377
rect 2249 372 2318 377
rect 2937 372 3230 377
rect 3329 372 3486 377
rect 3513 372 3750 377
rect 3921 372 4006 377
rect 1521 367 1526 372
rect 769 362 1006 367
rect 1225 362 1366 367
rect 1497 362 1526 367
rect 1593 367 1598 372
rect 3329 367 3334 372
rect 1593 362 1622 367
rect 2753 362 2910 367
rect 3081 362 3110 367
rect 3241 362 3334 367
rect 3481 367 3486 372
rect 4001 367 4006 372
rect 4081 372 4438 377
rect 4609 372 4670 377
rect 4713 372 4750 377
rect 4081 367 4086 372
rect 3481 362 3678 367
rect 1225 357 1230 362
rect 393 352 534 357
rect 649 352 726 357
rect 745 352 798 357
rect 1017 352 1230 357
rect 1361 357 1366 362
rect 1361 352 1486 357
rect 1633 352 1750 357
rect 2665 352 2710 357
rect 649 347 654 352
rect 177 342 414 347
rect 545 342 654 347
rect 721 347 726 352
rect 1481 347 1486 352
rect 1561 347 1638 352
rect 2753 347 2758 362
rect 721 342 750 347
rect 817 342 894 347
rect 1241 342 1350 347
rect 1481 342 1566 347
rect 1841 342 1974 347
rect 2105 342 2462 347
rect 2489 342 2646 347
rect 2729 342 2758 347
rect 2905 347 2910 362
rect 3105 357 3246 362
rect 3673 357 3678 362
rect 3737 362 3982 367
rect 4001 362 4086 367
rect 4273 362 4326 367
rect 3737 357 3742 362
rect 3345 352 3470 357
rect 3673 352 3742 357
rect 3889 352 3982 357
rect 4425 352 4470 357
rect 2905 342 3030 347
rect 3041 342 3142 347
rect 2489 337 2494 342
rect 129 332 174 337
rect 441 332 806 337
rect 905 332 974 337
rect 1585 332 1806 337
rect 1977 332 2094 337
rect 801 327 910 332
rect 2089 327 2094 332
rect 2193 332 2222 337
rect 2465 332 2494 337
rect 2641 337 2646 342
rect 3137 337 3142 342
rect 3233 342 3262 347
rect 3401 342 3526 347
rect 3569 342 3654 347
rect 3817 342 3910 347
rect 3945 342 4038 347
rect 4161 342 4230 347
rect 4361 342 4462 347
rect 3233 337 3238 342
rect 2641 332 2702 337
rect 2193 327 2198 332
rect 465 322 662 327
rect 1121 322 1182 327
rect 1321 322 1390 327
rect 1993 322 2038 327
rect 2089 322 2198 327
rect 2697 327 2702 332
rect 2769 332 2822 337
rect 2841 332 2894 337
rect 3137 332 3238 337
rect 3353 332 3462 337
rect 3657 332 3694 337
rect 3833 332 3918 337
rect 3929 332 3958 337
rect 4025 332 4174 337
rect 4697 332 4742 337
rect 2769 327 2774 332
rect 2697 322 2774 327
rect 2817 317 2822 332
rect 3017 322 3118 327
rect 3281 322 3398 327
rect 4073 322 4182 327
rect 4201 322 4350 327
rect 3017 317 3022 322
rect 3641 317 3734 322
rect 4345 317 4350 322
rect 4473 322 4582 327
rect 4473 317 4478 322
rect 297 312 342 317
rect 513 312 558 317
rect 577 312 694 317
rect 689 307 694 312
rect 833 312 870 317
rect 881 312 910 317
rect 1225 312 1294 317
rect 1329 312 1366 317
rect 1377 312 1454 317
rect 1473 312 1518 317
rect 1569 312 1790 317
rect 1905 312 1950 317
rect 2409 312 2478 317
rect 2489 312 2574 317
rect 2625 312 2662 317
rect 2817 312 3022 317
rect 3257 312 3294 317
rect 3361 312 3430 317
rect 3441 312 3646 317
rect 3729 312 3822 317
rect 833 307 838 312
rect 3817 307 3822 312
rect 3929 312 3990 317
rect 4001 312 4038 317
rect 4153 312 4182 317
rect 3929 307 3934 312
rect 329 302 358 307
rect 689 302 838 307
rect 1081 302 1430 307
rect 1769 302 1798 307
rect 3041 302 3198 307
rect 3273 302 3358 307
rect 3385 302 3486 307
rect 3657 302 3718 307
rect 3817 302 3934 307
rect 3985 307 3990 312
rect 4177 307 4182 312
rect 4241 312 4294 317
rect 4345 312 4478 317
rect 4241 307 4246 312
rect 3985 302 4086 307
rect 4177 302 4246 307
rect 1425 297 1614 302
rect 377 292 494 297
rect 1209 292 1278 297
rect 1345 292 1406 297
rect 377 287 382 292
rect 305 282 382 287
rect 489 287 494 292
rect 1609 287 1614 297
rect 1769 287 1774 302
rect 3153 292 3262 297
rect 3257 287 3262 292
rect 3409 292 3558 297
rect 3409 287 3414 292
rect 489 282 534 287
rect 553 282 670 287
rect 857 282 1198 287
rect 1289 282 1582 287
rect 1609 282 1774 287
rect 2281 282 2310 287
rect 2713 282 2878 287
rect 3105 282 3142 287
rect 3257 282 3414 287
rect 3465 282 3494 287
rect 4265 282 4326 287
rect 553 277 558 282
rect 1 272 294 277
rect 377 272 558 277
rect 665 277 670 282
rect 1193 277 1294 282
rect 665 272 694 277
rect 713 272 838 277
rect 1857 272 1974 277
rect 289 267 382 272
rect 713 267 718 272
rect 833 267 934 272
rect 1313 267 1566 272
rect 401 262 718 267
rect 929 262 958 267
rect 1065 262 1214 267
rect 1289 262 1318 267
rect 1561 262 1590 267
rect 1065 257 1070 262
rect 217 252 582 257
rect 689 252 1070 257
rect 1209 257 1214 262
rect 1857 257 1862 272
rect 1969 267 1974 272
rect 3137 267 3142 282
rect 3465 267 3470 282
rect 1969 262 2150 267
rect 3137 262 3470 267
rect 4065 262 4246 267
rect 4065 257 4070 262
rect 1209 252 1238 257
rect 1249 252 1862 257
rect 1873 252 1958 257
rect 3705 252 4070 257
rect 4241 257 4246 262
rect 4241 252 4550 257
rect 1249 247 1254 252
rect 337 242 382 247
rect 393 242 486 247
rect 593 242 766 247
rect 865 242 1254 247
rect 1273 242 1310 247
rect 1409 242 1574 247
rect 3033 242 3086 247
rect 4105 242 4222 247
rect 481 237 598 242
rect 1305 237 1414 242
rect 1641 237 1886 242
rect 4105 237 4110 242
rect 161 232 462 237
rect 881 232 1286 237
rect 1433 232 1526 237
rect 1617 232 1646 237
rect 1881 232 1910 237
rect 1929 232 1982 237
rect 2473 232 2526 237
rect 2561 232 2622 237
rect 2921 232 3086 237
rect 3417 232 3470 237
rect 3633 232 3678 237
rect 3961 232 4038 237
rect 4081 232 4110 237
rect 4217 237 4222 242
rect 4217 232 4270 237
rect 1617 227 1622 232
rect 2809 227 2894 232
rect 3961 227 3966 232
rect 129 222 174 227
rect 185 222 230 227
rect 297 222 342 227
rect 361 222 470 227
rect 545 222 670 227
rect 849 222 1070 227
rect 1065 217 1070 222
rect 1193 222 1222 227
rect 1401 222 1470 227
rect 1513 222 1622 227
rect 1673 222 1734 227
rect 1769 222 1902 227
rect 1929 222 1990 227
rect 2321 222 2414 227
rect 2457 222 2606 227
rect 2633 222 2726 227
rect 2753 222 2814 227
rect 2889 222 2918 227
rect 3145 222 3262 227
rect 3473 222 3526 227
rect 3537 222 3654 227
rect 3665 222 3862 227
rect 3937 222 3966 227
rect 4033 227 4038 232
rect 4033 222 4062 227
rect 4121 222 4230 227
rect 4249 222 4286 227
rect 4305 222 4606 227
rect 4705 222 4734 227
rect 1193 217 1198 222
rect 289 212 390 217
rect 649 212 758 217
rect 809 212 1046 217
rect 1065 212 1198 217
rect 1233 212 1462 217
rect 1609 212 1814 217
rect 1913 212 1998 217
rect 2481 212 2566 217
rect 2825 212 2854 217
rect 3377 212 3414 217
rect 3857 212 4078 217
rect 4137 212 4206 217
rect 409 202 782 207
rect 897 202 1006 207
rect 1041 202 1046 212
rect 1457 207 1462 212
rect 3665 207 3774 212
rect 4305 207 4310 222
rect 1457 202 1654 207
rect 1665 202 1750 207
rect 1857 202 1966 207
rect 2017 202 2102 207
rect 3257 202 3670 207
rect 3769 202 4310 207
rect 4601 207 4606 222
rect 4601 202 4782 207
rect 1649 197 1654 202
rect 2017 197 2022 202
rect 81 192 150 197
rect 217 192 254 197
rect 273 192 342 197
rect 377 192 430 197
rect 649 192 718 197
rect 729 192 790 197
rect 841 192 886 197
rect 225 182 254 187
rect 249 177 254 182
rect 393 182 422 187
rect 769 182 830 187
rect 393 177 398 182
rect 881 177 886 192
rect 1009 192 1038 197
rect 1153 192 1190 197
rect 1281 192 1470 197
rect 1561 192 1630 197
rect 1649 192 1846 197
rect 1897 192 1950 197
rect 1985 192 2022 197
rect 2097 197 2102 202
rect 2097 192 2126 197
rect 2145 192 2238 197
rect 2521 192 2566 197
rect 2617 192 2646 197
rect 2777 192 2822 197
rect 3065 192 3238 197
rect 3409 192 3446 197
rect 3681 192 3710 197
rect 3721 192 3758 197
rect 3905 192 3998 197
rect 4009 192 4054 197
rect 4089 192 4166 197
rect 4281 192 4590 197
rect 1009 177 1014 192
rect 1841 187 1846 192
rect 2145 187 2150 192
rect 1369 182 1406 187
rect 1401 177 1406 182
rect 1465 182 1494 187
rect 1601 182 1630 187
rect 1465 177 1470 182
rect 249 172 398 177
rect 529 172 774 177
rect 881 172 1014 177
rect 1345 172 1382 177
rect 1401 172 1470 177
rect 1625 177 1630 182
rect 1801 182 1830 187
rect 1841 182 1870 187
rect 1977 182 2150 187
rect 2233 187 2238 192
rect 2233 182 2342 187
rect 2505 182 2534 187
rect 2769 182 2942 187
rect 3441 182 3734 187
rect 3809 182 4110 187
rect 1801 177 1806 182
rect 1865 177 1982 182
rect 1625 172 1806 177
rect 2065 172 2086 177
rect 3433 172 3462 177
rect 3937 172 4694 177
rect 3457 167 3462 172
rect 3753 167 3942 172
rect 1905 162 1934 167
rect 1929 157 1934 162
rect 2073 162 2222 167
rect 2665 162 2750 167
rect 3457 162 3758 167
rect 2073 157 2078 162
rect 2665 157 2670 162
rect 1929 152 2078 157
rect 2641 152 2670 157
rect 2745 157 2750 162
rect 3961 157 4142 162
rect 2745 152 2782 157
rect 2905 152 3054 157
rect 3329 152 3366 157
rect 3873 152 3966 157
rect 4137 152 4318 157
rect 313 142 510 147
rect 569 142 686 147
rect 801 142 846 147
rect 937 142 982 147
rect 1137 142 1190 147
rect 1601 142 1878 147
rect 2097 142 2390 147
rect 2577 142 2662 147
rect 2705 142 2774 147
rect 2841 142 2902 147
rect 3369 142 3398 147
rect 3465 142 3494 147
rect 3513 142 3630 147
rect 3777 142 4142 147
rect 4425 142 4710 147
rect 841 132 902 137
rect 2633 132 2806 137
rect 2865 132 2990 137
rect 3673 132 3718 137
rect 4017 132 4118 137
rect 1153 122 1222 127
rect 1985 122 2062 127
rect 2657 122 2686 127
rect 2681 117 2686 122
rect 2777 122 2894 127
rect 2777 117 2782 122
rect 2889 117 2894 122
rect 3001 122 3038 127
rect 3001 117 3006 122
rect 193 112 238 117
rect 297 112 342 117
rect 553 112 598 117
rect 745 112 838 117
rect 849 112 894 117
rect 1105 112 1150 117
rect 1201 112 1270 117
rect 1289 112 1334 117
rect 1577 112 1622 117
rect 2001 112 2054 117
rect 2137 112 2166 117
rect 2681 112 2782 117
rect 2801 112 2870 117
rect 2889 112 3006 117
rect 3161 112 3262 117
rect 3401 112 3422 117
rect 3489 112 3662 117
rect 833 107 838 112
rect 3657 107 3662 112
rect 3729 112 3782 117
rect 3817 112 3870 117
rect 4017 112 4086 117
rect 4681 112 4734 117
rect 3729 107 3734 112
rect 833 102 862 107
rect 1257 102 1302 107
rect 2073 102 2110 107
rect 2249 102 2286 107
rect 3361 102 3414 107
rect 3657 102 3734 107
rect 793 92 822 97
rect 817 87 822 92
rect 905 92 1190 97
rect 905 87 910 92
rect 817 82 910 87
rect 1185 77 1190 92
rect 1345 92 1518 97
rect 2153 92 2182 97
rect 2273 92 2302 97
rect 1345 77 1350 92
rect 2089 82 2206 87
rect 1185 72 1350 77
rect 2017 32 2310 37
rect 2057 12 2086 17
rect 2081 7 2086 12
rect 2297 12 2326 17
rect 2361 12 2670 17
rect 2297 7 2302 12
rect 2081 2 2302 7
use M3_M2  M3_M2_0
timestamp 1677677812
transform 1 0 1652 0 1 4735
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1677677812
transform 1 0 3124 0 1 4735
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_0
timestamp 1677677812
transform 1 0 24 0 1 4717
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_2
timestamp 1677677812
transform 1 0 48 0 1 4693
box -10 -10 10 10
use M3_M2  M3_M2_2
timestamp 1677677812
transform 1 0 1172 0 1 4705
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1677677812
transform 1 0 2796 0 1 4705
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_1
timestamp 1677677812
transform 1 0 4843 0 1 4717
box -10 -10 10 10
use M3_M2  M3_M2_4
timestamp 1677677812
transform 1 0 2020 0 1 4685
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1677677812
transform 1 0 2476 0 1 4685
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_3
timestamp 1677677812
transform 1 0 4819 0 1 4693
box -10 -10 10 10
use top_level_VIA0  top_level_VIA0_0
timestamp 1677677812
transform 1 0 24 0 1 4670
box -10 -3 10 3
use M2_M1  M2_M1_1
timestamp 1677677812
transform 1 0 124 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1677677812
transform 1 0 92 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_57
timestamp 1677677812
transform 1 0 92 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_77
timestamp 1677677812
transform 1 0 180 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_2
timestamp 1677677812
transform 1 0 268 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_3
timestamp 1677677812
transform 1 0 316 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1677677812
transform 1 0 348 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_58
timestamp 1677677812
transform 1 0 324 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_59
timestamp 1677677812
transform 1 0 348 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_37
timestamp 1677677812
transform 1 0 380 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_4
timestamp 1677677812
transform 1 0 428 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1677677812
transform 1 0 404 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_38
timestamp 1677677812
transform 1 0 428 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1677677812
transform 1 0 404 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1677677812
transform 1 0 492 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_14
timestamp 1677677812
transform 1 0 548 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1677677812
transform 1 0 588 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_6
timestamp 1677677812
transform 1 0 548 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1677677812
transform 1 0 556 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_8
timestamp 1677677812
transform 1 0 588 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1677677812
transform 1 0 540 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_81
timestamp 1677677812
transform 1 0 636 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_61
timestamp 1677677812
transform 1 0 636 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_82
timestamp 1677677812
transform 1 0 652 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_16
timestamp 1677677812
transform 1 0 692 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1677677812
transform 1 0 732 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1677677812
transform 1 0 692 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_10
timestamp 1677677812
transform 1 0 732 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_11
timestamp 1677677812
transform 1 0 788 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1677677812
transform 1 0 708 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_62
timestamp 1677677812
transform 1 0 708 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_12
timestamp 1677677812
transform 1 0 860 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_84
timestamp 1677677812
transform 1 0 812 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_39
timestamp 1677677812
transform 1 0 860 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1677677812
transform 1 0 884 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_63
timestamp 1677677812
transform 1 0 812 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1677677812
transform 1 0 940 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_18
timestamp 1677677812
transform 1 0 1028 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_19
timestamp 1677677812
transform 1 0 1068 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_14
timestamp 1677677812
transform 1 0 1028 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_15
timestamp 1677677812
transform 1 0 1036 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_16
timestamp 1677677812
transform 1 0 1068 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_85
timestamp 1677677812
transform 1 0 1020 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1677677812
transform 1 0 1116 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_64
timestamp 1677677812
transform 1 0 1116 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_17
timestamp 1677677812
transform 1 0 1164 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1677677812
transform 1 0 1228 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1677677812
transform 1 0 1260 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_65
timestamp 1677677812
transform 1 0 1260 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_19
timestamp 1677677812
transform 1 0 1316 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_20
timestamp 1677677812
transform 1 0 1372 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_41
timestamp 1677677812
transform 1 0 1372 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_88
timestamp 1677677812
transform 1 0 1396 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_66
timestamp 1677677812
transform 1 0 1348 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_67
timestamp 1677677812
transform 1 0 1396 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1677677812
transform 1 0 1420 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_42
timestamp 1677677812
transform 1 0 1444 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_22
timestamp 1677677812
transform 1 0 1508 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1677677812
transform 1 0 1532 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_68
timestamp 1677677812
transform 1 0 1532 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_69
timestamp 1677677812
transform 1 0 1548 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1677677812
transform 1 0 1572 0 1 4645
box -3 -3 3 3
use M2_M1  M2_M1_23
timestamp 1677677812
transform 1 0 1620 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_90
timestamp 1677677812
transform 1 0 1588 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_70
timestamp 1677677812
transform 1 0 1588 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_24
timestamp 1677677812
transform 1 0 1676 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_6
timestamp 1677677812
transform 1 0 1868 0 1 4675
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1677677812
transform 1 0 1804 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1677677812
transform 1 0 1844 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_25
timestamp 1677677812
transform 1 0 1804 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1677677812
transform 1 0 1844 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1677677812
transform 1 0 1900 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1677677812
transform 1 0 1796 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_71
timestamp 1677677812
transform 1 0 1796 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_92
timestamp 1677677812
transform 1 0 1820 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_72
timestamp 1677677812
transform 1 0 1844 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1677677812
transform 1 0 1820 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_28
timestamp 1677677812
transform 1 0 1956 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1677677812
transform 1 0 1932 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_97
timestamp 1677677812
transform 1 0 1932 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_29
timestamp 1677677812
transform 1 0 2036 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_30
timestamp 1677677812
transform 1 0 2076 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_94
timestamp 1677677812
transform 1 0 2052 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_98
timestamp 1677677812
transform 1 0 2052 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_31
timestamp 1677677812
transform 1 0 2140 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_22
timestamp 1677677812
transform 1 0 2172 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1677677812
transform 1 0 2212 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_32
timestamp 1677677812
transform 1 0 2172 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_33
timestamp 1677677812
transform 1 0 2212 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1677677812
transform 1 0 2268 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1677677812
transform 1 0 2164 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_96
timestamp 1677677812
transform 1 0 2188 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_73
timestamp 1677677812
transform 1 0 2188 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_35
timestamp 1677677812
transform 1 0 2300 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1677677812
transform 1 0 2340 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_74
timestamp 1677677812
transform 1 0 2292 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_97
timestamp 1677677812
transform 1 0 2380 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_75
timestamp 1677677812
transform 1 0 2380 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_37
timestamp 1677677812
transform 1 0 2412 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1677677812
transform 1 0 2468 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1677677812
transform 1 0 2500 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1677677812
transform 1 0 2500 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1677677812
transform 1 0 2540 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1677677812
transform 1 0 2580 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_39
timestamp 1677677812
transform 1 0 2540 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1677677812
transform 1 0 2580 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_41
timestamp 1677677812
transform 1 0 2636 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1677677812
transform 1 0 2532 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_100
timestamp 1677677812
transform 1 0 2556 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_77
timestamp 1677677812
transform 1 0 2556 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_101
timestamp 1677677812
transform 1 0 2652 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_26
timestamp 1677677812
transform 1 0 2676 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_42
timestamp 1677677812
transform 1 0 2676 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_27
timestamp 1677677812
transform 1 0 2716 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1677677812
transform 1 0 2716 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1677677812
transform 1 0 2692 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_78
timestamp 1677677812
transform 1 0 2692 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1677677812
transform 1 0 2732 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_103
timestamp 1677677812
transform 1 0 2780 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_44
timestamp 1677677812
transform 1 0 2796 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1677677812
transform 1 0 2812 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_0
timestamp 1677677812
transform 1 0 2828 0 1 4625
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1677677812
transform 1 0 2820 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_80
timestamp 1677677812
transform 1 0 2820 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_28
timestamp 1677677812
transform 1 0 2852 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1677677812
transform 1 0 2876 0 1 4645
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1677677812
transform 1 0 2892 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_45
timestamp 1677677812
transform 1 0 2852 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1677677812
transform 1 0 2860 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_47
timestamp 1677677812
transform 1 0 2892 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_106
timestamp 1677677812
transform 1 0 2940 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_99
timestamp 1677677812
transform 1 0 2940 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_48
timestamp 1677677812
transform 1 0 3036 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1677677812
transform 1 0 2988 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_43
timestamp 1677677812
transform 1 0 3036 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1677677812
transform 1 0 2988 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_49
timestamp 1677677812
transform 1 0 3092 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1677677812
transform 1 0 3100 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1677677812
transform 1 0 3164 0 1 4675
box -3 -3 3 3
use M2_M1  M2_M1_50
timestamp 1677677812
transform 1 0 3172 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1677677812
transform 1 0 3140 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_82
timestamp 1677677812
transform 1 0 3140 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1677677812
transform 1 0 3132 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_51
timestamp 1677677812
transform 1 0 3244 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_45
timestamp 1677677812
transform 1 0 3268 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_52
timestamp 1677677812
transform 1 0 3308 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1677677812
transform 1 0 3364 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1677677812
transform 1 0 3372 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1677677812
transform 1 0 3284 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_46
timestamp 1677677812
transform 1 0 3308 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1677677812
transform 1 0 3284 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_55
timestamp 1677677812
transform 1 0 3436 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_47
timestamp 1677677812
transform 1 0 3436 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_110
timestamp 1677677812
transform 1 0 3460 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_84
timestamp 1677677812
transform 1 0 3460 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_10
timestamp 1677677812
transform 1 0 3484 0 1 4635
box -3 -3 3 3
use M2_M1  M2_M1_56
timestamp 1677677812
transform 1 0 3532 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_111
timestamp 1677677812
transform 1 0 3484 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1677677812
transform 1 0 3516 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1677677812
transform 1 0 3484 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1677677812
transform 1 0 3532 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1677677812
transform 1 0 3588 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_112
timestamp 1677677812
transform 1 0 3588 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_101
timestamp 1677677812
transform 1 0 3588 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1677677812
transform 1 0 3620 0 1 4625
box -3 -3 3 3
use M3_M2  M3_M2_31
timestamp 1677677812
transform 1 0 3644 0 1 4625
box -3 -3 3 3
use M2_M1  M2_M1_57
timestamp 1677677812
transform 1 0 3620 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_58
timestamp 1677677812
transform 1 0 3628 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_59
timestamp 1677677812
transform 1 0 3644 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1677677812
transform 1 0 3636 0 1 4605
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1677677812
transform 1 0 3652 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1677677812
transform 1 0 3636 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_102
timestamp 1677677812
transform 1 0 3628 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1677677812
transform 1 0 3684 0 1 4635
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1677677812
transform 1 0 3716 0 1 4635
box -3 -3 3 3
use M2_M1  M2_M1_60
timestamp 1677677812
transform 1 0 3732 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_115
timestamp 1677677812
transform 1 0 3684 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_49
timestamp 1677677812
transform 1 0 3732 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_50
timestamp 1677677812
transform 1 0 3756 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_103
timestamp 1677677812
transform 1 0 3724 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_61
timestamp 1677677812
transform 1 0 3780 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_104
timestamp 1677677812
transform 1 0 3788 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1677677812
transform 1 0 3820 0 1 4635
box -3 -3 3 3
use M2_M1  M2_M1_62
timestamp 1677677812
transform 1 0 3844 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1677677812
transform 1 0 3900 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1677677812
transform 1 0 3820 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1677677812
transform 1 0 3812 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_106
timestamp 1677677812
transform 1 0 3844 0 1 4585
box -3 -3 3 3
use M2_M1  M2_M1_64
timestamp 1677677812
transform 1 0 3932 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_51
timestamp 1677677812
transform 1 0 3940 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1677677812
transform 1 0 3956 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_65
timestamp 1677677812
transform 1 0 4004 0 1 4615
box -2 -2 2 2
use M3_M2  M3_M2_52
timestamp 1677677812
transform 1 0 4004 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_117
timestamp 1677677812
transform 1 0 4052 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_88
timestamp 1677677812
transform 1 0 4052 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_53
timestamp 1677677812
transform 1 0 4084 0 1 4605
box -3 -3 3 3
use M2_M1  M2_M1_66
timestamp 1677677812
transform 1 0 4124 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_67
timestamp 1677677812
transform 1 0 4180 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1677677812
transform 1 0 4100 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_54
timestamp 1677677812
transform 1 0 4124 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1677677812
transform 1 0 4100 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1677677812
transform 1 0 4116 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_68
timestamp 1677677812
transform 1 0 4244 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_69
timestamp 1677677812
transform 1 0 4300 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_119
timestamp 1677677812
transform 1 0 4220 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_91
timestamp 1677677812
transform 1 0 4220 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_70
timestamp 1677677812
transform 1 0 4364 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1677677812
transform 1 0 4420 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1677677812
transform 1 0 4340 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_92
timestamp 1677677812
transform 1 0 4340 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_107
timestamp 1677677812
transform 1 0 4332 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_108
timestamp 1677677812
transform 1 0 4364 0 1 4585
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1677677812
transform 1 0 4452 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_72
timestamp 1677677812
transform 1 0 4500 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1677677812
transform 1 0 4548 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1677677812
transform 1 0 4452 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_55
timestamp 1677677812
transform 1 0 4500 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1677677812
transform 1 0 4532 0 1 4605
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1677677812
transform 1 0 4452 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1677677812
transform 1 0 4660 0 1 4615
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1677677812
transform 1 0 4684 0 1 4615
box -3 -3 3 3
use M2_M1  M2_M1_74
timestamp 1677677812
transform 1 0 4708 0 1 4615
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1677677812
transform 1 0 4684 0 1 4605
box -2 -2 2 2
use M3_M2  M3_M2_94
timestamp 1677677812
transform 1 0 4684 0 1 4595
box -3 -3 3 3
use M3_M2  M3_M2_95
timestamp 1677677812
transform 1 0 4708 0 1 4595
box -3 -3 3 3
use M2_M1  M2_M1_75
timestamp 1677677812
transform 1 0 4780 0 1 4615
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_1
timestamp 1677677812
transform 1 0 4843 0 1 4670
box -10 -3 10 3
use top_level_VIA0  top_level_VIA0_2
timestamp 1677677812
transform 1 0 48 0 1 4570
box -10 -3 10 3
use FILL  FILL_0
timestamp 1677677812
transform 1 0 72 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1677677812
transform 1 0 80 0 1 4570
box -8 -3 104 105
use FILL  FILL_2
timestamp 1677677812
transform 1 0 176 0 1 4570
box -8 -3 16 105
use FILL  FILL_3
timestamp 1677677812
transform 1 0 184 0 1 4570
box -8 -3 16 105
use FILL  FILL_4
timestamp 1677677812
transform 1 0 192 0 1 4570
box -8 -3 16 105
use FILL  FILL_5
timestamp 1677677812
transform 1 0 200 0 1 4570
box -8 -3 16 105
use FILL  FILL_6
timestamp 1677677812
transform 1 0 208 0 1 4570
box -8 -3 16 105
use FILL  FILL_17
timestamp 1677677812
transform 1 0 216 0 1 4570
box -8 -3 16 105
use FILL  FILL_19
timestamp 1677677812
transform 1 0 224 0 1 4570
box -8 -3 16 105
use FILL  FILL_21
timestamp 1677677812
transform 1 0 232 0 1 4570
box -8 -3 16 105
use FILL  FILL_23
timestamp 1677677812
transform 1 0 240 0 1 4570
box -8 -3 16 105
use FILL  FILL_25
timestamp 1677677812
transform 1 0 248 0 1 4570
box -8 -3 16 105
use FILL  FILL_27
timestamp 1677677812
transform 1 0 256 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1677677812
transform -1 0 360 0 1 4570
box -8 -3 104 105
use FILL  FILL_28
timestamp 1677677812
transform 1 0 360 0 1 4570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1677677812
transform 1 0 368 0 1 4570
box -8 -3 16 105
use FILL  FILL_37
timestamp 1677677812
transform 1 0 376 0 1 4570
box -8 -3 16 105
use FILL  FILL_38
timestamp 1677677812
transform 1 0 384 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1677677812
transform 1 0 392 0 1 4570
box -8 -3 104 105
use FILL  FILL_39
timestamp 1677677812
transform 1 0 488 0 1 4570
box -8 -3 16 105
use FILL  FILL_40
timestamp 1677677812
transform 1 0 496 0 1 4570
box -8 -3 16 105
use FILL  FILL_46
timestamp 1677677812
transform 1 0 504 0 1 4570
box -8 -3 16 105
use FILL  FILL_48
timestamp 1677677812
transform 1 0 512 0 1 4570
box -8 -3 16 105
use FILL  FILL_50
timestamp 1677677812
transform 1 0 520 0 1 4570
box -8 -3 16 105
use FILL  FILL_51
timestamp 1677677812
transform 1 0 528 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1677677812
transform 1 0 536 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1677677812
transform -1 0 648 0 1 4570
box -8 -3 104 105
use FILL  FILL_52
timestamp 1677677812
transform 1 0 648 0 1 4570
box -8 -3 16 105
use FILL  FILL_53
timestamp 1677677812
transform 1 0 656 0 1 4570
box -8 -3 16 105
use FILL  FILL_62
timestamp 1677677812
transform 1 0 664 0 1 4570
box -8 -3 16 105
use FILL  FILL_64
timestamp 1677677812
transform 1 0 672 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_4
timestamp 1677677812
transform 1 0 680 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1677677812
transform 1 0 696 0 1 4570
box -8 -3 104 105
use FILL  FILL_66
timestamp 1677677812
transform 1 0 792 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1677677812
transform 1 0 800 0 1 4570
box -8 -3 104 105
use FILL  FILL_67
timestamp 1677677812
transform 1 0 896 0 1 4570
box -8 -3 16 105
use FILL  FILL_75
timestamp 1677677812
transform 1 0 904 0 1 4570
box -8 -3 16 105
use FILL  FILL_76
timestamp 1677677812
transform 1 0 912 0 1 4570
box -8 -3 16 105
use FILL  FILL_77
timestamp 1677677812
transform 1 0 920 0 1 4570
box -8 -3 16 105
use FILL  FILL_78
timestamp 1677677812
transform 1 0 928 0 1 4570
box -8 -3 16 105
use FILL  FILL_79
timestamp 1677677812
transform 1 0 936 0 1 4570
box -8 -3 16 105
use FILL  FILL_80
timestamp 1677677812
transform 1 0 944 0 1 4570
box -8 -3 16 105
use FILL  FILL_82
timestamp 1677677812
transform 1 0 952 0 1 4570
box -8 -3 16 105
use FILL  FILL_84
timestamp 1677677812
transform 1 0 960 0 1 4570
box -8 -3 16 105
use FILL  FILL_86
timestamp 1677677812
transform 1 0 968 0 1 4570
box -8 -3 16 105
use FILL  FILL_87
timestamp 1677677812
transform 1 0 976 0 1 4570
box -8 -3 16 105
use FILL  FILL_88
timestamp 1677677812
transform 1 0 984 0 1 4570
box -8 -3 16 105
use FILL  FILL_89
timestamp 1677677812
transform 1 0 992 0 1 4570
box -8 -3 16 105
use FILL  FILL_91
timestamp 1677677812
transform 1 0 1000 0 1 4570
box -8 -3 16 105
use FILL  FILL_93
timestamp 1677677812
transform 1 0 1008 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_7
timestamp 1677677812
transform 1 0 1016 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1677677812
transform -1 0 1128 0 1 4570
box -8 -3 104 105
use FILL  FILL_94
timestamp 1677677812
transform 1 0 1128 0 1 4570
box -8 -3 16 105
use FILL  FILL_95
timestamp 1677677812
transform 1 0 1136 0 1 4570
box -8 -3 16 105
use FILL  FILL_96
timestamp 1677677812
transform 1 0 1144 0 1 4570
box -8 -3 16 105
use FILL  FILL_97
timestamp 1677677812
transform 1 0 1152 0 1 4570
box -8 -3 16 105
use FILL  FILL_98
timestamp 1677677812
transform 1 0 1160 0 1 4570
box -8 -3 16 105
use FILL  FILL_99
timestamp 1677677812
transform 1 0 1168 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_8
timestamp 1677677812
transform -1 0 1272 0 1 4570
box -8 -3 104 105
use FILL  FILL_100
timestamp 1677677812
transform 1 0 1272 0 1 4570
box -8 -3 16 105
use FILL  FILL_101
timestamp 1677677812
transform 1 0 1280 0 1 4570
box -8 -3 16 105
use FILL  FILL_102
timestamp 1677677812
transform 1 0 1288 0 1 4570
box -8 -3 16 105
use FILL  FILL_103
timestamp 1677677812
transform 1 0 1296 0 1 4570
box -8 -3 16 105
use FILL  FILL_104
timestamp 1677677812
transform 1 0 1304 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1677677812
transform -1 0 1408 0 1 4570
box -8 -3 104 105
use FILL  FILL_105
timestamp 1677677812
transform 1 0 1408 0 1 4570
box -8 -3 16 105
use FILL  FILL_125
timestamp 1677677812
transform 1 0 1416 0 1 4570
box -8 -3 16 105
use FILL  FILL_126
timestamp 1677677812
transform 1 0 1424 0 1 4570
box -8 -3 16 105
use FILL  FILL_127
timestamp 1677677812
transform 1 0 1432 0 1 4570
box -8 -3 16 105
use FILL  FILL_128
timestamp 1677677812
transform 1 0 1440 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1677677812
transform -1 0 1544 0 1 4570
box -8 -3 104 105
use FILL  FILL_129
timestamp 1677677812
transform 1 0 1544 0 1 4570
box -8 -3 16 105
use FILL  FILL_137
timestamp 1677677812
transform 1 0 1552 0 1 4570
box -8 -3 16 105
use FILL  FILL_139
timestamp 1677677812
transform 1 0 1560 0 1 4570
box -8 -3 16 105
use FILL  FILL_141
timestamp 1677677812
transform 1 0 1568 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1677677812
transform 1 0 1576 0 1 4570
box -8 -3 104 105
use FILL  FILL_143
timestamp 1677677812
transform 1 0 1672 0 1 4570
box -8 -3 16 105
use FILL  FILL_144
timestamp 1677677812
transform 1 0 1680 0 1 4570
box -8 -3 16 105
use FILL  FILL_145
timestamp 1677677812
transform 1 0 1688 0 1 4570
box -8 -3 16 105
use FILL  FILL_146
timestamp 1677677812
transform 1 0 1696 0 1 4570
box -8 -3 16 105
use FILL  FILL_147
timestamp 1677677812
transform 1 0 1704 0 1 4570
box -8 -3 16 105
use FILL  FILL_148
timestamp 1677677812
transform 1 0 1712 0 1 4570
box -8 -3 16 105
use FILL  FILL_149
timestamp 1677677812
transform 1 0 1720 0 1 4570
box -8 -3 16 105
use FILL  FILL_150
timestamp 1677677812
transform 1 0 1728 0 1 4570
box -8 -3 16 105
use FILL  FILL_151
timestamp 1677677812
transform 1 0 1736 0 1 4570
box -8 -3 16 105
use FILL  FILL_152
timestamp 1677677812
transform 1 0 1744 0 1 4570
box -8 -3 16 105
use FILL  FILL_153
timestamp 1677677812
transform 1 0 1752 0 1 4570
box -8 -3 16 105
use FILL  FILL_154
timestamp 1677677812
transform 1 0 1760 0 1 4570
box -8 -3 16 105
use FILL  FILL_155
timestamp 1677677812
transform 1 0 1768 0 1 4570
box -8 -3 16 105
use FILL  FILL_156
timestamp 1677677812
transform 1 0 1776 0 1 4570
box -8 -3 16 105
use FILL  FILL_157
timestamp 1677677812
transform 1 0 1784 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_11
timestamp 1677677812
transform 1 0 1792 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1677677812
transform 1 0 1808 0 1 4570
box -8 -3 104 105
use FILL  FILL_158
timestamp 1677677812
transform 1 0 1904 0 1 4570
box -8 -3 16 105
use FILL  FILL_171
timestamp 1677677812
transform 1 0 1912 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1677677812
transform 1 0 1920 0 1 4570
box -8 -3 104 105
use FILL  FILL_173
timestamp 1677677812
transform 1 0 2016 0 1 4570
box -8 -3 16 105
use FILL  FILL_174
timestamp 1677677812
transform 1 0 2024 0 1 4570
box -8 -3 16 105
use FILL  FILL_175
timestamp 1677677812
transform 1 0 2032 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1677677812
transform 1 0 2040 0 1 4570
box -8 -3 104 105
use FILL  FILL_176
timestamp 1677677812
transform 1 0 2136 0 1 4570
box -8 -3 16 105
use FILL  FILL_177
timestamp 1677677812
transform 1 0 2144 0 1 4570
box -8 -3 16 105
use FILL  FILL_178
timestamp 1677677812
transform 1 0 2152 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_16
timestamp 1677677812
transform 1 0 2160 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1677677812
transform 1 0 2176 0 1 4570
box -8 -3 104 105
use FILL  FILL_179
timestamp 1677677812
transform 1 0 2272 0 1 4570
box -8 -3 16 105
use FILL  FILL_180
timestamp 1677677812
transform 1 0 2280 0 1 4570
box -8 -3 16 105
use FILL  FILL_181
timestamp 1677677812
transform 1 0 2288 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_17
timestamp 1677677812
transform -1 0 2392 0 1 4570
box -8 -3 104 105
use FILL  FILL_182
timestamp 1677677812
transform 1 0 2392 0 1 4570
box -8 -3 16 105
use FILL  FILL_183
timestamp 1677677812
transform 1 0 2400 0 1 4570
box -8 -3 16 105
use FILL  FILL_184
timestamp 1677677812
transform 1 0 2408 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1677677812
transform -1 0 2512 0 1 4570
box -8 -3 104 105
use FILL  FILL_185
timestamp 1677677812
transform 1 0 2512 0 1 4570
box -8 -3 16 105
use FILL  FILL_186
timestamp 1677677812
transform 1 0 2520 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_17
timestamp 1677677812
transform 1 0 2528 0 1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1677677812
transform 1 0 2544 0 1 4570
box -8 -3 104 105
use FILL  FILL_187
timestamp 1677677812
transform 1 0 2640 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_109
timestamp 1677677812
transform 1 0 2676 0 1 4575
box -3 -3 3 3
use INVX2  INVX2_18
timestamp 1677677812
transform 1 0 2648 0 1 4570
box -9 -3 26 105
use FILL  FILL_188
timestamp 1677677812
transform 1 0 2664 0 1 4570
box -8 -3 16 105
use FILL  FILL_189
timestamp 1677677812
transform 1 0 2672 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_110
timestamp 1677677812
transform 1 0 2780 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_20
timestamp 1677677812
transform 1 0 2680 0 1 4570
box -8 -3 104 105
use FILL  FILL_190
timestamp 1677677812
transform 1 0 2776 0 1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_4
timestamp 1677677812
transform 1 0 2784 0 1 4570
box -8 -3 34 105
use FILL  FILL_191
timestamp 1677677812
transform 1 0 2816 0 1 4570
box -8 -3 16 105
use FILL  FILL_192
timestamp 1677677812
transform 1 0 2824 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_111
timestamp 1677677812
transform 1 0 2844 0 1 4575
box -3 -3 3 3
use INVX2  INVX2_19
timestamp 1677677812
transform 1 0 2832 0 1 4570
box -9 -3 26 105
use FILL  FILL_193
timestamp 1677677812
transform 1 0 2848 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_112
timestamp 1677677812
transform 1 0 2876 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_21
timestamp 1677677812
transform -1 0 2952 0 1 4570
box -8 -3 104 105
use FILL  FILL_194
timestamp 1677677812
transform 1 0 2952 0 1 4570
box -8 -3 16 105
use FILL  FILL_195
timestamp 1677677812
transform 1 0 2960 0 1 4570
box -8 -3 16 105
use FILL  FILL_196
timestamp 1677677812
transform 1 0 2968 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1677677812
transform 1 0 2976 0 1 4570
box -8 -3 104 105
use FILL  FILL_197
timestamp 1677677812
transform 1 0 3072 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_20
timestamp 1677677812
transform 1 0 3080 0 1 4570
box -9 -3 26 105
use FILL  FILL_198
timestamp 1677677812
transform 1 0 3096 0 1 4570
box -8 -3 16 105
use FILL  FILL_199
timestamp 1677677812
transform 1 0 3104 0 1 4570
box -8 -3 16 105
use FILL  FILL_200
timestamp 1677677812
transform 1 0 3112 0 1 4570
box -8 -3 16 105
use FILL  FILL_201
timestamp 1677677812
transform 1 0 3120 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_23
timestamp 1677677812
transform 1 0 3128 0 1 4570
box -8 -3 104 105
use FILL  FILL_255
timestamp 1677677812
transform 1 0 3224 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_27
timestamp 1677677812
transform 1 0 3232 0 1 4570
box -9 -3 26 105
use FILL  FILL_264
timestamp 1677677812
transform 1 0 3248 0 1 4570
box -8 -3 16 105
use FILL  FILL_265
timestamp 1677677812
transform 1 0 3256 0 1 4570
box -8 -3 16 105
use FILL  FILL_266
timestamp 1677677812
transform 1 0 3264 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_113
timestamp 1677677812
transform 1 0 3284 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_24
timestamp 1677677812
transform 1 0 3272 0 1 4570
box -8 -3 104 105
use FILL  FILL_267
timestamp 1677677812
transform 1 0 3368 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_25
timestamp 1677677812
transform -1 0 3472 0 1 4570
box -8 -3 104 105
use M3_M2  M3_M2_114
timestamp 1677677812
transform 1 0 3508 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_26
timestamp 1677677812
transform 1 0 3472 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_28
timestamp 1677677812
transform 1 0 3568 0 1 4570
box -9 -3 26 105
use FILL  FILL_268
timestamp 1677677812
transform 1 0 3584 0 1 4570
box -8 -3 16 105
use FILL  FILL_269
timestamp 1677677812
transform 1 0 3592 0 1 4570
box -8 -3 16 105
use FILL  FILL_270
timestamp 1677677812
transform 1 0 3600 0 1 4570
box -8 -3 16 105
use FILL  FILL_271
timestamp 1677677812
transform 1 0 3608 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_115
timestamp 1677677812
transform 1 0 3628 0 1 4575
box -3 -3 3 3
use M3_M2  M3_M2_116
timestamp 1677677812
transform 1 0 3652 0 1 4575
box -3 -3 3 3
use OAI22X1  OAI22X1_11
timestamp 1677677812
transform 1 0 3616 0 1 4570
box -8 -3 46 105
use FILL  FILL_297
timestamp 1677677812
transform 1 0 3656 0 1 4570
box -8 -3 16 105
use FILL  FILL_298
timestamp 1677677812
transform 1 0 3664 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_117
timestamp 1677677812
transform 1 0 3772 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_27
timestamp 1677677812
transform 1 0 3672 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_31
timestamp 1677677812
transform 1 0 3768 0 1 4570
box -9 -3 26 105
use FILL  FILL_299
timestamp 1677677812
transform 1 0 3784 0 1 4570
box -8 -3 16 105
use FILL  FILL_312
timestamp 1677677812
transform 1 0 3792 0 1 4570
box -8 -3 16 105
use FILL  FILL_313
timestamp 1677677812
transform 1 0 3800 0 1 4570
box -8 -3 16 105
use M3_M2  M3_M2_118
timestamp 1677677812
transform 1 0 3828 0 1 4575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_28
timestamp 1677677812
transform 1 0 3808 0 1 4570
box -8 -3 104 105
use FILL  FILL_314
timestamp 1677677812
transform 1 0 3904 0 1 4570
box -8 -3 16 105
use FILL  FILL_323
timestamp 1677677812
transform 1 0 3912 0 1 4570
box -8 -3 16 105
use FILL  FILL_324
timestamp 1677677812
transform 1 0 3920 0 1 4570
box -8 -3 16 105
use FILL  FILL_325
timestamp 1677677812
transform 1 0 3928 0 1 4570
box -8 -3 16 105
use INVX2  INVX2_33
timestamp 1677677812
transform -1 0 3952 0 1 4570
box -9 -3 26 105
use FILL  FILL_326
timestamp 1677677812
transform 1 0 3952 0 1 4570
box -8 -3 16 105
use FILL  FILL_327
timestamp 1677677812
transform 1 0 3960 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1677677812
transform -1 0 4064 0 1 4570
box -8 -3 104 105
use FILL  FILL_328
timestamp 1677677812
transform 1 0 4064 0 1 4570
box -8 -3 16 105
use FILL  FILL_329
timestamp 1677677812
transform 1 0 4072 0 1 4570
box -8 -3 16 105
use FILL  FILL_330
timestamp 1677677812
transform 1 0 4080 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1677677812
transform 1 0 4088 0 1 4570
box -8 -3 104 105
use FILL  FILL_331
timestamp 1677677812
transform 1 0 4184 0 1 4570
box -8 -3 16 105
use FILL  FILL_350
timestamp 1677677812
transform 1 0 4192 0 1 4570
box -8 -3 16 105
use FILL  FILL_352
timestamp 1677677812
transform 1 0 4200 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_31
timestamp 1677677812
transform 1 0 4208 0 1 4570
box -8 -3 104 105
use FILL  FILL_354
timestamp 1677677812
transform 1 0 4304 0 1 4570
box -8 -3 16 105
use FILL  FILL_361
timestamp 1677677812
transform 1 0 4312 0 1 4570
box -8 -3 16 105
use FILL  FILL_362
timestamp 1677677812
transform 1 0 4320 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_32
timestamp 1677677812
transform 1 0 4328 0 1 4570
box -8 -3 104 105
use FILL  FILL_363
timestamp 1677677812
transform 1 0 4424 0 1 4570
box -8 -3 16 105
use FILL  FILL_364
timestamp 1677677812
transform 1 0 4432 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1677677812
transform 1 0 4440 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_36
timestamp 1677677812
transform 1 0 4536 0 1 4570
box -9 -3 26 105
use FILL  FILL_365
timestamp 1677677812
transform 1 0 4552 0 1 4570
box -8 -3 16 105
use FILL  FILL_366
timestamp 1677677812
transform 1 0 4560 0 1 4570
box -8 -3 16 105
use FILL  FILL_367
timestamp 1677677812
transform 1 0 4568 0 1 4570
box -8 -3 16 105
use FILL  FILL_368
timestamp 1677677812
transform 1 0 4576 0 1 4570
box -8 -3 16 105
use FILL  FILL_369
timestamp 1677677812
transform 1 0 4584 0 1 4570
box -8 -3 16 105
use FILL  FILL_370
timestamp 1677677812
transform 1 0 4592 0 1 4570
box -8 -3 16 105
use FILL  FILL_385
timestamp 1677677812
transform 1 0 4600 0 1 4570
box -8 -3 16 105
use FILL  FILL_387
timestamp 1677677812
transform 1 0 4608 0 1 4570
box -8 -3 16 105
use FILL  FILL_389
timestamp 1677677812
transform 1 0 4616 0 1 4570
box -8 -3 16 105
use FILL  FILL_391
timestamp 1677677812
transform 1 0 4624 0 1 4570
box -8 -3 16 105
use FILL  FILL_393
timestamp 1677677812
transform 1 0 4632 0 1 4570
box -8 -3 16 105
use FILL  FILL_395
timestamp 1677677812
transform 1 0 4640 0 1 4570
box -8 -3 16 105
use FILL  FILL_397
timestamp 1677677812
transform 1 0 4648 0 1 4570
box -8 -3 16 105
use FILL  FILL_399
timestamp 1677677812
transform 1 0 4656 0 1 4570
box -8 -3 16 105
use FILL  FILL_401
timestamp 1677677812
transform 1 0 4664 0 1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1677677812
transform 1 0 4672 0 1 4570
box -8 -3 104 105
use INVX2  INVX2_38
timestamp 1677677812
transform 1 0 4768 0 1 4570
box -9 -3 26 105
use FILL  FILL_402
timestamp 1677677812
transform 1 0 4784 0 1 4570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_3
timestamp 1677677812
transform 1 0 4819 0 1 4570
box -10 -3 10 3
use M2_M1  M2_M1_276
timestamp 1677677812
transform 1 0 124 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_153
timestamp 1677677812
transform 1 0 172 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_154
timestamp 1677677812
transform 1 0 188 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_127
timestamp 1677677812
transform 1 0 172 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1677677812
transform 1 0 180 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1677677812
transform 1 0 172 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_227
timestamp 1677677812
transform 1 0 180 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_278
timestamp 1677677812
transform 1 0 188 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_269
timestamp 1677677812
transform 1 0 172 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_279
timestamp 1677677812
transform 1 0 220 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1677677812
transform 1 0 228 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_280
timestamp 1677677812
transform 1 0 236 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_130
timestamp 1677677812
transform 1 0 276 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_129
timestamp 1677677812
transform 1 0 276 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1677677812
transform 1 0 292 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1677677812
transform 1 0 300 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_229
timestamp 1677677812
transform 1 0 268 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_281
timestamp 1677677812
transform 1 0 284 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_230
timestamp 1677677812
transform 1 0 292 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_282
timestamp 1677677812
transform 1 0 300 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_231
timestamp 1677677812
transform 1 0 308 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_283
timestamp 1677677812
transform 1 0 316 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_270
timestamp 1677677812
transform 1 0 300 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_132
timestamp 1677677812
transform 1 0 372 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_271
timestamp 1677677812
transform 1 0 372 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_131
timestamp 1677677812
transform 1 0 412 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1677677812
transform 1 0 396 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_133
timestamp 1677677812
transform 1 0 396 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1677677812
transform 1 0 412 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1677677812
transform 1 0 380 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1677677812
transform 1 0 388 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1677677812
transform 1 0 404 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_272
timestamp 1677677812
transform 1 0 404 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_319
timestamp 1677677812
transform 1 0 388 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_132
timestamp 1677677812
transform 1 0 428 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_320
timestamp 1677677812
transform 1 0 444 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_156
timestamp 1677677812
transform 1 0 492 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_135
timestamp 1677677812
transform 1 0 460 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1677677812
transform 1 0 476 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_137
timestamp 1677677812
transform 1 0 492 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1677677812
transform 1 0 452 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1677677812
transform 1 0 468 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1677677812
transform 1 0 492 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_273
timestamp 1677677812
transform 1 0 492 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_335
timestamp 1677677812
transform 1 0 476 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1677677812
transform 1 0 468 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_290
timestamp 1677677812
transform 1 0 508 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_321
timestamp 1677677812
transform 1 0 508 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_119
timestamp 1677677812
transform 1 0 540 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_120
timestamp 1677677812
transform 1 0 556 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_133
timestamp 1677677812
transform 1 0 556 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1677677812
transform 1 0 532 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_138
timestamp 1677677812
transform 1 0 540 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1677677812
transform 1 0 556 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1677677812
transform 1 0 532 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_292
timestamp 1677677812
transform 1 0 548 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_349
timestamp 1677677812
transform 1 0 556 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_293
timestamp 1677677812
transform 1 0 588 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1677677812
transform 1 0 612 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_196
timestamp 1677677812
transform 1 0 652 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_295
timestamp 1677677812
transform 1 0 636 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1677677812
transform 1 0 652 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_350
timestamp 1677677812
transform 1 0 652 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1677677812
transform 1 0 684 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1677677812
transform 1 0 724 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_140
timestamp 1677677812
transform 1 0 684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1677677812
transform 1 0 692 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1677677812
transform 1 0 708 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_197
timestamp 1677677812
transform 1 0 716 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_143
timestamp 1677677812
transform 1 0 724 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1677677812
transform 1 0 700 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1677677812
transform 1 0 716 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_274
timestamp 1677677812
transform 1 0 716 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1677677812
transform 1 0 700 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_144
timestamp 1677677812
transform 1 0 756 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_159
timestamp 1677677812
transform 1 0 780 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_299
timestamp 1677677812
transform 1 0 780 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_275
timestamp 1677677812
transform 1 0 780 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_145
timestamp 1677677812
transform 1 0 796 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_232
timestamp 1677677812
transform 1 0 796 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_300
timestamp 1677677812
transform 1 0 820 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_233
timestamp 1677677812
transform 1 0 836 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_301
timestamp 1677677812
transform 1 0 876 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_302
timestamp 1677677812
transform 1 0 884 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1677677812
transform 1 0 892 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_276
timestamp 1677677812
transform 1 0 820 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_134
timestamp 1677677812
transform 1 0 940 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_123
timestamp 1677677812
transform 1 0 948 0 1 4545
box -2 -2 2 2
use M2_M1  M2_M1_146
timestamp 1677677812
transform 1 0 908 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1677677812
transform 1 0 916 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_148
timestamp 1677677812
transform 1 0 940 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_234
timestamp 1677677812
transform 1 0 916 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_198
timestamp 1677677812
transform 1 0 948 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_304
timestamp 1677677812
transform 1 0 924 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1677677812
transform 1 0 940 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_277
timestamp 1677677812
transform 1 0 940 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_149
timestamp 1677677812
transform 1 0 964 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1677677812
transform 1 0 988 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_235
timestamp 1677677812
transform 1 0 988 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_160
timestamp 1677677812
transform 1 0 1004 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_199
timestamp 1677677812
transform 1 0 1012 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_151
timestamp 1677677812
transform 1 0 1036 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1677677812
transform 1 0 1004 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_307
timestamp 1677677812
transform 1 0 1012 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1677677812
transform 1 0 1028 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1677677812
transform 1 0 1044 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_278
timestamp 1677677812
transform 1 0 996 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1677677812
transform 1 0 1044 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_336
timestamp 1677677812
transform 1 0 1028 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_135
timestamp 1677677812
transform 1 0 1060 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_152
timestamp 1677677812
transform 1 0 1060 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_161
timestamp 1677677812
transform 1 0 1084 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_153
timestamp 1677677812
transform 1 0 1084 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1677677812
transform 1 0 1092 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_310
timestamp 1677677812
transform 1 0 1060 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1677677812
transform 1 0 1068 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1677677812
transform 1 0 1084 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_337
timestamp 1677677812
transform 1 0 1068 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1677677812
transform 1 0 1092 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1677677812
transform 1 0 1116 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_434
timestamp 1677677812
transform 1 0 1116 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1677677812
transform 1 0 1164 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_156
timestamp 1677677812
transform 1 0 1188 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_157
timestamp 1677677812
transform 1 0 1196 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1677677812
transform 1 0 1140 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1677677812
transform 1 0 1156 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1677677812
transform 1 0 1164 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1677677812
transform 1 0 1172 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_280
timestamp 1677677812
transform 1 0 1140 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_322
timestamp 1677677812
transform 1 0 1156 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_435
timestamp 1677677812
transform 1 0 1188 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1677677812
transform 1 0 1196 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1677677812
transform 1 0 1164 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_158
timestamp 1677677812
transform 1 0 1212 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_238
timestamp 1677677812
transform 1 0 1212 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_317
timestamp 1677677812
transform 1 0 1228 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1677677812
transform 1 0 1236 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1677677812
transform 1 0 1236 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_136
timestamp 1677677812
transform 1 0 1268 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_159
timestamp 1677677812
transform 1 0 1268 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_160
timestamp 1677677812
transform 1 0 1276 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_282
timestamp 1677677812
transform 1 0 1260 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_162
timestamp 1677677812
transform 1 0 1308 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_161
timestamp 1677677812
transform 1 0 1308 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1677677812
transform 1 0 1316 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_318
timestamp 1677677812
transform 1 0 1284 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_319
timestamp 1677677812
transform 1 0 1300 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_320
timestamp 1677677812
transform 1 0 1308 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_437
timestamp 1677677812
transform 1 0 1284 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_324
timestamp 1677677812
transform 1 0 1284 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_283
timestamp 1677677812
transform 1 0 1308 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_163
timestamp 1677677812
transform 1 0 1364 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_321
timestamp 1677677812
transform 1 0 1364 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_163
timestamp 1677677812
transform 1 0 1420 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1677677812
transform 1 0 1428 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_165
timestamp 1677677812
transform 1 0 1444 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_239
timestamp 1677677812
transform 1 0 1428 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_322
timestamp 1677677812
transform 1 0 1436 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_284
timestamp 1677677812
transform 1 0 1436 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_240
timestamp 1677677812
transform 1 0 1468 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_121
timestamp 1677677812
transform 1 0 1492 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_323
timestamp 1677677812
transform 1 0 1484 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_285
timestamp 1677677812
transform 1 0 1484 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_164
timestamp 1677677812
transform 1 0 1508 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_166
timestamp 1677677812
transform 1 0 1492 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1677677812
transform 1 0 1500 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_168
timestamp 1677677812
transform 1 0 1516 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_241
timestamp 1677677812
transform 1 0 1500 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_200
timestamp 1677677812
transform 1 0 1532 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1677677812
transform 1 0 1540 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_324
timestamp 1677677812
transform 1 0 1508 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_325
timestamp 1677677812
transform 1 0 1524 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_286
timestamp 1677677812
transform 1 0 1524 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_326
timestamp 1677677812
transform 1 0 1572 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_137
timestamp 1677677812
transform 1 0 1612 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_170
timestamp 1677677812
transform 1 0 1588 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_201
timestamp 1677677812
transform 1 0 1596 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_171
timestamp 1677677812
transform 1 0 1604 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_172
timestamp 1677677812
transform 1 0 1620 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1677677812
transform 1 0 1636 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_242
timestamp 1677677812
transform 1 0 1604 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_327
timestamp 1677677812
transform 1 0 1612 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_328
timestamp 1677677812
transform 1 0 1628 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_287
timestamp 1677677812
transform 1 0 1628 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_174
timestamp 1677677812
transform 1 0 1652 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_138
timestamp 1677677812
transform 1 0 1660 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_243
timestamp 1677677812
transform 1 0 1652 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_329
timestamp 1677677812
transform 1 0 1660 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_352
timestamp 1677677812
transform 1 0 1660 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1677677812
transform 1 0 1692 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1677677812
transform 1 0 1676 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_176
timestamp 1677677812
transform 1 0 1692 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1677677812
transform 1 0 1740 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1677677812
transform 1 0 1772 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1677677812
transform 1 0 1780 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_288
timestamp 1677677812
transform 1 0 1740 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_289
timestamp 1677677812
transform 1 0 1780 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_333
timestamp 1677677812
transform 1 0 1796 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_353
timestamp 1677677812
transform 1 0 1796 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1677677812
transform 1 0 1820 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1677677812
transform 1 0 1820 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_167
timestamp 1677677812
transform 1 0 1836 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1677677812
transform 1 0 1836 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_122
timestamp 1677677812
transform 1 0 1868 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_334
timestamp 1677677812
transform 1 0 1844 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_335
timestamp 1677677812
transform 1 0 1860 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1677677812
transform 1 0 1868 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1677677812
transform 1 0 1860 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_123
timestamp 1677677812
transform 1 0 1900 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_179
timestamp 1677677812
transform 1 0 1884 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_180
timestamp 1677677812
transform 1 0 1892 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_339
timestamp 1677677812
transform 1 0 1892 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1677677812
transform 1 0 1908 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_181
timestamp 1677677812
transform 1 0 1908 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1677677812
transform 1 0 1908 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_291
timestamp 1677677812
transform 1 0 1908 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_182
timestamp 1677677812
transform 1 0 1924 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_244
timestamp 1677677812
transform 1 0 1924 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1677677812
transform 1 0 1940 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_183
timestamp 1677677812
transform 1 0 1940 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1677677812
transform 1 0 1964 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_202
timestamp 1677677812
transform 1 0 1972 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_338
timestamp 1677677812
transform 1 0 1956 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1677677812
transform 1 0 1964 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_339
timestamp 1677677812
transform 1 0 1972 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_170
timestamp 1677677812
transform 1 0 2028 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_185
timestamp 1677677812
transform 1 0 2036 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1677677812
transform 1 0 2052 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_340
timestamp 1677677812
transform 1 0 2012 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_341
timestamp 1677677812
transform 1 0 2028 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_342
timestamp 1677677812
transform 1 0 2044 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_325
timestamp 1677677812
transform 1 0 2012 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1677677812
transform 1 0 2044 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_203
timestamp 1677677812
transform 1 0 2060 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_187
timestamp 1677677812
transform 1 0 2068 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1677677812
transform 1 0 2068 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_343
timestamp 1677677812
transform 1 0 2076 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_344
timestamp 1677677812
transform 1 0 2084 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_340
timestamp 1677677812
transform 1 0 2084 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1677677812
transform 1 0 2140 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_204
timestamp 1677677812
transform 1 0 2132 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_188
timestamp 1677677812
transform 1 0 2140 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1677677812
transform 1 0 2164 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_189
timestamp 1677677812
transform 1 0 2164 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1677677812
transform 1 0 2132 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_346
timestamp 1677677812
transform 1 0 2148 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_347
timestamp 1677677812
transform 1 0 2156 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_247
timestamp 1677677812
transform 1 0 2164 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_348
timestamp 1677677812
transform 1 0 2172 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_293
timestamp 1677677812
transform 1 0 2148 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1677677812
transform 1 0 2156 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_327
timestamp 1677677812
transform 1 0 2180 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_354
timestamp 1677677812
transform 1 0 2156 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_355
timestamp 1677677812
transform 1 0 2172 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1677677812
transform 1 0 2196 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_349
timestamp 1677677812
transform 1 0 2196 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_350
timestamp 1677677812
transform 1 0 2212 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_124
timestamp 1677677812
transform 1 0 2236 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_172
timestamp 1677677812
transform 1 0 2228 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1677677812
transform 1 0 2228 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1677677812
transform 1 0 2236 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_125
timestamp 1677677812
transform 1 0 2252 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_173
timestamp 1677677812
transform 1 0 2268 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_192
timestamp 1677677812
transform 1 0 2260 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_206
timestamp 1677677812
transform 1 0 2284 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_193
timestamp 1677677812
transform 1 0 2300 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_194
timestamp 1677677812
transform 1 0 2316 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1677677812
transform 1 0 2324 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1677677812
transform 1 0 2244 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1677677812
transform 1 0 2268 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_294
timestamp 1677677812
transform 1 0 2244 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_341
timestamp 1677677812
transform 1 0 2268 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_353
timestamp 1677677812
transform 1 0 2284 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_140
timestamp 1677677812
transform 1 0 2356 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_354
timestamp 1677677812
transform 1 0 2308 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_355
timestamp 1677677812
transform 1 0 2324 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1677677812
transform 1 0 2340 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1677677812
transform 1 0 2348 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1677677812
transform 1 0 2316 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1677677812
transform 1 0 2348 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_196
timestamp 1677677812
transform 1 0 2356 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_141
timestamp 1677677812
transform 1 0 2380 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_197
timestamp 1677677812
transform 1 0 2380 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_207
timestamp 1677677812
transform 1 0 2404 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_198
timestamp 1677677812
transform 1 0 2412 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1677677812
transform 1 0 2428 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1677677812
transform 1 0 2436 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1677677812
transform 1 0 2388 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1677677812
transform 1 0 2404 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1677677812
transform 1 0 2420 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1677677812
transform 1 0 2436 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_342
timestamp 1677677812
transform 1 0 2388 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1677677812
transform 1 0 2436 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_362
timestamp 1677677812
transform 1 0 2468 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1677677812
transform 1 0 2476 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_201
timestamp 1677677812
transform 1 0 2524 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_248
timestamp 1677677812
transform 1 0 2524 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_364
timestamp 1677677812
transform 1 0 2532 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_174
timestamp 1677677812
transform 1 0 2572 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_202
timestamp 1677677812
transform 1 0 2572 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1677677812
transform 1 0 2580 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_208
timestamp 1677677812
transform 1 0 2588 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_249
timestamp 1677677812
transform 1 0 2580 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_204
timestamp 1677677812
transform 1 0 2604 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1677677812
transform 1 0 2588 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1677677812
transform 1 0 2596 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_250
timestamp 1677677812
transform 1 0 2604 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_297
timestamp 1677677812
transform 1 0 2596 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1677677812
transform 1 0 2636 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1677677812
transform 1 0 2684 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1677677812
transform 1 0 2716 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_205
timestamp 1677677812
transform 1 0 2644 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_209
timestamp 1677677812
transform 1 0 2668 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_206
timestamp 1677677812
transform 1 0 2676 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1677677812
transform 1 0 2684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1677677812
transform 1 0 2700 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1677677812
transform 1 0 2644 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_210
timestamp 1677677812
transform 1 0 2708 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_209
timestamp 1677677812
transform 1 0 2716 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1677677812
transform 1 0 2652 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_368
timestamp 1677677812
transform 1 0 2668 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_369
timestamp 1677677812
transform 1 0 2676 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_252
timestamp 1677677812
transform 1 0 2684 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_370
timestamp 1677677812
transform 1 0 2692 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1677677812
transform 1 0 2700 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_142
timestamp 1677677812
transform 1 0 2756 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_124
timestamp 1677677812
transform 1 0 2756 0 1 4545
box -2 -2 2 2
use M3_M2  M3_M2_211
timestamp 1677677812
transform 1 0 2748 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_371
timestamp 1677677812
transform 1 0 2708 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1677677812
transform 1 0 2716 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1677677812
transform 1 0 2732 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_374
timestamp 1677677812
transform 1 0 2748 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_356
timestamp 1677677812
transform 1 0 2676 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_178
timestamp 1677677812
transform 1 0 2764 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_210
timestamp 1677677812
transform 1 0 2764 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_211
timestamp 1677677812
transform 1 0 2780 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_212
timestamp 1677677812
transform 1 0 2788 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_212
timestamp 1677677812
transform 1 0 2796 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_254
timestamp 1677677812
transform 1 0 2788 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1677677812
transform 1 0 2780 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1677677812
transform 1 0 2828 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1677677812
transform 1 0 2812 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1677677812
transform 1 0 2828 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_375
timestamp 1677677812
transform 1 0 2804 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1677677812
transform 1 0 2812 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_143
timestamp 1677677812
transform 1 0 2852 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_125
timestamp 1677677812
transform 1 0 2844 0 1 4545
box -2 -2 2 2
use M3_M2  M3_M2_179
timestamp 1677677812
transform 1 0 2860 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_213
timestamp 1677677812
transform 1 0 2844 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_214
timestamp 1677677812
transform 1 0 2852 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1677677812
transform 1 0 2860 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_215
timestamp 1677677812
transform 1 0 2868 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_377
timestamp 1677677812
transform 1 0 2860 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1677677812
transform 1 0 2868 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1677677812
transform 1 0 2836 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_298
timestamp 1677677812
transform 1 0 2844 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_216
timestamp 1677677812
transform 1 0 2916 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_299
timestamp 1677677812
transform 1 0 2932 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_439
timestamp 1677677812
transform 1 0 2940 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_329
timestamp 1677677812
transform 1 0 2940 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_217
timestamp 1677677812
transform 1 0 2972 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_127
timestamp 1677677812
transform 1 0 2980 0 1 4565
box -3 -3 3 3
use M2_M1  M2_M1_218
timestamp 1677677812
transform 1 0 2980 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_180
timestamp 1677677812
transform 1 0 3004 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_219
timestamp 1677677812
transform 1 0 3004 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1677677812
transform 1 0 3012 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_379
timestamp 1677677812
transform 1 0 2980 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_380
timestamp 1677677812
transform 1 0 2996 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_300
timestamp 1677677812
transform 1 0 2972 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_440
timestamp 1677677812
transform 1 0 2980 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_330
timestamp 1677677812
transform 1 0 2980 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_441
timestamp 1677677812
transform 1 0 3020 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_331
timestamp 1677677812
transform 1 0 3020 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_381
timestamp 1677677812
transform 1 0 3044 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1677677812
transform 1 0 3060 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_221
timestamp 1677677812
transform 1 0 3076 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_222
timestamp 1677677812
transform 1 0 3084 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1677677812
transform 1 0 3100 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1677677812
transform 1 0 3092 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_255
timestamp 1677677812
transform 1 0 3100 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_384
timestamp 1677677812
transform 1 0 3108 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_301
timestamp 1677677812
transform 1 0 3092 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_224
timestamp 1677677812
transform 1 0 3132 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_181
timestamp 1677677812
transform 1 0 3180 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_225
timestamp 1677677812
transform 1 0 3156 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_216
timestamp 1677677812
transform 1 0 3164 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_226
timestamp 1677677812
transform 1 0 3172 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_227
timestamp 1677677812
transform 1 0 3188 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1677677812
transform 1 0 3164 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_386
timestamp 1677677812
transform 1 0 3180 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_302
timestamp 1677677812
transform 1 0 3156 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_256
timestamp 1677677812
transform 1 0 3188 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1677677812
transform 1 0 3212 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_182
timestamp 1677677812
transform 1 0 3244 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_228
timestamp 1677677812
transform 1 0 3252 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_229
timestamp 1677677812
transform 1 0 3268 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_218
timestamp 1677677812
transform 1 0 3276 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_230
timestamp 1677677812
transform 1 0 3284 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_219
timestamp 1677677812
transform 1 0 3292 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_387
timestamp 1677677812
transform 1 0 3260 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1677677812
transform 1 0 3276 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_389
timestamp 1677677812
transform 1 0 3284 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_303
timestamp 1677677812
transform 1 0 3260 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_304
timestamp 1677677812
transform 1 0 3284 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1677677812
transform 1 0 3356 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_126
timestamp 1677677812
transform 1 0 3364 0 1 4545
box -2 -2 2 2
use M2_M1  M2_M1_231
timestamp 1677677812
transform 1 0 3372 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1677677812
transform 1 0 3388 0 1 4515
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1677677812
transform 1 0 3404 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_305
timestamp 1677677812
transform 1 0 3404 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1677677812
transform 1 0 3428 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1677677812
transform 1 0 3436 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_232
timestamp 1677677812
transform 1 0 3444 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1677677812
transform 1 0 3428 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_444
timestamp 1677677812
transform 1 0 3420 0 1 4505
box -2 -2 2 2
use M3_M2  M3_M2_344
timestamp 1677677812
transform 1 0 3420 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1677677812
transform 1 0 3436 0 1 4485
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1677677812
transform 1 0 3484 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_443
timestamp 1677677812
transform 1 0 3492 0 1 4515
box -2 -2 2 2
use M3_M2  M3_M2_183
timestamp 1677677812
transform 1 0 3532 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_233
timestamp 1677677812
transform 1 0 3516 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_234
timestamp 1677677812
transform 1 0 3532 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1677677812
transform 1 0 3540 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1677677812
transform 1 0 3508 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1677677812
transform 1 0 3524 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_306
timestamp 1677677812
transform 1 0 3524 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_307
timestamp 1677677812
transform 1 0 3540 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1677677812
transform 1 0 3556 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_145
timestamp 1677677812
transform 1 0 3604 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_236
timestamp 1677677812
transform 1 0 3604 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_394
timestamp 1677677812
transform 1 0 3572 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1677677812
transform 1 0 3588 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_332
timestamp 1677677812
transform 1 0 3572 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_184
timestamp 1677677812
transform 1 0 3652 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_237
timestamp 1677677812
transform 1 0 3644 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_396
timestamp 1677677812
transform 1 0 3644 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1677677812
transform 1 0 3652 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_398
timestamp 1677677812
transform 1 0 3668 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1677677812
transform 1 0 3684 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_308
timestamp 1677677812
transform 1 0 3644 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_333
timestamp 1677677812
transform 1 0 3652 0 1 4505
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1677677812
transform 1 0 3684 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1677677812
transform 1 0 3732 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_238
timestamp 1677677812
transform 1 0 3732 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1677677812
transform 1 0 3740 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_240
timestamp 1677677812
transform 1 0 3756 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1677677812
transform 1 0 3772 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_400
timestamp 1677677812
transform 1 0 3724 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_258
timestamp 1677677812
transform 1 0 3740 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_401
timestamp 1677677812
transform 1 0 3764 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_334
timestamp 1677677812
transform 1 0 3756 0 1 4505
box -3 -3 3 3
use M2_M1  M2_M1_242
timestamp 1677677812
transform 1 0 3796 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1677677812
transform 1 0 3812 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1677677812
transform 1 0 3828 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_402
timestamp 1677677812
transform 1 0 3788 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_403
timestamp 1677677812
transform 1 0 3820 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_404
timestamp 1677677812
transform 1 0 3836 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_245
timestamp 1677677812
transform 1 0 3852 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_405
timestamp 1677677812
transform 1 0 3860 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1677677812
transform 1 0 3900 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_186
timestamp 1677677812
transform 1 0 3932 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_187
timestamp 1677677812
transform 1 0 3956 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_247
timestamp 1677677812
transform 1 0 3924 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_248
timestamp 1677677812
transform 1 0 3940 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_249
timestamp 1677677812
transform 1 0 3956 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1677677812
transform 1 0 3964 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_259
timestamp 1677677812
transform 1 0 3924 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_406
timestamp 1677677812
transform 1 0 3932 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_310
timestamp 1677677812
transform 1 0 3964 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_345
timestamp 1677677812
transform 1 0 3964 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1677677812
transform 1 0 3988 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_251
timestamp 1677677812
transform 1 0 4020 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_252
timestamp 1677677812
transform 1 0 4036 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1677677812
transform 1 0 4004 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_408
timestamp 1677677812
transform 1 0 4028 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_311
timestamp 1677677812
transform 1 0 4004 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_261
timestamp 1677677812
transform 1 0 4036 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_146
timestamp 1677677812
transform 1 0 4076 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1677677812
transform 1 0 4084 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_222
timestamp 1677677812
transform 1 0 4092 0 1 4535
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1677677812
transform 1 0 4108 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_254
timestamp 1677677812
transform 1 0 4100 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1677677812
transform 1 0 4076 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1677677812
transform 1 0 4092 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_262
timestamp 1677677812
transform 1 0 4100 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_411
timestamp 1677677812
transform 1 0 4108 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_312
timestamp 1677677812
transform 1 0 4092 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1677677812
transform 1 0 4156 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_255
timestamp 1677677812
transform 1 0 4180 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_256
timestamp 1677677812
transform 1 0 4196 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1677677812
transform 1 0 4188 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_264
timestamp 1677677812
transform 1 0 4196 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_257
timestamp 1677677812
transform 1 0 4236 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1677677812
transform 1 0 4228 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1677677812
transform 1 0 4244 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_313
timestamp 1677677812
transform 1 0 4228 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_415
timestamp 1677677812
transform 1 0 4260 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_258
timestamp 1677677812
transform 1 0 4268 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_265
timestamp 1677677812
transform 1 0 4268 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_259
timestamp 1677677812
transform 1 0 4300 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_416
timestamp 1677677812
transform 1 0 4292 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_314
timestamp 1677677812
transform 1 0 4292 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_188
timestamp 1677677812
transform 1 0 4308 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_260
timestamp 1677677812
transform 1 0 4308 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_148
timestamp 1677677812
transform 1 0 4348 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_189
timestamp 1677677812
transform 1 0 4340 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1677677812
transform 1 0 4324 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_261
timestamp 1677677812
transform 1 0 4332 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1677677812
transform 1 0 4348 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1677677812
transform 1 0 4324 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1677677812
transform 1 0 4340 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_266
timestamp 1677677812
transform 1 0 4348 0 1 4525
box -3 -3 3 3
use M2_M1  M2_M1_263
timestamp 1677677812
transform 1 0 4364 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_419
timestamp 1677677812
transform 1 0 4372 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_190
timestamp 1677677812
transform 1 0 4404 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_264
timestamp 1677677812
transform 1 0 4404 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_191
timestamp 1677677812
transform 1 0 4428 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_265
timestamp 1677677812
transform 1 0 4420 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1677677812
transform 1 0 4396 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1677677812
transform 1 0 4412 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_315
timestamp 1677677812
transform 1 0 4412 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_358
timestamp 1677677812
transform 1 0 4396 0 1 4485
box -3 -3 3 3
use M2_M1  M2_M1_422
timestamp 1677677812
transform 1 0 4428 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_224
timestamp 1677677812
transform 1 0 4444 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_423
timestamp 1677677812
transform 1 0 4444 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1677677812
transform 1 0 4460 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_129
timestamp 1677677812
transform 1 0 4572 0 1 4565
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1677677812
transform 1 0 4548 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1677677812
transform 1 0 4564 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1677677812
transform 1 0 4548 0 1 4545
box -3 -3 3 3
use M3_M2  M3_M2_225
timestamp 1677677812
transform 1 0 4524 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_267
timestamp 1677677812
transform 1 0 4532 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1677677812
transform 1 0 4548 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_269
timestamp 1677677812
transform 1 0 4564 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_226
timestamp 1677677812
transform 1 0 4596 0 1 4535
box -3 -3 3 3
use M2_M1  M2_M1_270
timestamp 1677677812
transform 1 0 4604 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1677677812
transform 1 0 4612 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1677677812
transform 1 0 4524 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1677677812
transform 1 0 4540 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1677677812
transform 1 0 4556 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_427
timestamp 1677677812
transform 1 0 4572 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1677677812
transform 1 0 4588 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1677677812
transform 1 0 4596 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_316
timestamp 1677677812
transform 1 0 4556 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1677677812
transform 1 0 4612 0 1 4495
box -3 -3 3 3
use M3_M2  M3_M2_347
timestamp 1677677812
transform 1 0 4628 0 1 4495
box -3 -3 3 3
use M2_M1  M2_M1_430
timestamp 1677677812
transform 1 0 4652 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_267
timestamp 1677677812
transform 1 0 4660 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_151
timestamp 1677677812
transform 1 0 4692 0 1 4555
box -3 -3 3 3
use M3_M2  M3_M2_193
timestamp 1677677812
transform 1 0 4700 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_272
timestamp 1677677812
transform 1 0 4684 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1677677812
transform 1 0 4700 0 1 4535
box -2 -2 2 2
use M2_M1  M2_M1_431
timestamp 1677677812
transform 1 0 4676 0 1 4525
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1677677812
transform 1 0 4692 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_268
timestamp 1677677812
transform 1 0 4700 0 1 4525
box -3 -3 3 3
use M3_M2  M3_M2_317
timestamp 1677677812
transform 1 0 4676 0 1 4515
box -3 -3 3 3
use M2_M1  M2_M1_433
timestamp 1677677812
transform 1 0 4724 0 1 4525
box -2 -2 2 2
use M3_M2  M3_M2_318
timestamp 1677677812
transform 1 0 4724 0 1 4515
box -3 -3 3 3
use M3_M2  M3_M2_194
timestamp 1677677812
transform 1 0 4740 0 1 4545
box -3 -3 3 3
use M2_M1  M2_M1_274
timestamp 1677677812
transform 1 0 4740 0 1 4535
box -2 -2 2 2
use M3_M2  M3_M2_152
timestamp 1677677812
transform 1 0 4780 0 1 4555
box -3 -3 3 3
use M2_M1  M2_M1_275
timestamp 1677677812
transform 1 0 4772 0 1 4535
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_4
timestamp 1677677812
transform 1 0 24 0 1 4470
box -10 -3 10 3
use FILL  FILL_1
timestamp 1677677812
transform 1 0 72 0 -1 4570
box -8 -3 16 105
use FILL  FILL_7
timestamp 1677677812
transform 1 0 80 0 -1 4570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1677677812
transform 1 0 88 0 -1 4570
box -8 -3 16 105
use FILL  FILL_9
timestamp 1677677812
transform 1 0 96 0 -1 4570
box -8 -3 16 105
use FILL  FILL_10
timestamp 1677677812
transform 1 0 104 0 -1 4570
box -8 -3 16 105
use FILL  FILL_11
timestamp 1677677812
transform 1 0 112 0 -1 4570
box -8 -3 16 105
use FILL  FILL_12
timestamp 1677677812
transform 1 0 120 0 -1 4570
box -8 -3 16 105
use FILL  FILL_13
timestamp 1677677812
transform 1 0 128 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1677677812
transform -1 0 152 0 -1 4570
box -9 -3 26 105
use FILL  FILL_14
timestamp 1677677812
transform 1 0 152 0 -1 4570
box -8 -3 16 105
use FILL  FILL_15
timestamp 1677677812
transform 1 0 160 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_0
timestamp 1677677812
transform -1 0 208 0 -1 4570
box -8 -3 46 105
use FILL  FILL_16
timestamp 1677677812
transform 1 0 208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_18
timestamp 1677677812
transform 1 0 216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_20
timestamp 1677677812
transform 1 0 224 0 -1 4570
box -8 -3 16 105
use FILL  FILL_22
timestamp 1677677812
transform 1 0 232 0 -1 4570
box -8 -3 16 105
use FILL  FILL_24
timestamp 1677677812
transform 1 0 240 0 -1 4570
box -8 -3 16 105
use FILL  FILL_26
timestamp 1677677812
transform 1 0 248 0 -1 4570
box -8 -3 16 105
use FILL  FILL_29
timestamp 1677677812
transform 1 0 256 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1677677812
transform 1 0 264 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_1
timestamp 1677677812
transform 1 0 304 0 -1 4570
box -9 -3 26 105
use FILL  FILL_30
timestamp 1677677812
transform 1 0 320 0 -1 4570
box -8 -3 16 105
use FILL  FILL_31
timestamp 1677677812
transform 1 0 328 0 -1 4570
box -8 -3 16 105
use FILL  FILL_32
timestamp 1677677812
transform 1 0 336 0 -1 4570
box -8 -3 16 105
use FILL  FILL_33
timestamp 1677677812
transform 1 0 344 0 -1 4570
box -8 -3 16 105
use FILL  FILL_34
timestamp 1677677812
transform 1 0 352 0 -1 4570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1677677812
transform 1 0 360 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1677677812
transform 1 0 368 0 -1 4570
box -9 -3 26 105
use AOI22X1  AOI22X1_2
timestamp 1677677812
transform -1 0 424 0 -1 4570
box -8 -3 46 105
use FILL  FILL_41
timestamp 1677677812
transform 1 0 424 0 -1 4570
box -8 -3 16 105
use FILL  FILL_42
timestamp 1677677812
transform 1 0 432 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_359
timestamp 1677677812
transform 1 0 452 0 1 4475
box -3 -3 3 3
use FILL  FILL_43
timestamp 1677677812
transform 1 0 440 0 -1 4570
box -8 -3 16 105
use FILL  FILL_44
timestamp 1677677812
transform 1 0 448 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_360
timestamp 1677677812
transform 1 0 484 0 1 4475
box -3 -3 3 3
use OAI22X1  OAI22X1_0
timestamp 1677677812
transform -1 0 496 0 -1 4570
box -8 -3 46 105
use FILL  FILL_45
timestamp 1677677812
transform 1 0 496 0 -1 4570
box -8 -3 16 105
use FILL  FILL_47
timestamp 1677677812
transform 1 0 504 0 -1 4570
box -8 -3 16 105
use FILL  FILL_49
timestamp 1677677812
transform 1 0 512 0 -1 4570
box -8 -3 16 105
use FILL  FILL_54
timestamp 1677677812
transform 1 0 520 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_3
timestamp 1677677812
transform -1 0 568 0 -1 4570
box -8 -3 46 105
use FILL  FILL_55
timestamp 1677677812
transform 1 0 568 0 -1 4570
box -8 -3 16 105
use FILL  FILL_56
timestamp 1677677812
transform 1 0 576 0 -1 4570
box -8 -3 16 105
use FILL  FILL_57
timestamp 1677677812
transform 1 0 584 0 -1 4570
box -8 -3 16 105
use FILL  FILL_58
timestamp 1677677812
transform 1 0 592 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_361
timestamp 1677677812
transform 1 0 612 0 1 4475
box -3 -3 3 3
use FILL  FILL_59
timestamp 1677677812
transform 1 0 600 0 -1 4570
box -8 -3 16 105
use FILL  FILL_60
timestamp 1677677812
transform 1 0 608 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_4
timestamp 1677677812
transform 1 0 616 0 -1 4570
box -8 -3 46 105
use FILL  FILL_61
timestamp 1677677812
transform 1 0 656 0 -1 4570
box -8 -3 16 105
use FILL  FILL_63
timestamp 1677677812
transform 1 0 664 0 -1 4570
box -8 -3 16 105
use FILL  FILL_65
timestamp 1677677812
transform 1 0 672 0 -1 4570
box -8 -3 16 105
use FILL  FILL_68
timestamp 1677677812
transform 1 0 680 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_1
timestamp 1677677812
transform -1 0 728 0 -1 4570
box -8 -3 46 105
use FILL  FILL_69
timestamp 1677677812
transform 1 0 728 0 -1 4570
box -8 -3 16 105
use FILL  FILL_70
timestamp 1677677812
transform 1 0 736 0 -1 4570
box -8 -3 16 105
use FILL  FILL_71
timestamp 1677677812
transform 1 0 744 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_5
timestamp 1677677812
transform 1 0 752 0 -1 4570
box -9 -3 26 105
use FILL  FILL_72
timestamp 1677677812
transform 1 0 768 0 -1 4570
box -8 -3 16 105
use FILL  FILL_73
timestamp 1677677812
transform 1 0 776 0 -1 4570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1677677812
transform 1 0 784 0 -1 4570
box -8 -3 104 105
use M3_M2  M3_M2_362
timestamp 1677677812
transform 1 0 892 0 1 4475
box -3 -3 3 3
use INVX2  INVX2_6
timestamp 1677677812
transform -1 0 896 0 -1 4570
box -9 -3 26 105
use FILL  FILL_74
timestamp 1677677812
transform 1 0 896 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_5
timestamp 1677677812
transform 1 0 904 0 -1 4570
box -8 -3 46 105
use FILL  FILL_81
timestamp 1677677812
transform 1 0 944 0 -1 4570
box -8 -3 16 105
use FILL  FILL_83
timestamp 1677677812
transform 1 0 952 0 -1 4570
box -8 -3 16 105
use FILL  FILL_85
timestamp 1677677812
transform 1 0 960 0 -1 4570
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1677677812
transform 1 0 968 0 -1 4570
box -8 -3 32 105
use FILL  FILL_90
timestamp 1677677812
transform 1 0 992 0 -1 4570
box -8 -3 16 105
use FILL  FILL_92
timestamp 1677677812
transform 1 0 1000 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_6
timestamp 1677677812
transform 1 0 1008 0 -1 4570
box -8 -3 46 105
use FILL  FILL_106
timestamp 1677677812
transform 1 0 1048 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_363
timestamp 1677677812
transform 1 0 1092 0 1 4475
box -3 -3 3 3
use OAI21X1  OAI21X1_0
timestamp 1677677812
transform 1 0 1056 0 -1 4570
box -8 -3 34 105
use FILL  FILL_107
timestamp 1677677812
transform 1 0 1088 0 -1 4570
box -8 -3 16 105
use FILL  FILL_108
timestamp 1677677812
transform 1 0 1096 0 -1 4570
box -8 -3 16 105
use FILL  FILL_109
timestamp 1677677812
transform 1 0 1104 0 -1 4570
box -8 -3 16 105
use FILL  FILL_110
timestamp 1677677812
transform 1 0 1112 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_7
timestamp 1677677812
transform 1 0 1120 0 -1 4570
box -8 -3 46 105
use OAI21X1  OAI21X1_1
timestamp 1677677812
transform 1 0 1160 0 -1 4570
box -8 -3 34 105
use INVX2  INVX2_8
timestamp 1677677812
transform 1 0 1192 0 -1 4570
box -9 -3 26 105
use FILL  FILL_111
timestamp 1677677812
transform 1 0 1208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_112
timestamp 1677677812
transform 1 0 1216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_113
timestamp 1677677812
transform 1 0 1224 0 -1 4570
box -8 -3 16 105
use FILL  FILL_114
timestamp 1677677812
transform 1 0 1232 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_364
timestamp 1677677812
transform 1 0 1276 0 1 4475
box -3 -3 3 3
use OAI21X1  OAI21X1_2
timestamp 1677677812
transform -1 0 1272 0 -1 4570
box -8 -3 34 105
use FILL  FILL_115
timestamp 1677677812
transform 1 0 1272 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1677677812
transform -1 0 1312 0 -1 4570
box -8 -3 34 105
use FILL  FILL_116
timestamp 1677677812
transform 1 0 1312 0 -1 4570
box -8 -3 16 105
use FILL  FILL_117
timestamp 1677677812
transform 1 0 1320 0 -1 4570
box -8 -3 16 105
use FILL  FILL_118
timestamp 1677677812
transform 1 0 1328 0 -1 4570
box -8 -3 16 105
use FILL  FILL_119
timestamp 1677677812
transform 1 0 1336 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_9
timestamp 1677677812
transform 1 0 1344 0 -1 4570
box -9 -3 26 105
use FILL  FILL_120
timestamp 1677677812
transform 1 0 1360 0 -1 4570
box -8 -3 16 105
use FILL  FILL_121
timestamp 1677677812
transform 1 0 1368 0 -1 4570
box -8 -3 16 105
use FILL  FILL_122
timestamp 1677677812
transform 1 0 1376 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_10
timestamp 1677677812
transform -1 0 1400 0 -1 4570
box -9 -3 26 105
use FILL  FILL_123
timestamp 1677677812
transform 1 0 1400 0 -1 4570
box -8 -3 16 105
use FILL  FILL_124
timestamp 1677677812
transform 1 0 1408 0 -1 4570
box -8 -3 16 105
use FILL  FILL_130
timestamp 1677677812
transform 1 0 1416 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_2
timestamp 1677677812
transform -1 0 1464 0 -1 4570
box -8 -3 46 105
use FILL  FILL_131
timestamp 1677677812
transform 1 0 1464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_132
timestamp 1677677812
transform 1 0 1472 0 -1 4570
box -8 -3 16 105
use FILL  FILL_133
timestamp 1677677812
transform 1 0 1480 0 -1 4570
box -8 -3 16 105
use FILL  FILL_134
timestamp 1677677812
transform 1 0 1488 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_3
timestamp 1677677812
transform -1 0 1536 0 -1 4570
box -8 -3 46 105
use FILL  FILL_135
timestamp 1677677812
transform 1 0 1536 0 -1 4570
box -8 -3 16 105
use FILL  FILL_136
timestamp 1677677812
transform 1 0 1544 0 -1 4570
box -8 -3 16 105
use FILL  FILL_138
timestamp 1677677812
transform 1 0 1552 0 -1 4570
box -8 -3 16 105
use FILL  FILL_140
timestamp 1677677812
transform 1 0 1560 0 -1 4570
box -8 -3 16 105
use FILL  FILL_142
timestamp 1677677812
transform 1 0 1568 0 -1 4570
box -8 -3 16 105
use FILL  FILL_159
timestamp 1677677812
transform 1 0 1576 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_12
timestamp 1677677812
transform 1 0 1584 0 -1 4570
box -9 -3 26 105
use OAI22X1  OAI22X1_4
timestamp 1677677812
transform -1 0 1640 0 -1 4570
box -8 -3 46 105
use FILL  FILL_160
timestamp 1677677812
transform 1 0 1640 0 -1 4570
box -8 -3 16 105
use FILL  FILL_161
timestamp 1677677812
transform 1 0 1648 0 -1 4570
box -8 -3 16 105
use FILL  FILL_162
timestamp 1677677812
transform 1 0 1656 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_13
timestamp 1677677812
transform -1 0 1680 0 -1 4570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1677677812
transform 1 0 1680 0 -1 4570
box -8 -3 104 105
use FILL  FILL_163
timestamp 1677677812
transform 1 0 1776 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_14
timestamp 1677677812
transform -1 0 1800 0 -1 4570
box -9 -3 26 105
use FILL  FILL_164
timestamp 1677677812
transform 1 0 1800 0 -1 4570
box -8 -3 16 105
use FILL  FILL_165
timestamp 1677677812
transform 1 0 1808 0 -1 4570
box -8 -3 16 105
use FILL  FILL_166
timestamp 1677677812
transform 1 0 1816 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_8
timestamp 1677677812
transform 1 0 1824 0 -1 4570
box -8 -3 46 105
use FILL  FILL_167
timestamp 1677677812
transform 1 0 1864 0 -1 4570
box -8 -3 16 105
use FILL  FILL_168
timestamp 1677677812
transform 1 0 1872 0 -1 4570
box -8 -3 16 105
use FILL  FILL_169
timestamp 1677677812
transform 1 0 1880 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_15
timestamp 1677677812
transform 1 0 1888 0 -1 4570
box -9 -3 26 105
use FILL  FILL_170
timestamp 1677677812
transform 1 0 1904 0 -1 4570
box -8 -3 16 105
use FILL  FILL_172
timestamp 1677677812
transform 1 0 1912 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_21
timestamp 1677677812
transform 1 0 1920 0 -1 4570
box -9 -3 26 105
use INVX2  INVX2_22
timestamp 1677677812
transform 1 0 1936 0 -1 4570
box -9 -3 26 105
use FILL  FILL_202
timestamp 1677677812
transform 1 0 1952 0 -1 4570
box -8 -3 16 105
use FILL  FILL_203
timestamp 1677677812
transform 1 0 1960 0 -1 4570
box -8 -3 16 105
use FILL  FILL_204
timestamp 1677677812
transform 1 0 1968 0 -1 4570
box -8 -3 16 105
use FILL  FILL_205
timestamp 1677677812
transform 1 0 1976 0 -1 4570
box -8 -3 16 105
use FILL  FILL_206
timestamp 1677677812
transform 1 0 1984 0 -1 4570
box -8 -3 16 105
use FILL  FILL_207
timestamp 1677677812
transform 1 0 1992 0 -1 4570
box -8 -3 16 105
use FILL  FILL_208
timestamp 1677677812
transform 1 0 2000 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_9
timestamp 1677677812
transform 1 0 2008 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_23
timestamp 1677677812
transform 1 0 2048 0 -1 4570
box -9 -3 26 105
use FILL  FILL_209
timestamp 1677677812
transform 1 0 2064 0 -1 4570
box -8 -3 16 105
use FILL  FILL_210
timestamp 1677677812
transform 1 0 2072 0 -1 4570
box -8 -3 16 105
use FILL  FILL_211
timestamp 1677677812
transform 1 0 2080 0 -1 4570
box -8 -3 16 105
use FILL  FILL_212
timestamp 1677677812
transform 1 0 2088 0 -1 4570
box -8 -3 16 105
use FILL  FILL_213
timestamp 1677677812
transform 1 0 2096 0 -1 4570
box -8 -3 16 105
use FILL  FILL_214
timestamp 1677677812
transform 1 0 2104 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_10
timestamp 1677677812
transform 1 0 2112 0 -1 4570
box -8 -3 46 105
use AOI22X1  AOI22X1_11
timestamp 1677677812
transform 1 0 2152 0 -1 4570
box -8 -3 46 105
use FILL  FILL_215
timestamp 1677677812
transform 1 0 2192 0 -1 4570
box -8 -3 16 105
use FILL  FILL_216
timestamp 1677677812
transform 1 0 2200 0 -1 4570
box -8 -3 16 105
use FILL  FILL_217
timestamp 1677677812
transform 1 0 2208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_218
timestamp 1677677812
transform 1 0 2216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_219
timestamp 1677677812
transform 1 0 2224 0 -1 4570
box -8 -3 16 105
use FILL  FILL_220
timestamp 1677677812
transform 1 0 2232 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_5
timestamp 1677677812
transform 1 0 2240 0 -1 4570
box -8 -3 46 105
use FILL  FILL_221
timestamp 1677677812
transform 1 0 2280 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_365
timestamp 1677677812
transform 1 0 2324 0 1 4475
box -3 -3 3 3
use AOI22X1  AOI22X1_12
timestamp 1677677812
transform -1 0 2328 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_24
timestamp 1677677812
transform 1 0 2328 0 -1 4570
box -9 -3 26 105
use FILL  FILL_222
timestamp 1677677812
transform 1 0 2344 0 -1 4570
box -8 -3 16 105
use FILL  FILL_223
timestamp 1677677812
transform 1 0 2352 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_6
timestamp 1677677812
transform 1 0 2360 0 -1 4570
box -8 -3 46 105
use AOI22X1  AOI22X1_13
timestamp 1677677812
transform -1 0 2440 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_25
timestamp 1677677812
transform 1 0 2440 0 -1 4570
box -9 -3 26 105
use FILL  FILL_224
timestamp 1677677812
transform 1 0 2456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_225
timestamp 1677677812
transform 1 0 2464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_226
timestamp 1677677812
transform 1 0 2472 0 -1 4570
box -8 -3 16 105
use FILL  FILL_227
timestamp 1677677812
transform 1 0 2480 0 -1 4570
box -8 -3 16 105
use FILL  FILL_228
timestamp 1677677812
transform 1 0 2488 0 -1 4570
box -8 -3 16 105
use FILL  FILL_229
timestamp 1677677812
transform 1 0 2496 0 -1 4570
box -8 -3 16 105
use FILL  FILL_230
timestamp 1677677812
transform 1 0 2504 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_14
timestamp 1677677812
transform 1 0 2512 0 -1 4570
box -8 -3 46 105
use FILL  FILL_231
timestamp 1677677812
transform 1 0 2552 0 -1 4570
box -8 -3 16 105
use FILL  FILL_232
timestamp 1677677812
transform 1 0 2560 0 -1 4570
box -8 -3 16 105
use FILL  FILL_233
timestamp 1677677812
transform 1 0 2568 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_26
timestamp 1677677812
transform 1 0 2576 0 -1 4570
box -9 -3 26 105
use FILL  FILL_234
timestamp 1677677812
transform 1 0 2592 0 -1 4570
box -8 -3 16 105
use FILL  FILL_235
timestamp 1677677812
transform 1 0 2600 0 -1 4570
box -8 -3 16 105
use FILL  FILL_236
timestamp 1677677812
transform 1 0 2608 0 -1 4570
box -8 -3 16 105
use FILL  FILL_237
timestamp 1677677812
transform 1 0 2616 0 -1 4570
box -8 -3 16 105
use FILL  FILL_238
timestamp 1677677812
transform 1 0 2624 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_15
timestamp 1677677812
transform 1 0 2632 0 -1 4570
box -8 -3 46 105
use M3_M2  M3_M2_366
timestamp 1677677812
transform 1 0 2716 0 1 4475
box -3 -3 3 3
use AOI22X1  AOI22X1_16
timestamp 1677677812
transform 1 0 2672 0 -1 4570
box -8 -3 46 105
use AOI22X1  AOI22X1_17
timestamp 1677677812
transform 1 0 2712 0 -1 4570
box -8 -3 46 105
use FILL  FILL_239
timestamp 1677677812
transform 1 0 2752 0 -1 4570
box -8 -3 16 105
use FILL  FILL_240
timestamp 1677677812
transform 1 0 2760 0 -1 4570
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1677677812
transform 1 0 2768 0 -1 4570
box -8 -3 32 105
use FILL  FILL_241
timestamp 1677677812
transform 1 0 2792 0 -1 4570
box -8 -3 16 105
use FILL  FILL_242
timestamp 1677677812
transform 1 0 2800 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_5
timestamp 1677677812
transform 1 0 2808 0 -1 4570
box -8 -3 34 105
use NOR2X1  NOR2X1_2
timestamp 1677677812
transform 1 0 2840 0 -1 4570
box -8 -3 32 105
use FILL  FILL_243
timestamp 1677677812
transform 1 0 2864 0 -1 4570
box -8 -3 16 105
use FILL  FILL_244
timestamp 1677677812
transform 1 0 2872 0 -1 4570
box -8 -3 16 105
use FILL  FILL_245
timestamp 1677677812
transform 1 0 2880 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1677677812
transform 1 0 2888 0 -1 4570
box -8 -3 34 105
use FILL  FILL_246
timestamp 1677677812
transform 1 0 2920 0 -1 4570
box -8 -3 16 105
use FILL  FILL_247
timestamp 1677677812
transform 1 0 2928 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_367
timestamp 1677677812
transform 1 0 2964 0 1 4475
box -3 -3 3 3
use OAI21X1  OAI21X1_7
timestamp 1677677812
transform -1 0 2968 0 -1 4570
box -8 -3 34 105
use FILL  FILL_248
timestamp 1677677812
transform 1 0 2968 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_368
timestamp 1677677812
transform 1 0 3012 0 1 4475
box -3 -3 3 3
use OAI21X1  OAI21X1_8
timestamp 1677677812
transform -1 0 3008 0 -1 4570
box -8 -3 34 105
use FILL  FILL_249
timestamp 1677677812
transform 1 0 3008 0 -1 4570
box -8 -3 16 105
use FILL  FILL_250
timestamp 1677677812
transform 1 0 3016 0 -1 4570
box -8 -3 16 105
use FILL  FILL_251
timestamp 1677677812
transform 1 0 3024 0 -1 4570
box -8 -3 16 105
use FILL  FILL_252
timestamp 1677677812
transform 1 0 3032 0 -1 4570
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1677677812
transform -1 0 3072 0 -1 4570
box -8 -3 34 105
use FILL  FILL_253
timestamp 1677677812
transform 1 0 3072 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_7
timestamp 1677677812
transform -1 0 3120 0 -1 4570
box -8 -3 46 105
use FILL  FILL_254
timestamp 1677677812
transform 1 0 3120 0 -1 4570
box -8 -3 16 105
use FILL  FILL_256
timestamp 1677677812
transform 1 0 3128 0 -1 4570
box -8 -3 16 105
use FILL  FILL_257
timestamp 1677677812
transform 1 0 3136 0 -1 4570
box -8 -3 16 105
use FILL  FILL_258
timestamp 1677677812
transform 1 0 3144 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_8
timestamp 1677677812
transform 1 0 3152 0 -1 4570
box -8 -3 46 105
use FILL  FILL_259
timestamp 1677677812
transform 1 0 3192 0 -1 4570
box -8 -3 16 105
use FILL  FILL_260
timestamp 1677677812
transform 1 0 3200 0 -1 4570
box -8 -3 16 105
use FILL  FILL_261
timestamp 1677677812
transform 1 0 3208 0 -1 4570
box -8 -3 16 105
use FILL  FILL_262
timestamp 1677677812
transform 1 0 3216 0 -1 4570
box -8 -3 16 105
use FILL  FILL_263
timestamp 1677677812
transform 1 0 3224 0 -1 4570
box -8 -3 16 105
use FILL  FILL_272
timestamp 1677677812
transform 1 0 3232 0 -1 4570
box -8 -3 16 105
use FILL  FILL_273
timestamp 1677677812
transform 1 0 3240 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_9
timestamp 1677677812
transform -1 0 3288 0 -1 4570
box -8 -3 46 105
use INVX2  INVX2_29
timestamp 1677677812
transform -1 0 3304 0 -1 4570
box -9 -3 26 105
use FILL  FILL_274
timestamp 1677677812
transform 1 0 3304 0 -1 4570
box -8 -3 16 105
use FILL  FILL_275
timestamp 1677677812
transform 1 0 3312 0 -1 4570
box -8 -3 16 105
use FILL  FILL_276
timestamp 1677677812
transform 1 0 3320 0 -1 4570
box -8 -3 16 105
use FILL  FILL_277
timestamp 1677677812
transform 1 0 3328 0 -1 4570
box -8 -3 16 105
use FILL  FILL_278
timestamp 1677677812
transform 1 0 3336 0 -1 4570
box -8 -3 16 105
use FILL  FILL_279
timestamp 1677677812
transform 1 0 3344 0 -1 4570
box -8 -3 16 105
use FILL  FILL_280
timestamp 1677677812
transform 1 0 3352 0 -1 4570
box -8 -3 16 105
use FILL  FILL_281
timestamp 1677677812
transform 1 0 3360 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_30
timestamp 1677677812
transform 1 0 3368 0 -1 4570
box -9 -3 26 105
use FILL  FILL_282
timestamp 1677677812
transform 1 0 3384 0 -1 4570
box -8 -3 16 105
use FILL  FILL_283
timestamp 1677677812
transform 1 0 3392 0 -1 4570
box -8 -3 16 105
use FILL  FILL_284
timestamp 1677677812
transform 1 0 3400 0 -1 4570
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1677677812
transform -1 0 3440 0 -1 4570
box -8 -3 40 105
use FILL  FILL_285
timestamp 1677677812
transform 1 0 3440 0 -1 4570
box -8 -3 16 105
use FILL  FILL_286
timestamp 1677677812
transform 1 0 3448 0 -1 4570
box -8 -3 16 105
use FILL  FILL_287
timestamp 1677677812
transform 1 0 3456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_288
timestamp 1677677812
transform 1 0 3464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_289
timestamp 1677677812
transform 1 0 3472 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_369
timestamp 1677677812
transform 1 0 3492 0 1 4475
box -3 -3 3 3
use FILL  FILL_290
timestamp 1677677812
transform 1 0 3480 0 -1 4570
box -8 -3 16 105
use FILL  FILL_291
timestamp 1677677812
transform 1 0 3488 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_10
timestamp 1677677812
transform 1 0 3496 0 -1 4570
box -8 -3 46 105
use FILL  FILL_292
timestamp 1677677812
transform 1 0 3536 0 -1 4570
box -8 -3 16 105
use FILL  FILL_293
timestamp 1677677812
transform 1 0 3544 0 -1 4570
box -8 -3 16 105
use FILL  FILL_294
timestamp 1677677812
transform 1 0 3552 0 -1 4570
box -8 -3 16 105
use FILL  FILL_295
timestamp 1677677812
transform 1 0 3560 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_18
timestamp 1677677812
transform -1 0 3608 0 -1 4570
box -8 -3 46 105
use FILL  FILL_296
timestamp 1677677812
transform 1 0 3608 0 -1 4570
box -8 -3 16 105
use FILL  FILL_300
timestamp 1677677812
transform 1 0 3616 0 -1 4570
box -8 -3 16 105
use FILL  FILL_301
timestamp 1677677812
transform 1 0 3624 0 -1 4570
box -8 -3 16 105
use FILL  FILL_302
timestamp 1677677812
transform 1 0 3632 0 -1 4570
box -8 -3 16 105
use FILL  FILL_303
timestamp 1677677812
transform 1 0 3640 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_19
timestamp 1677677812
transform -1 0 3688 0 -1 4570
box -8 -3 46 105
use FILL  FILL_304
timestamp 1677677812
transform 1 0 3688 0 -1 4570
box -8 -3 16 105
use FILL  FILL_305
timestamp 1677677812
transform 1 0 3696 0 -1 4570
box -8 -3 16 105
use FILL  FILL_306
timestamp 1677677812
transform 1 0 3704 0 -1 4570
box -8 -3 16 105
use FILL  FILL_307
timestamp 1677677812
transform 1 0 3712 0 -1 4570
box -8 -3 16 105
use FILL  FILL_308
timestamp 1677677812
transform 1 0 3720 0 -1 4570
box -8 -3 16 105
use M3_M2  M3_M2_370
timestamp 1677677812
transform 1 0 3740 0 1 4475
box -3 -3 3 3
use FILL  FILL_309
timestamp 1677677812
transform 1 0 3728 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_12
timestamp 1677677812
transform 1 0 3736 0 -1 4570
box -8 -3 46 105
use FILL  FILL_310
timestamp 1677677812
transform 1 0 3776 0 -1 4570
box -8 -3 16 105
use FILL  FILL_311
timestamp 1677677812
transform 1 0 3784 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_13
timestamp 1677677812
transform 1 0 3792 0 -1 4570
box -8 -3 46 105
use FILL  FILL_315
timestamp 1677677812
transform 1 0 3832 0 -1 4570
box -8 -3 16 105
use FILL  FILL_316
timestamp 1677677812
transform 1 0 3840 0 -1 4570
box -8 -3 16 105
use FILL  FILL_317
timestamp 1677677812
transform 1 0 3848 0 -1 4570
box -8 -3 16 105
use FILL  FILL_318
timestamp 1677677812
transform 1 0 3856 0 -1 4570
box -8 -3 16 105
use FILL  FILL_319
timestamp 1677677812
transform 1 0 3864 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_32
timestamp 1677677812
transform -1 0 3888 0 -1 4570
box -9 -3 26 105
use FILL  FILL_320
timestamp 1677677812
transform 1 0 3888 0 -1 4570
box -8 -3 16 105
use FILL  FILL_321
timestamp 1677677812
transform 1 0 3896 0 -1 4570
box -8 -3 16 105
use FILL  FILL_322
timestamp 1677677812
transform 1 0 3904 0 -1 4570
box -8 -3 16 105
use FILL  FILL_332
timestamp 1677677812
transform 1 0 3912 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_14
timestamp 1677677812
transform -1 0 3960 0 -1 4570
box -8 -3 46 105
use FILL  FILL_333
timestamp 1677677812
transform 1 0 3960 0 -1 4570
box -8 -3 16 105
use FILL  FILL_334
timestamp 1677677812
transform 1 0 3968 0 -1 4570
box -8 -3 16 105
use FILL  FILL_335
timestamp 1677677812
transform 1 0 3976 0 -1 4570
box -8 -3 16 105
use FILL  FILL_336
timestamp 1677677812
transform 1 0 3984 0 -1 4570
box -8 -3 16 105
use FILL  FILL_337
timestamp 1677677812
transform 1 0 3992 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_15
timestamp 1677677812
transform 1 0 4000 0 -1 4570
box -8 -3 46 105
use FILL  FILL_338
timestamp 1677677812
transform 1 0 4040 0 -1 4570
box -8 -3 16 105
use FILL  FILL_339
timestamp 1677677812
transform 1 0 4048 0 -1 4570
box -8 -3 16 105
use FILL  FILL_340
timestamp 1677677812
transform 1 0 4056 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_16
timestamp 1677677812
transform -1 0 4104 0 -1 4570
box -8 -3 46 105
use FILL  FILL_341
timestamp 1677677812
transform 1 0 4104 0 -1 4570
box -8 -3 16 105
use FILL  FILL_342
timestamp 1677677812
transform 1 0 4112 0 -1 4570
box -8 -3 16 105
use FILL  FILL_343
timestamp 1677677812
transform 1 0 4120 0 -1 4570
box -8 -3 16 105
use FILL  FILL_344
timestamp 1677677812
transform 1 0 4128 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_34
timestamp 1677677812
transform -1 0 4152 0 -1 4570
box -9 -3 26 105
use FILL  FILL_345
timestamp 1677677812
transform 1 0 4152 0 -1 4570
box -8 -3 16 105
use FILL  FILL_346
timestamp 1677677812
transform 1 0 4160 0 -1 4570
box -8 -3 16 105
use FILL  FILL_347
timestamp 1677677812
transform 1 0 4168 0 -1 4570
box -8 -3 16 105
use FILL  FILL_348
timestamp 1677677812
transform 1 0 4176 0 -1 4570
box -8 -3 16 105
use FILL  FILL_349
timestamp 1677677812
transform 1 0 4184 0 -1 4570
box -8 -3 16 105
use FILL  FILL_351
timestamp 1677677812
transform 1 0 4192 0 -1 4570
box -8 -3 16 105
use FILL  FILL_353
timestamp 1677677812
transform 1 0 4200 0 -1 4570
box -8 -3 16 105
use FILL  FILL_355
timestamp 1677677812
transform 1 0 4208 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_17
timestamp 1677677812
transform 1 0 4216 0 -1 4570
box -8 -3 46 105
use FILL  FILL_356
timestamp 1677677812
transform 1 0 4256 0 -1 4570
box -8 -3 16 105
use FILL  FILL_357
timestamp 1677677812
transform 1 0 4264 0 -1 4570
box -8 -3 16 105
use FILL  FILL_358
timestamp 1677677812
transform 1 0 4272 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_35
timestamp 1677677812
transform -1 0 4296 0 -1 4570
box -9 -3 26 105
use FILL  FILL_359
timestamp 1677677812
transform 1 0 4296 0 -1 4570
box -8 -3 16 105
use FILL  FILL_360
timestamp 1677677812
transform 1 0 4304 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_18
timestamp 1677677812
transform 1 0 4312 0 -1 4570
box -8 -3 46 105
use FILL  FILL_371
timestamp 1677677812
transform 1 0 4352 0 -1 4570
box -8 -3 16 105
use FILL  FILL_372
timestamp 1677677812
transform 1 0 4360 0 -1 4570
box -8 -3 16 105
use FILL  FILL_373
timestamp 1677677812
transform 1 0 4368 0 -1 4570
box -8 -3 16 105
use AOI22X1  AOI22X1_20
timestamp 1677677812
transform -1 0 4416 0 -1 4570
box -8 -3 46 105
use FILL  FILL_374
timestamp 1677677812
transform 1 0 4416 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_37
timestamp 1677677812
transform 1 0 4424 0 -1 4570
box -9 -3 26 105
use FILL  FILL_375
timestamp 1677677812
transform 1 0 4440 0 -1 4570
box -8 -3 16 105
use FILL  FILL_376
timestamp 1677677812
transform 1 0 4448 0 -1 4570
box -8 -3 16 105
use FILL  FILL_377
timestamp 1677677812
transform 1 0 4456 0 -1 4570
box -8 -3 16 105
use FILL  FILL_378
timestamp 1677677812
transform 1 0 4464 0 -1 4570
box -8 -3 16 105
use FILL  FILL_379
timestamp 1677677812
transform 1 0 4472 0 -1 4570
box -8 -3 16 105
use FILL  FILL_380
timestamp 1677677812
transform 1 0 4480 0 -1 4570
box -8 -3 16 105
use FILL  FILL_381
timestamp 1677677812
transform 1 0 4488 0 -1 4570
box -8 -3 16 105
use FILL  FILL_382
timestamp 1677677812
transform 1 0 4496 0 -1 4570
box -8 -3 16 105
use FILL  FILL_383
timestamp 1677677812
transform 1 0 4504 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_19
timestamp 1677677812
transform 1 0 4512 0 -1 4570
box -8 -3 46 105
use AOI22X1  AOI22X1_21
timestamp 1677677812
transform 1 0 4552 0 -1 4570
box -8 -3 46 105
use FILL  FILL_384
timestamp 1677677812
transform 1 0 4592 0 -1 4570
box -8 -3 16 105
use FILL  FILL_386
timestamp 1677677812
transform 1 0 4600 0 -1 4570
box -8 -3 16 105
use FILL  FILL_388
timestamp 1677677812
transform 1 0 4608 0 -1 4570
box -8 -3 16 105
use FILL  FILL_390
timestamp 1677677812
transform 1 0 4616 0 -1 4570
box -8 -3 16 105
use FILL  FILL_392
timestamp 1677677812
transform 1 0 4624 0 -1 4570
box -8 -3 16 105
use FILL  FILL_394
timestamp 1677677812
transform 1 0 4632 0 -1 4570
box -8 -3 16 105
use FILL  FILL_396
timestamp 1677677812
transform 1 0 4640 0 -1 4570
box -8 -3 16 105
use FILL  FILL_398
timestamp 1677677812
transform 1 0 4648 0 -1 4570
box -8 -3 16 105
use FILL  FILL_400
timestamp 1677677812
transform 1 0 4656 0 -1 4570
box -8 -3 16 105
use OAI22X1  OAI22X1_20
timestamp 1677677812
transform 1 0 4664 0 -1 4570
box -8 -3 46 105
use FILL  FILL_403
timestamp 1677677812
transform 1 0 4704 0 -1 4570
box -8 -3 16 105
use FILL  FILL_404
timestamp 1677677812
transform 1 0 4712 0 -1 4570
box -8 -3 16 105
use FILL  FILL_405
timestamp 1677677812
transform 1 0 4720 0 -1 4570
box -8 -3 16 105
use INVX2  INVX2_39
timestamp 1677677812
transform -1 0 4744 0 -1 4570
box -9 -3 26 105
use FILL  FILL_406
timestamp 1677677812
transform 1 0 4744 0 -1 4570
box -8 -3 16 105
use FILL  FILL_407
timestamp 1677677812
transform 1 0 4752 0 -1 4570
box -8 -3 16 105
use FILL  FILL_408
timestamp 1677677812
transform 1 0 4760 0 -1 4570
box -8 -3 16 105
use FILL  FILL_409
timestamp 1677677812
transform 1 0 4768 0 -1 4570
box -8 -3 16 105
use FILL  FILL_410
timestamp 1677677812
transform 1 0 4776 0 -1 4570
box -8 -3 16 105
use FILL  FILL_411
timestamp 1677677812
transform 1 0 4784 0 -1 4570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_5
timestamp 1677677812
transform 1 0 4843 0 1 4470
box -10 -3 10 3
use M3_M2  M3_M2_398
timestamp 1677677812
transform 1 0 164 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_423
timestamp 1677677812
transform 1 0 132 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_424
timestamp 1677677812
transform 1 0 172 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_472
timestamp 1677677812
transform 1 0 124 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_464
timestamp 1677677812
transform 1 0 132 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_465
timestamp 1677677812
transform 1 0 164 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1677677812
transform 1 0 172 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_582
timestamp 1677677812
transform 1 0 84 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_390
timestamp 1677677812
transform 1 0 220 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1677677812
transform 1 0 196 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_467
timestamp 1677677812
transform 1 0 180 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1677677812
transform 1 0 204 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_473
timestamp 1677677812
transform 1 0 212 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_469
timestamp 1677677812
transform 1 0 220 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_583
timestamp 1677677812
transform 1 0 188 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_584
timestamp 1677677812
transform 1 0 196 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1677677812
transform 1 0 220 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_586
timestamp 1677677812
transform 1 0 228 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_512
timestamp 1677677812
transform 1 0 220 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_400
timestamp 1677677812
transform 1 0 268 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1677677812
transform 1 0 260 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_470
timestamp 1677677812
transform 1 0 244 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1677677812
transform 1 0 260 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_587
timestamp 1677677812
transform 1 0 252 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_492
timestamp 1677677812
transform 1 0 260 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_588
timestamp 1677677812
transform 1 0 268 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_426
timestamp 1677677812
transform 1 0 284 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_474
timestamp 1677677812
transform 1 0 332 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_472
timestamp 1677677812
transform 1 0 388 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_427
timestamp 1677677812
transform 1 0 452 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1677677812
transform 1 0 484 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_473
timestamp 1677677812
transform 1 0 452 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1677677812
transform 1 0 460 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_474
timestamp 1677677812
transform 1 0 468 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1677677812
transform 1 0 484 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1677677812
transform 1 0 452 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1677677812
transform 1 0 460 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1677677812
transform 1 0 476 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1677677812
transform 1 0 476 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_476
timestamp 1677677812
transform 1 0 500 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1677677812
transform 1 0 556 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1677677812
transform 1 0 524 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1677677812
transform 1 0 532 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1677677812
transform 1 0 548 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1677677812
transform 1 0 564 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1677677812
transform 1 0 572 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_514
timestamp 1677677812
transform 1 0 548 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_371
timestamp 1677677812
transform 1 0 588 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_428
timestamp 1677677812
transform 1 0 580 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_535
timestamp 1677677812
transform 1 0 572 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_478
timestamp 1677677812
transform 1 0 596 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_536
timestamp 1677677812
transform 1 0 588 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_429
timestamp 1677677812
transform 1 0 644 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_479
timestamp 1677677812
transform 1 0 612 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1677677812
transform 1 0 628 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_476
timestamp 1677677812
transform 1 0 636 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_481
timestamp 1677677812
transform 1 0 644 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1677677812
transform 1 0 620 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_537
timestamp 1677677812
transform 1 0 628 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_477
timestamp 1677677812
transform 1 0 660 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_482
timestamp 1677677812
transform 1 0 692 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_391
timestamp 1677677812
transform 1 0 756 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_483
timestamp 1677677812
transform 1 0 756 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_598
timestamp 1677677812
transform 1 0 780 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_493
timestamp 1677677812
transform 1 0 796 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_686
timestamp 1677677812
transform 1 0 796 0 1 4395
box -2 -2 2 2
use M3_M2  M3_M2_392
timestamp 1677677812
transform 1 0 884 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1677677812
transform 1 0 868 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_484
timestamp 1677677812
transform 1 0 860 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_485
timestamp 1677677812
transform 1 0 868 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1677677812
transform 1 0 884 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1677677812
transform 1 0 892 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_599
timestamp 1677677812
transform 1 0 868 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_600
timestamp 1677677812
transform 1 0 876 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1677677812
transform 1 0 892 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_602
timestamp 1677677812
transform 1 0 900 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_538
timestamp 1677677812
transform 1 0 860 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_603
timestamp 1677677812
transform 1 0 916 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_430
timestamp 1677677812
transform 1 0 956 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_487
timestamp 1677677812
transform 1 0 940 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_479
timestamp 1677677812
transform 1 0 948 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_488
timestamp 1677677812
transform 1 0 956 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_604
timestamp 1677677812
transform 1 0 948 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_605
timestamp 1677677812
transform 1 0 972 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_539
timestamp 1677677812
transform 1 0 972 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_687
timestamp 1677677812
transform 1 0 980 0 1 4395
box -2 -2 2 2
use M3_M2  M3_M2_383
timestamp 1677677812
transform 1 0 1012 0 1 4455
box -3 -3 3 3
use M2_M1  M2_M1_448
timestamp 1677677812
transform 1 0 1004 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_606
timestamp 1677677812
transform 1 0 1012 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1677677812
transform 1 0 1036 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_480
timestamp 1677677812
transform 1 0 1044 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_372
timestamp 1677677812
transform 1 0 1084 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1677677812
transform 1 0 1108 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_449
timestamp 1677677812
transform 1 0 1092 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1677677812
transform 1 0 1100 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_431
timestamp 1677677812
transform 1 0 1116 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_490
timestamp 1677677812
transform 1 0 1052 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_491
timestamp 1677677812
transform 1 0 1068 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_481
timestamp 1677677812
transform 1 0 1092 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1677677812
transform 1 0 1108 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_492
timestamp 1677677812
transform 1 0 1116 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_607
timestamp 1677677812
transform 1 0 1044 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_688
timestamp 1677677812
transform 1 0 1028 0 1 4395
box -2 -2 2 2
use M3_M2  M3_M2_494
timestamp 1677677812
transform 1 0 1052 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_608
timestamp 1677677812
transform 1 0 1060 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_495
timestamp 1677677812
transform 1 0 1076 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_609
timestamp 1677677812
transform 1 0 1084 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_610
timestamp 1677677812
transform 1 0 1092 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_540
timestamp 1677677812
transform 1 0 1100 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_611
timestamp 1677677812
transform 1 0 1132 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_496
timestamp 1677677812
transform 1 0 1140 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_612
timestamp 1677677812
transform 1 0 1148 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1677677812
transform 1 0 1140 0 1 4395
box -2 -2 2 2
use M2_M1  M2_M1_493
timestamp 1677677812
transform 1 0 1180 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_494
timestamp 1677677812
transform 1 0 1188 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_403
timestamp 1677677812
transform 1 0 1236 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_451
timestamp 1677677812
transform 1 0 1236 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_393
timestamp 1677677812
transform 1 0 1300 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1677677812
transform 1 0 1268 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_405
timestamp 1677677812
transform 1 0 1292 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_452
timestamp 1677677812
transform 1 0 1268 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_453
timestamp 1677677812
transform 1 0 1300 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1677677812
transform 1 0 1268 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_496
timestamp 1677677812
transform 1 0 1284 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1677677812
transform 1 0 1260 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_614
timestamp 1677677812
transform 1 0 1268 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_497
timestamp 1677677812
transform 1 0 1284 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_432
timestamp 1677677812
transform 1 0 1308 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_433
timestamp 1677677812
transform 1 0 1324 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_497
timestamp 1677677812
transform 1 0 1316 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1677677812
transform 1 0 1292 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1677677812
transform 1 0 1300 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_498
timestamp 1677677812
transform 1 0 1316 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_498
timestamp 1677677812
transform 1 0 1388 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1677677812
transform 1 0 1324 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_618
timestamp 1677677812
transform 1 0 1340 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_541
timestamp 1677677812
transform 1 0 1300 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1677677812
transform 1 0 1388 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1677677812
transform 1 0 1436 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_499
timestamp 1677677812
transform 1 0 1436 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1677677812
transform 1 0 1468 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_435
timestamp 1677677812
transform 1 0 1484 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_500
timestamp 1677677812
transform 1 0 1484 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1677677812
transform 1 0 1492 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_516
timestamp 1677677812
transform 1 0 1492 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_501
timestamp 1677677812
transform 1 0 1516 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1677677812
transform 1 0 1532 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_406
timestamp 1677677812
transform 1 0 1644 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1677677812
transform 1 0 1628 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_502
timestamp 1677677812
transform 1 0 1596 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1677677812
transform 1 0 1548 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_517
timestamp 1677677812
transform 1 0 1596 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_503
timestamp 1677677812
transform 1 0 1644 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_623
timestamp 1677677812
transform 1 0 1652 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_407
timestamp 1677677812
transform 1 0 1692 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_437
timestamp 1677677812
transform 1 0 1708 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_504
timestamp 1677677812
transform 1 0 1692 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_505
timestamp 1677677812
transform 1 0 1708 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1677677812
transform 1 0 1700 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_518
timestamp 1677677812
transform 1 0 1700 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_483
timestamp 1677677812
transform 1 0 1724 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_625
timestamp 1677677812
transform 1 0 1724 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_438
timestamp 1677677812
transform 1 0 1748 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_506
timestamp 1677677812
transform 1 0 1748 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_507
timestamp 1677677812
transform 1 0 1756 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1677677812
transform 1 0 1740 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_439
timestamp 1677677812
transform 1 0 1772 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1677677812
transform 1 0 1812 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1677677812
transform 1 0 1836 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1677677812
transform 1 0 1828 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_508
timestamp 1677677812
transform 1 0 1804 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_509
timestamp 1677677812
transform 1 0 1820 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1677677812
transform 1 0 1812 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1677677812
transform 1 0 1828 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_519
timestamp 1677677812
transform 1 0 1804 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_510
timestamp 1677677812
transform 1 0 1860 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_373
timestamp 1677677812
transform 1 0 1892 0 1 4465
box -3 -3 3 3
use M2_M1  M2_M1_511
timestamp 1677677812
transform 1 0 1892 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_512
timestamp 1677677812
transform 1 0 1908 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1677677812
transform 1 0 1900 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_441
timestamp 1677677812
transform 1 0 1996 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_513
timestamp 1677677812
transform 1 0 1988 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_514
timestamp 1677677812
transform 1 0 2004 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_499
timestamp 1677677812
transform 1 0 1988 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_442
timestamp 1677677812
transform 1 0 2028 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_515
timestamp 1677677812
transform 1 0 2028 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_630
timestamp 1677677812
transform 1 0 1996 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_631
timestamp 1677677812
transform 1 0 2012 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1677677812
transform 1 0 2020 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_500
timestamp 1677677812
transform 1 0 2028 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1677677812
transform 1 0 2020 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_374
timestamp 1677677812
transform 1 0 2084 0 1 4465
box -3 -3 3 3
use M2_M1  M2_M1_516
timestamp 1677677812
transform 1 0 2068 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_501
timestamp 1677677812
transform 1 0 2044 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_502
timestamp 1677677812
transform 1 0 2068 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_633
timestamp 1677677812
transform 1 0 2116 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_521
timestamp 1677677812
transform 1 0 2036 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_443
timestamp 1677677812
transform 1 0 2188 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_410
timestamp 1677677812
transform 1 0 2260 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1677677812
transform 1 0 2252 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_517
timestamp 1677677812
transform 1 0 2164 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1677677812
transform 1 0 2220 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_519
timestamp 1677677812
transform 1 0 2236 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_520
timestamp 1677677812
transform 1 0 2252 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1677677812
transform 1 0 2140 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1677677812
transform 1 0 2228 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_636
timestamp 1677677812
transform 1 0 2244 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_522
timestamp 1677677812
transform 1 0 2228 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_445
timestamp 1677677812
transform 1 0 2268 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_637
timestamp 1677677812
transform 1 0 2268 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1677677812
transform 1 0 2276 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_542
timestamp 1677677812
transform 1 0 2276 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_446
timestamp 1677677812
transform 1 0 2292 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_521
timestamp 1677677812
transform 1 0 2292 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_384
timestamp 1677677812
transform 1 0 2316 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_447
timestamp 1677677812
transform 1 0 2332 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_522
timestamp 1677677812
transform 1 0 2332 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1677677812
transform 1 0 2388 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1677677812
transform 1 0 2308 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1677677812
transform 1 0 2396 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_543
timestamp 1677677812
transform 1 0 2324 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_375
timestamp 1677677812
transform 1 0 2436 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_376
timestamp 1677677812
transform 1 0 2500 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1677677812
transform 1 0 2428 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_448
timestamp 1677677812
transform 1 0 2420 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_449
timestamp 1677677812
transform 1 0 2460 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_524
timestamp 1677677812
transform 1 0 2420 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1677677812
transform 1 0 2428 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_526
timestamp 1677677812
transform 1 0 2460 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1677677812
transform 1 0 2508 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_642
timestamp 1677677812
transform 1 0 2540 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_450
timestamp 1677677812
transform 1 0 2564 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_527
timestamp 1677677812
transform 1 0 2564 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_451
timestamp 1677677812
transform 1 0 2604 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_528
timestamp 1677677812
transform 1 0 2604 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1677677812
transform 1 0 2660 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1677677812
transform 1 0 2580 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_503
timestamp 1677677812
transform 1 0 2644 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_544
timestamp 1677677812
transform 1 0 2660 0 1 4385
box -3 -3 3 3
use M2_M1  M2_M1_644
timestamp 1677677812
transform 1 0 2684 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_452
timestamp 1677677812
transform 1 0 2700 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_530
timestamp 1677677812
transform 1 0 2700 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_453
timestamp 1677677812
transform 1 0 2740 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_531
timestamp 1677677812
transform 1 0 2740 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1677677812
transform 1 0 2796 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1677677812
transform 1 0 2716 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_646
timestamp 1677677812
transform 1 0 2804 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_545
timestamp 1677677812
transform 1 0 2804 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1677677812
transform 1 0 2828 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_533
timestamp 1677677812
transform 1 0 2828 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_411
timestamp 1677677812
transform 1 0 2852 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_647
timestamp 1677677812
transform 1 0 2852 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1677677812
transform 1 0 2860 0 1 4395
box -2 -2 2 2
use M3_M2  M3_M2_412
timestamp 1677677812
transform 1 0 2876 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_454
timestamp 1677677812
transform 1 0 2876 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_394
timestamp 1677677812
transform 1 0 2900 0 1 4445
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1677677812
transform 1 0 2916 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_534
timestamp 1677677812
transform 1 0 2908 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1677677812
transform 1 0 2916 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1677677812
transform 1 0 2932 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_648
timestamp 1677677812
transform 1 0 2900 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_649
timestamp 1677677812
transform 1 0 2908 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_504
timestamp 1677677812
transform 1 0 2916 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_455
timestamp 1677677812
transform 1 0 2964 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_650
timestamp 1677677812
transform 1 0 2964 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_386
timestamp 1677677812
transform 1 0 2996 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_413
timestamp 1677677812
transform 1 0 3004 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_456
timestamp 1677677812
transform 1 0 2972 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_456
timestamp 1677677812
transform 1 0 2988 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_537
timestamp 1677677812
transform 1 0 2988 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1677677812
transform 1 0 2996 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_652
timestamp 1677677812
transform 1 0 3004 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1677677812
transform 1 0 3012 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_457
timestamp 1677677812
transform 1 0 3028 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_538
timestamp 1677677812
transform 1 0 3028 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_414
timestamp 1677677812
transform 1 0 3076 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_458
timestamp 1677677812
transform 1 0 3092 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1677677812
transform 1 0 3068 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_539
timestamp 1677677812
transform 1 0 3076 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1677677812
transform 1 0 3092 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_415
timestamp 1677677812
transform 1 0 3108 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_653
timestamp 1677677812
transform 1 0 3060 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_654
timestamp 1677677812
transform 1 0 3068 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1677677812
transform 1 0 3084 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1677677812
transform 1 0 3100 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_546
timestamp 1677677812
transform 1 0 3060 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1677677812
transform 1 0 3084 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_657
timestamp 1677677812
transform 1 0 3116 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_541
timestamp 1677677812
transform 1 0 3164 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_658
timestamp 1677677812
transform 1 0 3140 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_524
timestamp 1677677812
transform 1 0 3164 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_485
timestamp 1677677812
transform 1 0 3228 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_547
timestamp 1677677812
transform 1 0 3244 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_387
timestamp 1677677812
transform 1 0 3260 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1677677812
transform 1 0 3260 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_542
timestamp 1677677812
transform 1 0 3260 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_543
timestamp 1677677812
transform 1 0 3308 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_659
timestamp 1677677812
transform 1 0 3284 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1677677812
transform 1 0 3404 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1677677812
transform 1 0 3404 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_548
timestamp 1677677812
transform 1 0 3404 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1677677812
transform 1 0 3420 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1677677812
transform 1 0 3428 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_445
timestamp 1677677812
transform 1 0 3428 0 1 4435
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1677677812
transform 1 0 3436 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_416
timestamp 1677677812
transform 1 0 3476 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1677677812
transform 1 0 3508 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_389
timestamp 1677677812
transform 1 0 3588 0 1 4455
box -3 -3 3 3
use M3_M2  M3_M2_396
timestamp 1677677812
transform 1 0 3500 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_446
timestamp 1677677812
transform 1 0 3492 0 1 4435
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1677677812
transform 1 0 3476 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1677677812
transform 1 0 3484 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1677677812
transform 1 0 3508 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1677677812
transform 1 0 3500 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1677677812
transform 1 0 3516 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1677677812
transform 1 0 3572 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1677677812
transform 1 0 3596 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_417
timestamp 1677677812
transform 1 0 3668 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_549
timestamp 1677677812
transform 1 0 3684 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_505
timestamp 1677677812
transform 1 0 3700 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1677677812
transform 1 0 3724 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_378
timestamp 1677677812
transform 1 0 3756 0 1 4465
box -3 -3 3 3
use M2_M1  M2_M1_550
timestamp 1677677812
transform 1 0 3724 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1677677812
transform 1 0 3740 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1677677812
transform 1 0 3756 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_661
timestamp 1677677812
transform 1 0 3732 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_525
timestamp 1677677812
transform 1 0 3732 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_662
timestamp 1677677812
transform 1 0 3764 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_461
timestamp 1677677812
transform 1 0 3804 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_553
timestamp 1677677812
transform 1 0 3788 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_486
timestamp 1677677812
transform 1 0 3796 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1677677812
transform 1 0 3836 0 1 4465
box -3 -3 3 3
use M2_M1  M2_M1_554
timestamp 1677677812
transform 1 0 3836 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_418
timestamp 1677677812
transform 1 0 3868 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1677677812
transform 1 0 3884 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_555
timestamp 1677677812
transform 1 0 3868 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1677677812
transform 1 0 3884 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1677677812
transform 1 0 3852 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_664
timestamp 1677677812
transform 1 0 3860 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1677677812
transform 1 0 3908 0 1 4425
box -2 -2 2 2
use M3_M2  M3_M2_463
timestamp 1677677812
transform 1 0 3924 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_665
timestamp 1677677812
transform 1 0 3924 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_447
timestamp 1677677812
transform 1 0 3940 0 1 4435
box -2 -2 2 2
use M3_M2  M3_M2_419
timestamp 1677677812
transform 1 0 3948 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_463
timestamp 1677677812
transform 1 0 3948 0 1 4425
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1677677812
transform 1 0 3948 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_549
timestamp 1677677812
transform 1 0 3948 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1677677812
transform 1 0 3964 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_558
timestamp 1677677812
transform 1 0 3964 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_559
timestamp 1677677812
transform 1 0 3996 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_465
timestamp 1677677812
transform 1 0 4020 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_560
timestamp 1677677812
transform 1 0 4012 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_487
timestamp 1677677812
transform 1 0 4020 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_526
timestamp 1677677812
transform 1 0 4012 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_561
timestamp 1677677812
transform 1 0 4028 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_666
timestamp 1677677812
transform 1 0 4028 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_466
timestamp 1677677812
transform 1 0 4092 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_562
timestamp 1677677812
transform 1 0 4092 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_667
timestamp 1677677812
transform 1 0 4140 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_527
timestamp 1677677812
transform 1 0 4116 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_528
timestamp 1677677812
transform 1 0 4140 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_563
timestamp 1677677812
transform 1 0 4172 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1677677812
transform 1 0 4164 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_506
timestamp 1677677812
transform 1 0 4172 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1677677812
transform 1 0 4164 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1677677812
transform 1 0 4196 0 1 4445
box -3 -3 3 3
use M2_M1  M2_M1_564
timestamp 1677677812
transform 1 0 4196 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_420
timestamp 1677677812
transform 1 0 4220 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_565
timestamp 1677677812
transform 1 0 4220 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_669
timestamp 1677677812
transform 1 0 4236 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1677677812
transform 1 0 4252 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_530
timestamp 1677677812
transform 1 0 4252 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_488
timestamp 1677677812
transform 1 0 4276 0 1 4415
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1677677812
transform 1 0 4276 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_670
timestamp 1677677812
transform 1 0 4284 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_671
timestamp 1677677812
transform 1 0 4292 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1677677812
transform 1 0 4308 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_421
timestamp 1677677812
transform 1 0 4380 0 1 4435
box -3 -3 3 3
use M2_M1  M2_M1_567
timestamp 1677677812
transform 1 0 4340 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_568
timestamp 1677677812
transform 1 0 4348 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1677677812
transform 1 0 4364 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_489
timestamp 1677677812
transform 1 0 4372 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_570
timestamp 1677677812
transform 1 0 4380 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_673
timestamp 1677677812
transform 1 0 4356 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1677677812
transform 1 0 4372 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_380
timestamp 1677677812
transform 1 0 4436 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_422
timestamp 1677677812
transform 1 0 4412 0 1 4435
box -3 -3 3 3
use M3_M2  M3_M2_490
timestamp 1677677812
transform 1 0 4412 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_571
timestamp 1677677812
transform 1 0 4420 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_572
timestamp 1677677812
transform 1 0 4436 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_573
timestamp 1677677812
transform 1 0 4444 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1677677812
transform 1 0 4412 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_507
timestamp 1677677812
transform 1 0 4428 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_550
timestamp 1677677812
transform 1 0 4420 0 1 4385
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1677677812
transform 1 0 4452 0 1 4425
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1677677812
transform 1 0 4444 0 1 4405
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1677677812
transform 1 0 4484 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_574
timestamp 1677677812
transform 1 0 4484 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_469
timestamp 1677677812
transform 1 0 4500 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_575
timestamp 1677677812
transform 1 0 4500 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1677677812
transform 1 0 4452 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1677677812
transform 1 0 4460 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1677677812
transform 1 0 4476 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1677677812
transform 1 0 4492 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1677677812
transform 1 0 4460 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_576
timestamp 1677677812
transform 1 0 4524 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_509
timestamp 1677677812
transform 1 0 4524 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_680
timestamp 1677677812
transform 1 0 4532 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_491
timestamp 1677677812
transform 1 0 4540 0 1 4415
box -3 -3 3 3
use M2_M1  M2_M1_681
timestamp 1677677812
transform 1 0 4540 0 1 4405
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1677677812
transform 1 0 4564 0 1 4415
box -2 -2 2 2
use M3_M2  M3_M2_510
timestamp 1677677812
transform 1 0 4564 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_682
timestamp 1677677812
transform 1 0 4572 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_381
timestamp 1677677812
transform 1 0 4588 0 1 4465
box -3 -3 3 3
use M3_M2  M3_M2_470
timestamp 1677677812
transform 1 0 4604 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_578
timestamp 1677677812
transform 1 0 4604 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_579
timestamp 1677677812
transform 1 0 4620 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_683
timestamp 1677677812
transform 1 0 4612 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_511
timestamp 1677677812
transform 1 0 4620 0 1 4405
box -3 -3 3 3
use M2_M1  M2_M1_684
timestamp 1677677812
transform 1 0 4628 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1677677812
transform 1 0 4612 0 1 4395
box -3 -3 3 3
use M2_M1  M2_M1_580
timestamp 1677677812
transform 1 0 4692 0 1 4415
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1677677812
transform 1 0 4668 0 1 4405
box -2 -2 2 2
use M3_M2  M3_M2_534
timestamp 1677677812
transform 1 0 4692 0 1 4395
box -3 -3 3 3
use M3_M2  M3_M2_471
timestamp 1677677812
transform 1 0 4780 0 1 4425
box -3 -3 3 3
use M2_M1  M2_M1_581
timestamp 1677677812
transform 1 0 4780 0 1 4415
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_6
timestamp 1677677812
transform 1 0 48 0 1 4370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_35
timestamp 1677677812
transform 1 0 72 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_40
timestamp 1677677812
transform -1 0 184 0 1 4370
box -9 -3 26 105
use AOI22X1  AOI22X1_22
timestamp 1677677812
transform -1 0 224 0 1 4370
box -8 -3 46 105
use FILL  FILL_412
timestamp 1677677812
transform 1 0 224 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_21
timestamp 1677677812
transform 1 0 232 0 1 4370
box -8 -3 46 105
use FILL  FILL_413
timestamp 1677677812
transform 1 0 272 0 1 4370
box -8 -3 16 105
use FILL  FILL_414
timestamp 1677677812
transform 1 0 280 0 1 4370
box -8 -3 16 105
use FILL  FILL_415
timestamp 1677677812
transform 1 0 288 0 1 4370
box -8 -3 16 105
use FILL  FILL_416
timestamp 1677677812
transform 1 0 296 0 1 4370
box -8 -3 16 105
use FILL  FILL_417
timestamp 1677677812
transform 1 0 304 0 1 4370
box -8 -3 16 105
use FILL  FILL_418
timestamp 1677677812
transform 1 0 312 0 1 4370
box -8 -3 16 105
use FILL  FILL_426
timestamp 1677677812
transform 1 0 320 0 1 4370
box -8 -3 16 105
use FILL  FILL_427
timestamp 1677677812
transform 1 0 328 0 1 4370
box -8 -3 16 105
use FILL  FILL_428
timestamp 1677677812
transform 1 0 336 0 1 4370
box -8 -3 16 105
use FILL  FILL_429
timestamp 1677677812
transform 1 0 344 0 1 4370
box -8 -3 16 105
use FILL  FILL_430
timestamp 1677677812
transform 1 0 352 0 1 4370
box -8 -3 16 105
use FILL  FILL_431
timestamp 1677677812
transform 1 0 360 0 1 4370
box -8 -3 16 105
use FILL  FILL_432
timestamp 1677677812
transform 1 0 368 0 1 4370
box -8 -3 16 105
use FILL  FILL_433
timestamp 1677677812
transform 1 0 376 0 1 4370
box -8 -3 16 105
use FILL  FILL_434
timestamp 1677677812
transform 1 0 384 0 1 4370
box -8 -3 16 105
use FILL  FILL_435
timestamp 1677677812
transform 1 0 392 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_42
timestamp 1677677812
transform -1 0 416 0 1 4370
box -9 -3 26 105
use FILL  FILL_436
timestamp 1677677812
transform 1 0 416 0 1 4370
box -8 -3 16 105
use FILL  FILL_437
timestamp 1677677812
transform 1 0 424 0 1 4370
box -8 -3 16 105
use FILL  FILL_440
timestamp 1677677812
transform 1 0 432 0 1 4370
box -8 -3 16 105
use FILL  FILL_442
timestamp 1677677812
transform 1 0 440 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_24
timestamp 1677677812
transform -1 0 488 0 1 4370
box -8 -3 46 105
use FILL  FILL_443
timestamp 1677677812
transform 1 0 488 0 1 4370
box -8 -3 16 105
use FILL  FILL_444
timestamp 1677677812
transform 1 0 496 0 1 4370
box -8 -3 16 105
use FILL  FILL_445
timestamp 1677677812
transform 1 0 504 0 1 4370
box -8 -3 16 105
use FILL  FILL_446
timestamp 1677677812
transform 1 0 512 0 1 4370
box -8 -3 16 105
use FILL  FILL_447
timestamp 1677677812
transform 1 0 520 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_23
timestamp 1677677812
transform 1 0 528 0 1 4370
box -8 -3 46 105
use FILL  FILL_448
timestamp 1677677812
transform 1 0 568 0 1 4370
box -8 -3 16 105
use FILL  FILL_452
timestamp 1677677812
transform 1 0 576 0 1 4370
box -8 -3 16 105
use FILL  FILL_454
timestamp 1677677812
transform 1 0 584 0 1 4370
box -8 -3 16 105
use FILL  FILL_455
timestamp 1677677812
transform 1 0 592 0 1 4370
box -8 -3 16 105
use FILL  FILL_456
timestamp 1677677812
transform 1 0 600 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_25
timestamp 1677677812
transform 1 0 608 0 1 4370
box -8 -3 46 105
use FILL  FILL_457
timestamp 1677677812
transform 1 0 648 0 1 4370
box -8 -3 16 105
use FILL  FILL_462
timestamp 1677677812
transform 1 0 656 0 1 4370
box -8 -3 16 105
use FILL  FILL_463
timestamp 1677677812
transform 1 0 664 0 1 4370
box -8 -3 16 105
use FILL  FILL_464
timestamp 1677677812
transform 1 0 672 0 1 4370
box -8 -3 16 105
use FILL  FILL_466
timestamp 1677677812
transform 1 0 680 0 1 4370
box -8 -3 16 105
use FILL  FILL_468
timestamp 1677677812
transform 1 0 688 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_39
timestamp 1677677812
transform -1 0 792 0 1 4370
box -8 -3 104 105
use FILL  FILL_469
timestamp 1677677812
transform 1 0 792 0 1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_3
timestamp 1677677812
transform 1 0 800 0 1 4370
box -8 -3 32 105
use FILL  FILL_482
timestamp 1677677812
transform 1 0 824 0 1 4370
box -8 -3 16 105
use FILL  FILL_483
timestamp 1677677812
transform 1 0 832 0 1 4370
box -8 -3 16 105
use FILL  FILL_484
timestamp 1677677812
transform 1 0 840 0 1 4370
box -8 -3 16 105
use FILL  FILL_485
timestamp 1677677812
transform 1 0 848 0 1 4370
box -8 -3 16 105
use FILL  FILL_486
timestamp 1677677812
transform 1 0 856 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_27
timestamp 1677677812
transform 1 0 864 0 1 4370
box -8 -3 46 105
use FILL  FILL_487
timestamp 1677677812
transform 1 0 904 0 1 4370
box -8 -3 16 105
use FILL  FILL_488
timestamp 1677677812
transform 1 0 912 0 1 4370
box -8 -3 16 105
use FILL  FILL_489
timestamp 1677677812
transform 1 0 920 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_46
timestamp 1677677812
transform 1 0 928 0 1 4370
box -9 -3 26 105
use OAI21X1  OAI21X1_10
timestamp 1677677812
transform 1 0 944 0 1 4370
box -8 -3 34 105
use FILL  FILL_494
timestamp 1677677812
transform 1 0 976 0 1 4370
box -8 -3 16 105
use FILL  FILL_495
timestamp 1677677812
transform 1 0 984 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_551
timestamp 1677677812
transform 1 0 1004 0 1 4375
box -3 -3 3 3
use FILL  FILL_496
timestamp 1677677812
transform 1 0 992 0 1 4370
box -8 -3 16 105
use FILL  FILL_497
timestamp 1677677812
transform 1 0 1000 0 1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1677677812
transform 1 0 1008 0 1 4370
box -8 -3 32 105
use NOR2X1  NOR2X1_5
timestamp 1677677812
transform 1 0 1032 0 1 4370
box -8 -3 32 105
use OAI21X1  OAI21X1_11
timestamp 1677677812
transform 1 0 1056 0 1 4370
box -8 -3 34 105
use FILL  FILL_498
timestamp 1677677812
transform 1 0 1088 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_12
timestamp 1677677812
transform -1 0 1128 0 1 4370
box -8 -3 34 105
use FILL  FILL_499
timestamp 1677677812
transform 1 0 1128 0 1 4370
box -8 -3 16 105
use FILL  FILL_510
timestamp 1677677812
transform 1 0 1136 0 1 4370
box -8 -3 16 105
use FILL  FILL_512
timestamp 1677677812
transform 1 0 1144 0 1 4370
box -8 -3 16 105
use FILL  FILL_514
timestamp 1677677812
transform 1 0 1152 0 1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1677677812
transform 1 0 1160 0 1 4370
box -8 -3 32 105
use FILL  FILL_515
timestamp 1677677812
transform 1 0 1184 0 1 4370
box -8 -3 16 105
use FILL  FILL_516
timestamp 1677677812
transform 1 0 1192 0 1 4370
box -8 -3 16 105
use FILL  FILL_517
timestamp 1677677812
transform 1 0 1200 0 1 4370
box -8 -3 16 105
use FILL  FILL_518
timestamp 1677677812
transform 1 0 1208 0 1 4370
box -8 -3 16 105
use FILL  FILL_519
timestamp 1677677812
transform 1 0 1216 0 1 4370
box -8 -3 16 105
use FILL  FILL_520
timestamp 1677677812
transform 1 0 1224 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_552
timestamp 1677677812
transform 1 0 1268 0 1 4375
box -3 -3 3 3
use OAI21X1  OAI21X1_14
timestamp 1677677812
transform -1 0 1264 0 1 4370
box -8 -3 34 105
use OAI21X1  OAI21X1_15
timestamp 1677677812
transform -1 0 1296 0 1 4370
box -8 -3 34 105
use OAI21X1  OAI21X1_16
timestamp 1677677812
transform -1 0 1328 0 1 4370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1677677812
transform 1 0 1328 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_48
timestamp 1677677812
transform 1 0 1424 0 1 4370
box -9 -3 26 105
use FILL  FILL_521
timestamp 1677677812
transform 1 0 1440 0 1 4370
box -8 -3 16 105
use FILL  FILL_522
timestamp 1677677812
transform 1 0 1448 0 1 4370
box -8 -3 16 105
use FILL  FILL_529
timestamp 1677677812
transform 1 0 1456 0 1 4370
box -8 -3 16 105
use FILL  FILL_530
timestamp 1677677812
transform 1 0 1464 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_24
timestamp 1677677812
transform -1 0 1512 0 1 4370
box -8 -3 46 105
use FILL  FILL_531
timestamp 1677677812
transform 1 0 1512 0 1 4370
box -8 -3 16 105
use FILL  FILL_535
timestamp 1677677812
transform 1 0 1520 0 1 4370
box -8 -3 16 105
use FILL  FILL_536
timestamp 1677677812
transform 1 0 1528 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_553
timestamp 1677677812
transform 1 0 1548 0 1 4375
box -3 -3 3 3
use M3_M2  M3_M2_554
timestamp 1677677812
transform 1 0 1620 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_44
timestamp 1677677812
transform 1 0 1536 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_51
timestamp 1677677812
transform 1 0 1632 0 1 4370
box -9 -3 26 105
use FILL  FILL_537
timestamp 1677677812
transform 1 0 1648 0 1 4370
box -8 -3 16 105
use FILL  FILL_541
timestamp 1677677812
transform 1 0 1656 0 1 4370
box -8 -3 16 105
use FILL  FILL_543
timestamp 1677677812
transform 1 0 1664 0 1 4370
box -8 -3 16 105
use FILL  FILL_544
timestamp 1677677812
transform 1 0 1672 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_26
timestamp 1677677812
transform -1 0 1720 0 1 4370
box -8 -3 46 105
use FILL  FILL_545
timestamp 1677677812
transform 1 0 1720 0 1 4370
box -8 -3 16 105
use FILL  FILL_546
timestamp 1677677812
transform 1 0 1728 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_53
timestamp 1677677812
transform 1 0 1736 0 1 4370
box -9 -3 26 105
use FILL  FILL_547
timestamp 1677677812
transform 1 0 1752 0 1 4370
box -8 -3 16 105
use FILL  FILL_548
timestamp 1677677812
transform 1 0 1760 0 1 4370
box -8 -3 16 105
use FILL  FILL_549
timestamp 1677677812
transform 1 0 1768 0 1 4370
box -8 -3 16 105
use FILL  FILL_550
timestamp 1677677812
transform 1 0 1776 0 1 4370
box -8 -3 16 105
use FILL  FILL_551
timestamp 1677677812
transform 1 0 1784 0 1 4370
box -8 -3 16 105
use FILL  FILL_554
timestamp 1677677812
transform 1 0 1792 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_30
timestamp 1677677812
transform 1 0 1800 0 1 4370
box -8 -3 46 105
use FILL  FILL_556
timestamp 1677677812
transform 1 0 1840 0 1 4370
box -8 -3 16 105
use FILL  FILL_557
timestamp 1677677812
transform 1 0 1848 0 1 4370
box -8 -3 16 105
use FILL  FILL_558
timestamp 1677677812
transform 1 0 1856 0 1 4370
box -8 -3 16 105
use FILL  FILL_559
timestamp 1677677812
transform 1 0 1864 0 1 4370
box -8 -3 16 105
use FILL  FILL_564
timestamp 1677677812
transform 1 0 1872 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_555
timestamp 1677677812
transform 1 0 1924 0 1 4375
box -3 -3 3 3
use OAI22X1  OAI22X1_27
timestamp 1677677812
transform 1 0 1880 0 1 4370
box -8 -3 46 105
use FILL  FILL_566
timestamp 1677677812
transform 1 0 1920 0 1 4370
box -8 -3 16 105
use FILL  FILL_567
timestamp 1677677812
transform 1 0 1928 0 1 4370
box -8 -3 16 105
use FILL  FILL_568
timestamp 1677677812
transform 1 0 1936 0 1 4370
box -8 -3 16 105
use FILL  FILL_569
timestamp 1677677812
transform 1 0 1944 0 1 4370
box -8 -3 16 105
use FILL  FILL_574
timestamp 1677677812
transform 1 0 1952 0 1 4370
box -8 -3 16 105
use FILL  FILL_576
timestamp 1677677812
transform 1 0 1960 0 1 4370
box -8 -3 16 105
use FILL  FILL_578
timestamp 1677677812
transform 1 0 1968 0 1 4370
box -8 -3 16 105
use FILL  FILL_580
timestamp 1677677812
transform 1 0 1976 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_32
timestamp 1677677812
transform -1 0 2024 0 1 4370
box -8 -3 46 105
use FILL  FILL_581
timestamp 1677677812
transform 1 0 2024 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1677677812
transform -1 0 2128 0 1 4370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1677677812
transform 1 0 2128 0 1 4370
box -8 -3 104 105
use OAI22X1  OAI22X1_29
timestamp 1677677812
transform 1 0 2224 0 1 4370
box -8 -3 46 105
use FILL  FILL_582
timestamp 1677677812
transform 1 0 2264 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_55
timestamp 1677677812
transform 1 0 2272 0 1 4370
box -9 -3 26 105
use FILL  FILL_583
timestamp 1677677812
transform 1 0 2288 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1677677812
transform 1 0 2296 0 1 4370
box -8 -3 104 105
use INVX2  INVX2_60
timestamp 1677677812
transform 1 0 2392 0 1 4370
box -9 -3 26 105
use FILL  FILL_599
timestamp 1677677812
transform 1 0 2408 0 1 4370
box -8 -3 16 105
use FILL  FILL_600
timestamp 1677677812
transform 1 0 2416 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_51
timestamp 1677677812
transform -1 0 2520 0 1 4370
box -8 -3 104 105
use FILL  FILL_601
timestamp 1677677812
transform 1 0 2520 0 1 4370
box -8 -3 16 105
use FILL  FILL_616
timestamp 1677677812
transform 1 0 2528 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_61
timestamp 1677677812
transform 1 0 2536 0 1 4370
box -9 -3 26 105
use FILL  FILL_617
timestamp 1677677812
transform 1 0 2552 0 1 4370
box -8 -3 16 105
use FILL  FILL_618
timestamp 1677677812
transform 1 0 2560 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_52
timestamp 1677677812
transform 1 0 2568 0 1 4370
box -8 -3 104 105
use FILL  FILL_619
timestamp 1677677812
transform 1 0 2664 0 1 4370
box -8 -3 16 105
use FILL  FILL_620
timestamp 1677677812
transform 1 0 2672 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_63
timestamp 1677677812
transform 1 0 2680 0 1 4370
box -9 -3 26 105
use FILL  FILL_628
timestamp 1677677812
transform 1 0 2696 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_556
timestamp 1677677812
transform 1 0 2796 0 1 4375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_53
timestamp 1677677812
transform 1 0 2704 0 1 4370
box -8 -3 104 105
use FILL  FILL_629
timestamp 1677677812
transform 1 0 2800 0 1 4370
box -8 -3 16 105
use FILL  FILL_634
timestamp 1677677812
transform 1 0 2808 0 1 4370
box -8 -3 16 105
use FILL  FILL_636
timestamp 1677677812
transform 1 0 2816 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_18
timestamp 1677677812
transform 1 0 2824 0 1 4370
box -8 -3 34 105
use M3_M2  M3_M2_557
timestamp 1677677812
transform 1 0 2868 0 1 4375
box -3 -3 3 3
use FILL  FILL_637
timestamp 1677677812
transform 1 0 2856 0 1 4370
box -8 -3 16 105
use FILL  FILL_638
timestamp 1677677812
transform 1 0 2864 0 1 4370
box -8 -3 16 105
use FILL  FILL_639
timestamp 1677677812
transform 1 0 2872 0 1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_7
timestamp 1677677812
transform 1 0 2880 0 1 4370
box -8 -3 32 105
use OAI21X1  OAI21X1_19
timestamp 1677677812
transform 1 0 2904 0 1 4370
box -8 -3 34 105
use FILL  FILL_640
timestamp 1677677812
transform 1 0 2936 0 1 4370
box -8 -3 16 105
use FILL  FILL_647
timestamp 1677677812
transform 1 0 2944 0 1 4370
box -8 -3 16 105
use FILL  FILL_648
timestamp 1677677812
transform 1 0 2952 0 1 4370
box -8 -3 16 105
use FILL  FILL_649
timestamp 1677677812
transform 1 0 2960 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_21
timestamp 1677677812
transform -1 0 3000 0 1 4370
box -8 -3 34 105
use FILL  FILL_650
timestamp 1677677812
transform 1 0 3000 0 1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_22
timestamp 1677677812
transform -1 0 3040 0 1 4370
box -8 -3 34 105
use FILL  FILL_656
timestamp 1677677812
transform 1 0 3040 0 1 4370
box -8 -3 16 105
use FILL  FILL_658
timestamp 1677677812
transform 1 0 3048 0 1 4370
box -8 -3 16 105
use FILL  FILL_660
timestamp 1677677812
transform 1 0 3056 0 1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_31
timestamp 1677677812
transform 1 0 3064 0 1 4370
box -8 -3 46 105
use FILL  FILL_662
timestamp 1677677812
transform 1 0 3104 0 1 4370
box -8 -3 16 105
use FILL  FILL_663
timestamp 1677677812
transform 1 0 3112 0 1 4370
box -8 -3 16 105
use FILL  FILL_664
timestamp 1677677812
transform 1 0 3120 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1677677812
transform 1 0 3128 0 1 4370
box -8 -3 104 105
use FILL  FILL_665
timestamp 1677677812
transform 1 0 3224 0 1 4370
box -8 -3 16 105
use FILL  FILL_666
timestamp 1677677812
transform 1 0 3232 0 1 4370
box -8 -3 16 105
use FILL  FILL_667
timestamp 1677677812
transform 1 0 3240 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_64
timestamp 1677677812
transform 1 0 3248 0 1 4370
box -9 -3 26 105
use FILL  FILL_668
timestamp 1677677812
transform 1 0 3264 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_57
timestamp 1677677812
transform 1 0 3272 0 1 4370
box -8 -3 104 105
use FILL  FILL_676
timestamp 1677677812
transform 1 0 3368 0 1 4370
box -8 -3 16 105
use FILL  FILL_677
timestamp 1677677812
transform 1 0 3376 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_66
timestamp 1677677812
transform 1 0 3384 0 1 4370
box -9 -3 26 105
use FILL  FILL_678
timestamp 1677677812
transform 1 0 3400 0 1 4370
box -8 -3 16 105
use FILL  FILL_684
timestamp 1677677812
transform 1 0 3408 0 1 4370
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1677677812
transform -1 0 3448 0 1 4370
box -8 -3 40 105
use FILL  FILL_685
timestamp 1677677812
transform 1 0 3448 0 1 4370
box -8 -3 16 105
use FILL  FILL_686
timestamp 1677677812
transform 1 0 3456 0 1 4370
box -8 -3 16 105
use FILL  FILL_687
timestamp 1677677812
transform 1 0 3464 0 1 4370
box -8 -3 16 105
use FILL  FILL_688
timestamp 1677677812
transform 1 0 3472 0 1 4370
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1677677812
transform -1 0 3512 0 1 4370
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_59
timestamp 1677677812
transform -1 0 3608 0 1 4370
box -8 -3 104 105
use FILL  FILL_689
timestamp 1677677812
transform 1 0 3608 0 1 4370
box -8 -3 16 105
use FILL  FILL_702
timestamp 1677677812
transform 1 0 3616 0 1 4370
box -8 -3 16 105
use FILL  FILL_704
timestamp 1677677812
transform 1 0 3624 0 1 4370
box -8 -3 16 105
use FILL  FILL_706
timestamp 1677677812
transform 1 0 3632 0 1 4370
box -8 -3 16 105
use FILL  FILL_708
timestamp 1677677812
transform 1 0 3640 0 1 4370
box -8 -3 16 105
use FILL  FILL_709
timestamp 1677677812
transform 1 0 3648 0 1 4370
box -8 -3 16 105
use FILL  FILL_710
timestamp 1677677812
transform 1 0 3656 0 1 4370
box -8 -3 16 105
use FILL  FILL_711
timestamp 1677677812
transform 1 0 3664 0 1 4370
box -8 -3 16 105
use FILL  FILL_712
timestamp 1677677812
transform 1 0 3672 0 1 4370
box -8 -3 16 105
use FILL  FILL_713
timestamp 1677677812
transform 1 0 3680 0 1 4370
box -8 -3 16 105
use FILL  FILL_715
timestamp 1677677812
transform 1 0 3688 0 1 4370
box -8 -3 16 105
use FILL  FILL_717
timestamp 1677677812
transform 1 0 3696 0 1 4370
box -8 -3 16 105
use FILL  FILL_719
timestamp 1677677812
transform 1 0 3704 0 1 4370
box -8 -3 16 105
use FILL  FILL_720
timestamp 1677677812
transform 1 0 3712 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_38
timestamp 1677677812
transform 1 0 3720 0 1 4370
box -8 -3 46 105
use FILL  FILL_721
timestamp 1677677812
transform 1 0 3760 0 1 4370
box -8 -3 16 105
use FILL  FILL_722
timestamp 1677677812
transform 1 0 3768 0 1 4370
box -8 -3 16 105
use FILL  FILL_723
timestamp 1677677812
transform 1 0 3776 0 1 4370
box -8 -3 16 105
use FILL  FILL_724
timestamp 1677677812
transform 1 0 3784 0 1 4370
box -8 -3 16 105
use FILL  FILL_725
timestamp 1677677812
transform 1 0 3792 0 1 4370
box -8 -3 16 105
use FILL  FILL_726
timestamp 1677677812
transform 1 0 3800 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_68
timestamp 1677677812
transform -1 0 3824 0 1 4370
box -9 -3 26 105
use FILL  FILL_727
timestamp 1677677812
transform 1 0 3824 0 1 4370
box -8 -3 16 105
use FILL  FILL_728
timestamp 1677677812
transform 1 0 3832 0 1 4370
box -8 -3 16 105
use FILL  FILL_732
timestamp 1677677812
transform 1 0 3840 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_39
timestamp 1677677812
transform -1 0 3888 0 1 4370
box -8 -3 46 105
use FILL  FILL_733
timestamp 1677677812
transform 1 0 3888 0 1 4370
box -8 -3 16 105
use FILL  FILL_734
timestamp 1677677812
transform 1 0 3896 0 1 4370
box -8 -3 16 105
use FILL  FILL_735
timestamp 1677677812
transform 1 0 3904 0 1 4370
box -8 -3 16 105
use FILL  FILL_740
timestamp 1677677812
transform 1 0 3912 0 1 4370
box -8 -3 16 105
use FILL  FILL_742
timestamp 1677677812
transform 1 0 3920 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_558
timestamp 1677677812
transform 1 0 3940 0 1 4375
box -3 -3 3 3
use NAND3X1  NAND3X1_3
timestamp 1677677812
transform -1 0 3960 0 1 4370
box -8 -3 40 105
use FILL  FILL_743
timestamp 1677677812
transform 1 0 3960 0 1 4370
box -8 -3 16 105
use FILL  FILL_748
timestamp 1677677812
transform 1 0 3968 0 1 4370
box -8 -3 16 105
use FILL  FILL_750
timestamp 1677677812
transform 1 0 3976 0 1 4370
box -8 -3 16 105
use FILL  FILL_751
timestamp 1677677812
transform 1 0 3984 0 1 4370
box -8 -3 16 105
use FILL  FILL_752
timestamp 1677677812
transform 1 0 3992 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_71
timestamp 1677677812
transform -1 0 4016 0 1 4370
box -9 -3 26 105
use FILL  FILL_753
timestamp 1677677812
transform 1 0 4016 0 1 4370
box -8 -3 16 105
use FILL  FILL_754
timestamp 1677677812
transform 1 0 4024 0 1 4370
box -8 -3 16 105
use FILL  FILL_755
timestamp 1677677812
transform 1 0 4032 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_72
timestamp 1677677812
transform -1 0 4056 0 1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_62
timestamp 1677677812
transform -1 0 4152 0 1 4370
box -8 -3 104 105
use FILL  FILL_756
timestamp 1677677812
transform 1 0 4152 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_559
timestamp 1677677812
transform 1 0 4172 0 1 4375
box -3 -3 3 3
use FILL  FILL_757
timestamp 1677677812
transform 1 0 4160 0 1 4370
box -8 -3 16 105
use FILL  FILL_758
timestamp 1677677812
transform 1 0 4168 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_40
timestamp 1677677812
transform -1 0 4216 0 1 4370
box -8 -3 46 105
use FILL  FILL_759
timestamp 1677677812
transform 1 0 4216 0 1 4370
box -8 -3 16 105
use FILL  FILL_760
timestamp 1677677812
transform 1 0 4224 0 1 4370
box -8 -3 16 105
use FILL  FILL_761
timestamp 1677677812
transform 1 0 4232 0 1 4370
box -8 -3 16 105
use FILL  FILL_762
timestamp 1677677812
transform 1 0 4240 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_73
timestamp 1677677812
transform -1 0 4264 0 1 4370
box -9 -3 26 105
use FILL  FILL_763
timestamp 1677677812
transform 1 0 4264 0 1 4370
box -8 -3 16 105
use FILL  FILL_764
timestamp 1677677812
transform 1 0 4272 0 1 4370
box -8 -3 16 105
use FILL  FILL_765
timestamp 1677677812
transform 1 0 4280 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_74
timestamp 1677677812
transform 1 0 4288 0 1 4370
box -9 -3 26 105
use FILL  FILL_766
timestamp 1677677812
transform 1 0 4304 0 1 4370
box -8 -3 16 105
use FILL  FILL_767
timestamp 1677677812
transform 1 0 4312 0 1 4370
box -8 -3 16 105
use FILL  FILL_768
timestamp 1677677812
transform 1 0 4320 0 1 4370
box -8 -3 16 105
use FILL  FILL_777
timestamp 1677677812
transform 1 0 4328 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_560
timestamp 1677677812
transform 1 0 4372 0 1 4375
box -3 -3 3 3
use OAI22X1  OAI22X1_37
timestamp 1677677812
transform 1 0 4336 0 1 4370
box -8 -3 46 105
use FILL  FILL_778
timestamp 1677677812
transform 1 0 4376 0 1 4370
box -8 -3 16 105
use FILL  FILL_779
timestamp 1677677812
transform 1 0 4384 0 1 4370
box -8 -3 16 105
use FILL  FILL_780
timestamp 1677677812
transform 1 0 4392 0 1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_41
timestamp 1677677812
transform 1 0 4400 0 1 4370
box -8 -3 46 105
use FILL  FILL_781
timestamp 1677677812
transform 1 0 4440 0 1 4370
box -8 -3 16 105
use FILL  FILL_782
timestamp 1677677812
transform 1 0 4448 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_561
timestamp 1677677812
transform 1 0 4492 0 1 4375
box -3 -3 3 3
use OAI22X1  OAI22X1_38
timestamp 1677677812
transform 1 0 4456 0 1 4370
box -8 -3 46 105
use FILL  FILL_783
timestamp 1677677812
transform 1 0 4496 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_76
timestamp 1677677812
transform -1 0 4520 0 1 4370
box -9 -3 26 105
use FILL  FILL_784
timestamp 1677677812
transform 1 0 4520 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_562
timestamp 1677677812
transform 1 0 4540 0 1 4375
box -3 -3 3 3
use FILL  FILL_785
timestamp 1677677812
transform 1 0 4528 0 1 4370
box -8 -3 16 105
use FILL  FILL_786
timestamp 1677677812
transform 1 0 4536 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_563
timestamp 1677677812
transform 1 0 4572 0 1 4375
box -3 -3 3 3
use INVX2  INVX2_77
timestamp 1677677812
transform 1 0 4544 0 1 4370
box -9 -3 26 105
use FILL  FILL_790
timestamp 1677677812
transform 1 0 4560 0 1 4370
box -8 -3 16 105
use FILL  FILL_791
timestamp 1677677812
transform 1 0 4568 0 1 4370
box -8 -3 16 105
use FILL  FILL_792
timestamp 1677677812
transform 1 0 4576 0 1 4370
box -8 -3 16 105
use FILL  FILL_793
timestamp 1677677812
transform 1 0 4584 0 1 4370
box -8 -3 16 105
use M3_M2  M3_M2_564
timestamp 1677677812
transform 1 0 4604 0 1 4375
box -3 -3 3 3
use OAI22X1  OAI22X1_39
timestamp 1677677812
transform -1 0 4632 0 1 4370
box -8 -3 46 105
use FILL  FILL_794
timestamp 1677677812
transform 1 0 4632 0 1 4370
box -8 -3 16 105
use FILL  FILL_795
timestamp 1677677812
transform 1 0 4640 0 1 4370
box -8 -3 16 105
use FILL  FILL_802
timestamp 1677677812
transform 1 0 4648 0 1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_67
timestamp 1677677812
transform 1 0 4656 0 1 4370
box -8 -3 104 105
use FILL  FILL_804
timestamp 1677677812
transform 1 0 4752 0 1 4370
box -8 -3 16 105
use FILL  FILL_805
timestamp 1677677812
transform 1 0 4760 0 1 4370
box -8 -3 16 105
use INVX2  INVX2_79
timestamp 1677677812
transform 1 0 4768 0 1 4370
box -9 -3 26 105
use FILL  FILL_806
timestamp 1677677812
transform 1 0 4784 0 1 4370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_7
timestamp 1677677812
transform 1 0 4819 0 1 4370
box -10 -3 10 3
use M2_M1  M2_M1_695
timestamp 1677677812
transform 1 0 92 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1677677812
transform 1 0 140 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1677677812
transform 1 0 172 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_796
timestamp 1677677812
transform 1 0 180 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1677677812
transform 1 0 188 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_678
timestamp 1677677812
transform 1 0 140 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1677677812
transform 1 0 180 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_699
timestamp 1677677812
transform 1 0 172 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_565
timestamp 1677677812
transform 1 0 236 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_696
timestamp 1677677812
transform 1 0 204 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_697
timestamp 1677677812
transform 1 0 212 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_698
timestamp 1677677812
transform 1 0 228 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_699
timestamp 1677677812
transform 1 0 236 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_798
timestamp 1677677812
transform 1 0 204 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1677677812
transform 1 0 220 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_700
timestamp 1677677812
transform 1 0 212 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_700
timestamp 1677677812
transform 1 0 252 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_701
timestamp 1677677812
transform 1 0 252 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1677677812
transform 1 0 268 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_581
timestamp 1677677812
transform 1 0 292 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_701
timestamp 1677677812
transform 1 0 292 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_626
timestamp 1677677812
transform 1 0 300 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_702
timestamp 1677677812
transform 1 0 308 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_800
timestamp 1677677812
transform 1 0 284 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1677677812
transform 1 0 300 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1677677812
transform 1 0 412 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1677677812
transform 1 0 332 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_803
timestamp 1677677812
transform 1 0 388 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_649
timestamp 1677677812
transform 1 0 412 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_704
timestamp 1677677812
transform 1 0 460 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_627
timestamp 1677677812
transform 1 0 540 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_650
timestamp 1677677812
transform 1 0 460 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1677677812
transform 1 0 484 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_804
timestamp 1677677812
transform 1 0 508 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1677677812
transform 1 0 540 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1677677812
transform 1 0 548 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_680
timestamp 1677677812
transform 1 0 508 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1677677812
transform 1 0 548 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_628
timestamp 1677677812
transform 1 0 564 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_807
timestamp 1677677812
transform 1 0 580 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1677677812
transform 1 0 588 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_682
timestamp 1677677812
transform 1 0 588 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_702
timestamp 1677677812
transform 1 0 580 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_706
timestamp 1677677812
transform 1 0 604 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_629
timestamp 1677677812
transform 1 0 612 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_707
timestamp 1677677812
transform 1 0 620 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1677677812
transform 1 0 628 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1677677812
transform 1 0 612 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_652
timestamp 1677677812
transform 1 0 620 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_683
timestamp 1677677812
transform 1 0 612 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1677677812
transform 1 0 636 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_709
timestamp 1677677812
transform 1 0 660 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1677677812
transform 1 0 676 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_653
timestamp 1677677812
transform 1 0 676 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_809
timestamp 1677677812
transform 1 0 756 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1677677812
transform 1 0 788 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_596
timestamp 1677677812
transform 1 0 916 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_711
timestamp 1677677812
transform 1 0 836 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1677677812
transform 1 0 836 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1677677812
transform 1 0 860 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_811
timestamp 1677677812
transform 1 0 884 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_656
timestamp 1677677812
transform 1 0 900 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_812
timestamp 1677677812
transform 1 0 916 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1677677812
transform 1 0 924 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_684
timestamp 1677677812
transform 1 0 884 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_685
timestamp 1677677812
transform 1 0 924 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_582
timestamp 1677677812
transform 1 0 980 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_597
timestamp 1677677812
transform 1 0 996 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_712
timestamp 1677677812
transform 1 0 972 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1677677812
transform 1 0 980 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1677677812
transform 1 0 996 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1677677812
transform 1 0 972 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_657
timestamp 1677677812
transform 1 0 980 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_815
timestamp 1677677812
transform 1 0 988 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1677677812
transform 1 0 1004 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_658
timestamp 1677677812
transform 1 0 1028 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_566
timestamp 1677677812
transform 1 0 1092 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_598
timestamp 1677677812
transform 1 0 1084 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_715
timestamp 1677677812
transform 1 0 1076 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1677677812
transform 1 0 1060 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_659
timestamp 1677677812
transform 1 0 1076 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_716
timestamp 1677677812
transform 1 0 1092 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_717
timestamp 1677677812
transform 1 0 1100 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1677677812
transform 1 0 1116 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1677677812
transform 1 0 1124 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_818
timestamp 1677677812
transform 1 0 1108 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_911
timestamp 1677677812
transform 1 0 1084 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_686
timestamp 1677677812
transform 1 0 1100 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1677677812
transform 1 0 1116 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_819
timestamp 1677677812
transform 1 0 1140 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_705
timestamp 1677677812
transform 1 0 1132 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1677677812
transform 1 0 1236 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_584
timestamp 1677677812
transform 1 0 1276 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_599
timestamp 1677677812
transform 1 0 1268 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1677677812
transform 1 0 1164 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_631
timestamp 1677677812
transform 1 0 1204 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_720
timestamp 1677677812
transform 1 0 1252 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1677677812
transform 1 0 1268 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_820
timestamp 1677677812
transform 1 0 1156 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_821
timestamp 1677677812
transform 1 0 1164 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_822
timestamp 1677677812
transform 1 0 1172 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1677677812
transform 1 0 1204 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_706
timestamp 1677677812
transform 1 0 1172 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_824
timestamp 1677677812
transform 1 0 1292 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_912
timestamp 1677677812
transform 1 0 1276 0 1 4315
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1677677812
transform 1 0 1316 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_660
timestamp 1677677812
transform 1 0 1316 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_687
timestamp 1677677812
transform 1 0 1308 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_600
timestamp 1677677812
transform 1 0 1380 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_723
timestamp 1677677812
transform 1 0 1332 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1677677812
transform 1 0 1380 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_707
timestamp 1677677812
transform 1 0 1332 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_661
timestamp 1677677812
transform 1 0 1436 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_826
timestamp 1677677812
transform 1 0 1444 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_708
timestamp 1677677812
transform 1 0 1428 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_601
timestamp 1677677812
transform 1 0 1484 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_724
timestamp 1677677812
transform 1 0 1468 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_725
timestamp 1677677812
transform 1 0 1484 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_662
timestamp 1677677812
transform 1 0 1468 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_827
timestamp 1677677812
transform 1 0 1476 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1677677812
transform 1 0 1508 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_585
timestamp 1677677812
transform 1 0 1524 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_727
timestamp 1677677812
transform 1 0 1524 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_828
timestamp 1677677812
transform 1 0 1516 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_728
timestamp 1677677812
transform 1 0 1620 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_829
timestamp 1677677812
transform 1 0 1532 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1677677812
transform 1 0 1540 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1677677812
transform 1 0 1580 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_709
timestamp 1677677812
transform 1 0 1532 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_710
timestamp 1677677812
transform 1 0 1580 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_602
timestamp 1677677812
transform 1 0 1756 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_729
timestamp 1677677812
transform 1 0 1676 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_632
timestamp 1677677812
transform 1 0 1724 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1677677812
transform 1 0 1764 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_832
timestamp 1677677812
transform 1 0 1724 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_833
timestamp 1677677812
transform 1 0 1756 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_834
timestamp 1677677812
transform 1 0 1764 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_729
timestamp 1677677812
transform 1 0 1676 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_730
timestamp 1677677812
transform 1 0 1732 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1677677812
transform 1 0 1780 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_835
timestamp 1677677812
transform 1 0 1780 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1677677812
transform 1 0 1812 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_711
timestamp 1677677812
transform 1 0 1812 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_603
timestamp 1677677812
transform 1 0 1852 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_730
timestamp 1677677812
transform 1 0 1828 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1677677812
transform 1 0 1836 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1677677812
transform 1 0 1852 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1677677812
transform 1 0 1844 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_837
timestamp 1677677812
transform 1 0 1860 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_838
timestamp 1677677812
transform 1 0 1876 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1677677812
transform 1 0 1892 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_587
timestamp 1677677812
transform 1 0 1908 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_733
timestamp 1677677812
transform 1 0 1924 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_840
timestamp 1677677812
transform 1 0 1908 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1677677812
transform 1 0 1932 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_712
timestamp 1677677812
transform 1 0 1948 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_723
timestamp 1677677812
transform 1 0 1948 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_604
timestamp 1677677812
transform 1 0 1972 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_734
timestamp 1677677812
transform 1 0 1972 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1677677812
transform 1 0 1980 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_567
timestamp 1677677812
transform 1 0 1996 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_736
timestamp 1677677812
transform 1 0 1996 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_842
timestamp 1677677812
transform 1 0 1996 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_713
timestamp 1677677812
transform 1 0 1996 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1677677812
transform 1 0 2012 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_605
timestamp 1677677812
transform 1 0 2020 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_737
timestamp 1677677812
transform 1 0 2012 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1677677812
transform 1 0 2004 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_569
timestamp 1677677812
transform 1 0 2036 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_844
timestamp 1677677812
transform 1 0 2028 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_606
timestamp 1677677812
transform 1 0 2052 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1677677812
transform 1 0 2132 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_738
timestamp 1677677812
transform 1 0 2132 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1677677812
transform 1 0 2044 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_846
timestamp 1677677812
transform 1 0 2052 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_847
timestamp 1677677812
transform 1 0 2084 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_714
timestamp 1677677812
transform 1 0 2084 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_848
timestamp 1677677812
transform 1 0 2164 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_570
timestamp 1677677812
transform 1 0 2180 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_691
timestamp 1677677812
transform 1 0 2220 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_739
timestamp 1677677812
transform 1 0 2220 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1677677812
transform 1 0 2212 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_663
timestamp 1677677812
transform 1 0 2220 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_740
timestamp 1677677812
transform 1 0 2228 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_571
timestamp 1677677812
transform 1 0 2260 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_741
timestamp 1677677812
transform 1 0 2260 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_664
timestamp 1677677812
transform 1 0 2244 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_850
timestamp 1677677812
transform 1 0 2252 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_851
timestamp 1677677812
transform 1 0 2268 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_731
timestamp 1677677812
transform 1 0 2268 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_634
timestamp 1677677812
transform 1 0 2284 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_608
timestamp 1677677812
transform 1 0 2308 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_852
timestamp 1677677812
transform 1 0 2300 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_715
timestamp 1677677812
transform 1 0 2300 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_635
timestamp 1677677812
transform 1 0 2340 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_853
timestamp 1677677812
transform 1 0 2324 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_665
timestamp 1677677812
transform 1 0 2332 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_854
timestamp 1677677812
transform 1 0 2340 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_724
timestamp 1677677812
transform 1 0 2332 0 1 4295
box -3 -3 3 3
use M2_M1  M2_M1_855
timestamp 1677677812
transform 1 0 2356 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_716
timestamp 1677677812
transform 1 0 2356 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1677677812
transform 1 0 2348 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_572
timestamp 1677677812
transform 1 0 2388 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_742
timestamp 1677677812
transform 1 0 2380 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_743
timestamp 1677677812
transform 1 0 2388 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1677677812
transform 1 0 2404 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_573
timestamp 1677677812
transform 1 0 2436 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_609
timestamp 1677677812
transform 1 0 2428 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_744
timestamp 1677677812
transform 1 0 2428 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_745
timestamp 1677677812
transform 1 0 2436 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1677677812
transform 1 0 2436 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_610
timestamp 1677677812
transform 1 0 2492 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_746
timestamp 1677677812
transform 1 0 2476 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_747
timestamp 1677677812
transform 1 0 2492 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1677677812
transform 1 0 2468 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_859
timestamp 1677677812
transform 1 0 2484 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_717
timestamp 1677677812
transform 1 0 2476 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_636
timestamp 1677677812
transform 1 0 2500 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_860
timestamp 1677677812
transform 1 0 2500 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1677677812
transform 1 0 2532 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_666
timestamp 1677677812
transform 1 0 2532 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_637
timestamp 1677677812
transform 1 0 2564 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_861
timestamp 1677677812
transform 1 0 2548 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1677677812
transform 1 0 2564 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1677677812
transform 1 0 2572 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_732
timestamp 1677677812
transform 1 0 2572 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_611
timestamp 1677677812
transform 1 0 2604 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_749
timestamp 1677677812
transform 1 0 2604 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_750
timestamp 1677677812
transform 1 0 2612 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_751
timestamp 1677677812
transform 1 0 2628 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_752
timestamp 1677677812
transform 1 0 2636 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_667
timestamp 1677677812
transform 1 0 2612 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_864
timestamp 1677677812
transform 1 0 2620 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_668
timestamp 1677677812
transform 1 0 2628 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_638
timestamp 1677677812
transform 1 0 2644 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_865
timestamp 1677677812
transform 1 0 2644 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_612
timestamp 1677677812
transform 1 0 2660 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1677677812
transform 1 0 2676 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1677677812
transform 1 0 2692 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_866
timestamp 1677677812
transform 1 0 2692 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1677677812
transform 1 0 2708 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_641
timestamp 1677677812
transform 1 0 2732 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_867
timestamp 1677677812
transform 1 0 2732 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_669
timestamp 1677677812
transform 1 0 2780 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_692
timestamp 1677677812
transform 1 0 2796 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_868
timestamp 1677677812
transform 1 0 2788 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_733
timestamp 1677677812
transform 1 0 2708 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_734
timestamp 1677677812
transform 1 0 2756 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1677677812
transform 1 0 2828 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_693
timestamp 1677677812
transform 1 0 2844 0 1 4345
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1677677812
transform 1 0 2860 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_755
timestamp 1677677812
transform 1 0 2868 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1677677812
transform 1 0 2876 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_869
timestamp 1677677812
transform 1 0 2852 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_726
timestamp 1677677812
transform 1 0 2844 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1677677812
transform 1 0 2876 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_613
timestamp 1677677812
transform 1 0 2892 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_870
timestamp 1677677812
transform 1 0 2892 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_588
timestamp 1677677812
transform 1 0 2932 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_614
timestamp 1677677812
transform 1 0 2924 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_757
timestamp 1677677812
transform 1 0 2924 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1677677812
transform 1 0 2908 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1677677812
transform 1 0 2932 0 1 4345
box -2 -2 2 2
use M3_M2  M3_M2_671
timestamp 1677677812
transform 1 0 2940 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_914
timestamp 1677677812
transform 1 0 2940 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_718
timestamp 1677677812
transform 1 0 2932 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_758
timestamp 1677677812
transform 1 0 2956 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1677677812
transform 1 0 2972 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1677677812
transform 1 0 2964 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_727
timestamp 1677677812
transform 1 0 2956 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_672
timestamp 1677677812
transform 1 0 2972 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_873
timestamp 1677677812
transform 1 0 3028 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1677677812
transform 1 0 3012 0 1 4315
box -2 -2 2 2
use M3_M2  M3_M2_642
timestamp 1677677812
transform 1 0 3068 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_760
timestamp 1677677812
transform 1 0 3076 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_874
timestamp 1677677812
transform 1 0 3068 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_689
timestamp 1677677812
transform 1 0 3076 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1677677812
transform 1 0 3140 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_615
timestamp 1677677812
transform 1 0 3092 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1677677812
transform 1 0 3140 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_761
timestamp 1677677812
transform 1 0 3092 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_673
timestamp 1677677812
transform 1 0 3092 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_875
timestamp 1677677812
transform 1 0 3132 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_690
timestamp 1677677812
transform 1 0 3124 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_876
timestamp 1677677812
transform 1 0 3188 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1677677812
transform 1 0 3196 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_691
timestamp 1677677812
transform 1 0 3188 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_574
timestamp 1677677812
transform 1 0 3236 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_762
timestamp 1677677812
transform 1 0 3220 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_763
timestamp 1677677812
transform 1 0 3236 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1677677812
transform 1 0 3252 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1677677812
transform 1 0 3212 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_879
timestamp 1677677812
transform 1 0 3244 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_692
timestamp 1677677812
transform 1 0 3244 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_590
timestamp 1677677812
transform 1 0 3284 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_575
timestamp 1677677812
transform 1 0 3308 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1677677812
transform 1 0 3308 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_765
timestamp 1677677812
transform 1 0 3308 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1677677812
transform 1 0 3332 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1677677812
transform 1 0 3388 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_693
timestamp 1677677812
transform 1 0 3332 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_766
timestamp 1677677812
transform 1 0 3420 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1677677812
transform 1 0 3460 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1677677812
transform 1 0 3500 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_767
timestamp 1677677812
transform 1 0 3516 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_617
timestamp 1677677812
transform 1 0 3572 0 1 4345
box -3 -3 3 3
use M3_M2  M3_M2_618
timestamp 1677677812
transform 1 0 3612 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_768
timestamp 1677677812
transform 1 0 3604 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1677677812
transform 1 0 3620 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_885
timestamp 1677677812
transform 1 0 3628 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_694
timestamp 1677677812
transform 1 0 3628 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_592
timestamp 1677677812
transform 1 0 3644 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_769
timestamp 1677677812
transform 1 0 3644 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_770
timestamp 1677677812
transform 1 0 3660 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_771
timestamp 1677677812
transform 1 0 3676 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_886
timestamp 1677677812
transform 1 0 3668 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_674
timestamp 1677677812
transform 1 0 3676 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_735
timestamp 1677677812
transform 1 0 3652 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1677677812
transform 1 0 3788 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_619
timestamp 1677677812
transform 1 0 3764 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1677677812
transform 1 0 3716 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1677677812
transform 1 0 3764 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1677677812
transform 1 0 3716 0 1 4305
box -3 -3 3 3
use M2_M1  M2_M1_773
timestamp 1677677812
transform 1 0 3852 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1677677812
transform 1 0 3860 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_577
timestamp 1677677812
transform 1 0 3892 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_593
timestamp 1677677812
transform 1 0 3900 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_620
timestamp 1677677812
transform 1 0 3884 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_774
timestamp 1677677812
transform 1 0 3884 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_775
timestamp 1677677812
transform 1 0 3900 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1677677812
transform 1 0 3876 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1677677812
transform 1 0 3892 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1677677812
transform 1 0 3924 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1677677812
transform 1 0 3956 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_777
timestamp 1677677812
transform 1 0 3964 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_594
timestamp 1677677812
transform 1 0 3988 0 1 4355
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1677677812
transform 1 0 4004 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_778
timestamp 1677677812
transform 1 0 3988 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1677677812
transform 1 0 4004 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1677677812
transform 1 0 4020 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1677677812
transform 1 0 3996 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1677677812
transform 1 0 4012 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1677677812
transform 1 0 4028 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_622
timestamp 1677677812
transform 1 0 4068 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_781
timestamp 1677677812
transform 1 0 4116 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1677677812
transform 1 0 4068 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_720
timestamp 1677677812
transform 1 0 4084 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1677677812
transform 1 0 4132 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_623
timestamp 1677677812
transform 1 0 4156 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_782
timestamp 1677677812
transform 1 0 4140 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1677677812
transform 1 0 4132 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_643
timestamp 1677677812
transform 1 0 4148 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_783
timestamp 1677677812
transform 1 0 4156 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_784
timestamp 1677677812
transform 1 0 4172 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_897
timestamp 1677677812
transform 1 0 4164 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_736
timestamp 1677677812
transform 1 0 4172 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1677677812
transform 1 0 4188 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_624
timestamp 1677677812
transform 1 0 4228 0 1 4345
box -3 -3 3 3
use M2_M1  M2_M1_785
timestamp 1677677812
transform 1 0 4204 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1677677812
transform 1 0 4228 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_675
timestamp 1677677812
transform 1 0 4268 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_644
timestamp 1677677812
transform 1 0 4292 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_899
timestamp 1677677812
transform 1 0 4284 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_728
timestamp 1677677812
transform 1 0 4268 0 1 4295
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1677677812
transform 1 0 4300 0 1 4355
box -3 -3 3 3
use M2_M1  M2_M1_786
timestamp 1677677812
transform 1 0 4300 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_721
timestamp 1677677812
transform 1 0 4300 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_645
timestamp 1677677812
transform 1 0 4324 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_900
timestamp 1677677812
transform 1 0 4316 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_901
timestamp 1677677812
transform 1 0 4324 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_696
timestamp 1677677812
transform 1 0 4316 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_579
timestamp 1677677812
transform 1 0 4348 0 1 4365
box -3 -3 3 3
use M3_M2  M3_M2_646
timestamp 1677677812
transform 1 0 4356 0 1 4335
box -3 -3 3 3
use M3_M2  M3_M2_647
timestamp 1677677812
transform 1 0 4396 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_787
timestamp 1677677812
transform 1 0 4420 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1677677812
transform 1 0 4396 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_676
timestamp 1677677812
transform 1 0 4420 0 1 4325
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1677677812
transform 1 0 4348 0 1 4315
box -3 -3 3 3
use M3_M2  M3_M2_722
timestamp 1677677812
transform 1 0 4396 0 1 4305
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1677677812
transform 1 0 4380 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1677677812
transform 1 0 4412 0 1 4285
box -3 -3 3 3
use M3_M2  M3_M2_580
timestamp 1677677812
transform 1 0 4444 0 1 4365
box -3 -3 3 3
use M2_M1  M2_M1_788
timestamp 1677677812
transform 1 0 4452 0 1 4335
box -2 -2 2 2
use M3_M2  M3_M2_677
timestamp 1677677812
transform 1 0 4452 0 1 4325
box -3 -3 3 3
use M2_M1  M2_M1_789
timestamp 1677677812
transform 1 0 4540 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_903
timestamp 1677677812
transform 1 0 4476 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_904
timestamp 1677677812
transform 1 0 4532 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_905
timestamp 1677677812
transform 1 0 4548 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_790
timestamp 1677677812
transform 1 0 4572 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1677677812
transform 1 0 4564 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_907
timestamp 1677677812
transform 1 0 4580 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_648
timestamp 1677677812
transform 1 0 4596 0 1 4335
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1677677812
transform 1 0 4604 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1677677812
transform 1 0 4596 0 1 4325
box -2 -2 2 2
use M3_M2  M3_M2_698
timestamp 1677677812
transform 1 0 4596 0 1 4315
box -3 -3 3 3
use M2_M1  M2_M1_792
timestamp 1677677812
transform 1 0 4684 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_793
timestamp 1677677812
transform 1 0 4700 0 1 4335
box -2 -2 2 2
use M2_M1  M2_M1_909
timestamp 1677677812
transform 1 0 4724 0 1 4325
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1677677812
transform 1 0 4780 0 1 4325
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_8
timestamp 1677677812
transform 1 0 24 0 1 4270
box -10 -3 10 3
use FILL  FILL_419
timestamp 1677677812
transform 1 0 72 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_36
timestamp 1677677812
transform 1 0 80 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_41
timestamp 1677677812
transform -1 0 192 0 -1 4370
box -9 -3 26 105
use FILL  FILL_420
timestamp 1677677812
transform 1 0 192 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_23
timestamp 1677677812
transform -1 0 240 0 -1 4370
box -8 -3 46 105
use FILL  FILL_421
timestamp 1677677812
transform 1 0 240 0 -1 4370
box -8 -3 16 105
use FILL  FILL_422
timestamp 1677677812
transform 1 0 248 0 -1 4370
box -8 -3 16 105
use FILL  FILL_423
timestamp 1677677812
transform 1 0 256 0 -1 4370
box -8 -3 16 105
use FILL  FILL_424
timestamp 1677677812
transform 1 0 264 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_22
timestamp 1677677812
transform -1 0 312 0 -1 4370
box -8 -3 46 105
use FILL  FILL_425
timestamp 1677677812
transform 1 0 312 0 -1 4370
box -8 -3 16 105
use FILL  FILL_438
timestamp 1677677812
transform 1 0 320 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1677677812
transform -1 0 424 0 -1 4370
box -8 -3 104 105
use FILL  FILL_439
timestamp 1677677812
transform 1 0 424 0 -1 4370
box -8 -3 16 105
use FILL  FILL_441
timestamp 1677677812
transform 1 0 432 0 -1 4370
box -8 -3 16 105
use FILL  FILL_449
timestamp 1677677812
transform 1 0 440 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1677677812
transform 1 0 448 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_43
timestamp 1677677812
transform -1 0 560 0 -1 4370
box -9 -3 26 105
use FILL  FILL_450
timestamp 1677677812
transform 1 0 560 0 -1 4370
box -8 -3 16 105
use FILL  FILL_451
timestamp 1677677812
transform 1 0 568 0 -1 4370
box -8 -3 16 105
use FILL  FILL_453
timestamp 1677677812
transform 1 0 576 0 -1 4370
box -8 -3 16 105
use FILL  FILL_458
timestamp 1677677812
transform 1 0 584 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_26
timestamp 1677677812
transform -1 0 632 0 -1 4370
box -8 -3 46 105
use FILL  FILL_459
timestamp 1677677812
transform 1 0 632 0 -1 4370
box -8 -3 16 105
use FILL  FILL_460
timestamp 1677677812
transform 1 0 640 0 -1 4370
box -8 -3 16 105
use FILL  FILL_461
timestamp 1677677812
transform 1 0 648 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_44
timestamp 1677677812
transform 1 0 656 0 -1 4370
box -9 -3 26 105
use FILL  FILL_465
timestamp 1677677812
transform 1 0 672 0 -1 4370
box -8 -3 16 105
use FILL  FILL_467
timestamp 1677677812
transform 1 0 680 0 -1 4370
box -8 -3 16 105
use FILL  FILL_470
timestamp 1677677812
transform 1 0 688 0 -1 4370
box -8 -3 16 105
use FILL  FILL_471
timestamp 1677677812
transform 1 0 696 0 -1 4370
box -8 -3 16 105
use FILL  FILL_472
timestamp 1677677812
transform 1 0 704 0 -1 4370
box -8 -3 16 105
use FILL  FILL_473
timestamp 1677677812
transform 1 0 712 0 -1 4370
box -8 -3 16 105
use FILL  FILL_474
timestamp 1677677812
transform 1 0 720 0 -1 4370
box -8 -3 16 105
use FILL  FILL_475
timestamp 1677677812
transform 1 0 728 0 -1 4370
box -8 -3 16 105
use FILL  FILL_476
timestamp 1677677812
transform 1 0 736 0 -1 4370
box -8 -3 16 105
use FILL  FILL_477
timestamp 1677677812
transform 1 0 744 0 -1 4370
box -8 -3 16 105
use FILL  FILL_478
timestamp 1677677812
transform 1 0 752 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_45
timestamp 1677677812
transform 1 0 760 0 -1 4370
box -9 -3 26 105
use FILL  FILL_479
timestamp 1677677812
transform 1 0 776 0 -1 4370
box -8 -3 16 105
use FILL  FILL_480
timestamp 1677677812
transform 1 0 784 0 -1 4370
box -8 -3 16 105
use FILL  FILL_481
timestamp 1677677812
transform 1 0 792 0 -1 4370
box -8 -3 16 105
use FILL  FILL_490
timestamp 1677677812
transform 1 0 800 0 -1 4370
box -8 -3 16 105
use FILL  FILL_491
timestamp 1677677812
transform 1 0 808 0 -1 4370
box -8 -3 16 105
use FILL  FILL_492
timestamp 1677677812
transform 1 0 816 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1677677812
transform 1 0 824 0 -1 4370
box -8 -3 104 105
use FILL  FILL_493
timestamp 1677677812
transform 1 0 920 0 -1 4370
box -8 -3 16 105
use FILL  FILL_500
timestamp 1677677812
transform 1 0 928 0 -1 4370
box -8 -3 16 105
use FILL  FILL_501
timestamp 1677677812
transform 1 0 936 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_47
timestamp 1677677812
transform -1 0 960 0 -1 4370
box -9 -3 26 105
use M3_M2  M3_M2_739
timestamp 1677677812
transform 1 0 972 0 1 4275
box -3 -3 3 3
use FILL  FILL_502
timestamp 1677677812
transform 1 0 960 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_28
timestamp 1677677812
transform 1 0 968 0 -1 4370
box -8 -3 46 105
use FILL  FILL_503
timestamp 1677677812
transform 1 0 1008 0 -1 4370
box -8 -3 16 105
use FILL  FILL_504
timestamp 1677677812
transform 1 0 1016 0 -1 4370
box -8 -3 16 105
use FILL  FILL_505
timestamp 1677677812
transform 1 0 1024 0 -1 4370
box -8 -3 16 105
use FILL  FILL_506
timestamp 1677677812
transform 1 0 1032 0 -1 4370
box -8 -3 16 105
use FILL  FILL_507
timestamp 1677677812
transform 1 0 1040 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_13
timestamp 1677677812
transform 1 0 1048 0 -1 4370
box -8 -3 34 105
use FILL  FILL_508
timestamp 1677677812
transform 1 0 1080 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_29
timestamp 1677677812
transform 1 0 1088 0 -1 4370
box -8 -3 46 105
use FILL  FILL_509
timestamp 1677677812
transform 1 0 1128 0 -1 4370
box -8 -3 16 105
use FILL  FILL_511
timestamp 1677677812
transform 1 0 1136 0 -1 4370
box -8 -3 16 105
use FILL  FILL_513
timestamp 1677677812
transform 1 0 1144 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_49
timestamp 1677677812
transform 1 0 1152 0 -1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1677677812
transform -1 0 1264 0 -1 4370
box -8 -3 104 105
use FILL  FILL_523
timestamp 1677677812
transform 1 0 1264 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_17
timestamp 1677677812
transform -1 0 1304 0 -1 4370
box -8 -3 34 105
use FILL  FILL_524
timestamp 1677677812
transform 1 0 1304 0 -1 4370
box -8 -3 16 105
use FILL  FILL_525
timestamp 1677677812
transform 1 0 1312 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1677677812
transform 1 0 1320 0 -1 4370
box -8 -3 104 105
use FILL  FILL_526
timestamp 1677677812
transform 1 0 1416 0 -1 4370
box -8 -3 16 105
use FILL  FILL_527
timestamp 1677677812
transform 1 0 1424 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_50
timestamp 1677677812
transform 1 0 1432 0 -1 4370
box -9 -3 26 105
use FILL  FILL_528
timestamp 1677677812
transform 1 0 1448 0 -1 4370
box -8 -3 16 105
use FILL  FILL_532
timestamp 1677677812
transform 1 0 1456 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_25
timestamp 1677677812
transform -1 0 1504 0 -1 4370
box -8 -3 46 105
use FILL  FILL_533
timestamp 1677677812
transform 1 0 1504 0 -1 4370
box -8 -3 16 105
use FILL  FILL_534
timestamp 1677677812
transform 1 0 1512 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_52
timestamp 1677677812
transform 1 0 1520 0 -1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1677677812
transform -1 0 1632 0 -1 4370
box -8 -3 104 105
use FILL  FILL_538
timestamp 1677677812
transform 1 0 1632 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_740
timestamp 1677677812
transform 1 0 1660 0 1 4275
box -3 -3 3 3
use FILL  FILL_539
timestamp 1677677812
transform 1 0 1640 0 -1 4370
box -8 -3 16 105
use FILL  FILL_540
timestamp 1677677812
transform 1 0 1648 0 -1 4370
box -8 -3 16 105
use FILL  FILL_542
timestamp 1677677812
transform 1 0 1656 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1677677812
transform 1 0 1664 0 -1 4370
box -8 -3 104 105
use FILL  FILL_552
timestamp 1677677812
transform 1 0 1760 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_54
timestamp 1677677812
transform -1 0 1784 0 -1 4370
box -9 -3 26 105
use FILL  FILL_553
timestamp 1677677812
transform 1 0 1784 0 -1 4370
box -8 -3 16 105
use FILL  FILL_555
timestamp 1677677812
transform 1 0 1792 0 -1 4370
box -8 -3 16 105
use FILL  FILL_560
timestamp 1677677812
transform 1 0 1800 0 -1 4370
box -8 -3 16 105
use FILL  FILL_561
timestamp 1677677812
transform 1 0 1808 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_741
timestamp 1677677812
transform 1 0 1828 0 1 4275
box -3 -3 3 3
use FILL  FILL_562
timestamp 1677677812
transform 1 0 1816 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_31
timestamp 1677677812
transform 1 0 1824 0 -1 4370
box -8 -3 46 105
use FILL  FILL_563
timestamp 1677677812
transform 1 0 1864 0 -1 4370
box -8 -3 16 105
use FILL  FILL_565
timestamp 1677677812
transform 1 0 1872 0 -1 4370
box -8 -3 16 105
use FILL  FILL_570
timestamp 1677677812
transform 1 0 1880 0 -1 4370
box -8 -3 16 105
use FILL  FILL_571
timestamp 1677677812
transform 1 0 1888 0 -1 4370
box -8 -3 16 105
use FILL  FILL_572
timestamp 1677677812
transform 1 0 1896 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_28
timestamp 1677677812
transform 1 0 1904 0 -1 4370
box -8 -3 46 105
use FILL  FILL_573
timestamp 1677677812
transform 1 0 1944 0 -1 4370
box -8 -3 16 105
use FILL  FILL_575
timestamp 1677677812
transform 1 0 1952 0 -1 4370
box -8 -3 16 105
use FILL  FILL_577
timestamp 1677677812
transform 1 0 1960 0 -1 4370
box -8 -3 16 105
use FILL  FILL_579
timestamp 1677677812
transform 1 0 1968 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_56
timestamp 1677677812
transform 1 0 1976 0 -1 4370
box -9 -3 26 105
use INVX2  INVX2_57
timestamp 1677677812
transform 1 0 1992 0 -1 4370
box -9 -3 26 105
use FILL  FILL_584
timestamp 1677677812
transform 1 0 2008 0 -1 4370
box -8 -3 16 105
use FILL  FILL_585
timestamp 1677677812
transform 1 0 2016 0 -1 4370
box -8 -3 16 105
use FILL  FILL_586
timestamp 1677677812
transform 1 0 2024 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_58
timestamp 1677677812
transform 1 0 2032 0 -1 4370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1677677812
transform -1 0 2144 0 -1 4370
box -8 -3 104 105
use FILL  FILL_587
timestamp 1677677812
transform 1 0 2144 0 -1 4370
box -8 -3 16 105
use FILL  FILL_588
timestamp 1677677812
transform 1 0 2152 0 -1 4370
box -8 -3 16 105
use FILL  FILL_589
timestamp 1677677812
transform 1 0 2160 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_59
timestamp 1677677812
transform -1 0 2184 0 -1 4370
box -9 -3 26 105
use FILL  FILL_590
timestamp 1677677812
transform 1 0 2184 0 -1 4370
box -8 -3 16 105
use FILL  FILL_591
timestamp 1677677812
transform 1 0 2192 0 -1 4370
box -8 -3 16 105
use FILL  FILL_592
timestamp 1677677812
transform 1 0 2200 0 -1 4370
box -8 -3 16 105
use FILL  FILL_593
timestamp 1677677812
transform 1 0 2208 0 -1 4370
box -8 -3 16 105
use FILL  FILL_594
timestamp 1677677812
transform 1 0 2216 0 -1 4370
box -8 -3 16 105
use FILL  FILL_595
timestamp 1677677812
transform 1 0 2224 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_33
timestamp 1677677812
transform -1 0 2272 0 -1 4370
box -8 -3 46 105
use FILL  FILL_596
timestamp 1677677812
transform 1 0 2272 0 -1 4370
box -8 -3 16 105
use FILL  FILL_597
timestamp 1677677812
transform 1 0 2280 0 -1 4370
box -8 -3 16 105
use FILL  FILL_598
timestamp 1677677812
transform 1 0 2288 0 -1 4370
box -8 -3 16 105
use FILL  FILL_602
timestamp 1677677812
transform 1 0 2296 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_34
timestamp 1677677812
transform 1 0 2304 0 -1 4370
box -8 -3 46 105
use FILL  FILL_603
timestamp 1677677812
transform 1 0 2344 0 -1 4370
box -8 -3 16 105
use FILL  FILL_604
timestamp 1677677812
transform 1 0 2352 0 -1 4370
box -8 -3 16 105
use FILL  FILL_605
timestamp 1677677812
transform 1 0 2360 0 -1 4370
box -8 -3 16 105
use FILL  FILL_606
timestamp 1677677812
transform 1 0 2368 0 -1 4370
box -8 -3 16 105
use FILL  FILL_607
timestamp 1677677812
transform 1 0 2376 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_35
timestamp 1677677812
transform 1 0 2384 0 -1 4370
box -8 -3 46 105
use FILL  FILL_608
timestamp 1677677812
transform 1 0 2424 0 -1 4370
box -8 -3 16 105
use FILL  FILL_609
timestamp 1677677812
transform 1 0 2432 0 -1 4370
box -8 -3 16 105
use FILL  FILL_610
timestamp 1677677812
transform 1 0 2440 0 -1 4370
box -8 -3 16 105
use FILL  FILL_611
timestamp 1677677812
transform 1 0 2448 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_30
timestamp 1677677812
transform -1 0 2496 0 -1 4370
box -8 -3 46 105
use FILL  FILL_612
timestamp 1677677812
transform 1 0 2496 0 -1 4370
box -8 -3 16 105
use FILL  FILL_613
timestamp 1677677812
transform 1 0 2504 0 -1 4370
box -8 -3 16 105
use FILL  FILL_614
timestamp 1677677812
transform 1 0 2512 0 -1 4370
box -8 -3 16 105
use FILL  FILL_615
timestamp 1677677812
transform 1 0 2520 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_36
timestamp 1677677812
transform 1 0 2528 0 -1 4370
box -8 -3 46 105
use FILL  FILL_621
timestamp 1677677812
transform 1 0 2568 0 -1 4370
box -8 -3 16 105
use FILL  FILL_622
timestamp 1677677812
transform 1 0 2576 0 -1 4370
box -8 -3 16 105
use FILL  FILL_623
timestamp 1677677812
transform 1 0 2584 0 -1 4370
box -8 -3 16 105
use FILL  FILL_624
timestamp 1677677812
transform 1 0 2592 0 -1 4370
box -8 -3 16 105
use AOI22X1  AOI22X1_37
timestamp 1677677812
transform 1 0 2600 0 -1 4370
box -8 -3 46 105
use FILL  FILL_625
timestamp 1677677812
transform 1 0 2640 0 -1 4370
box -8 -3 16 105
use FILL  FILL_626
timestamp 1677677812
transform 1 0 2648 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_62
timestamp 1677677812
transform 1 0 2656 0 -1 4370
box -9 -3 26 105
use FILL  FILL_627
timestamp 1677677812
transform 1 0 2672 0 -1 4370
box -8 -3 16 105
use FILL  FILL_630
timestamp 1677677812
transform 1 0 2680 0 -1 4370
box -8 -3 16 105
use FILL  FILL_631
timestamp 1677677812
transform 1 0 2688 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_54
timestamp 1677677812
transform 1 0 2696 0 -1 4370
box -8 -3 104 105
use FILL  FILL_632
timestamp 1677677812
transform 1 0 2792 0 -1 4370
box -8 -3 16 105
use FILL  FILL_633
timestamp 1677677812
transform 1 0 2800 0 -1 4370
box -8 -3 16 105
use FILL  FILL_635
timestamp 1677677812
transform 1 0 2808 0 -1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_8
timestamp 1677677812
transform 1 0 2816 0 -1 4370
box -8 -3 32 105
use FILL  FILL_641
timestamp 1677677812
transform 1 0 2840 0 -1 4370
box -8 -3 16 105
use FILL  FILL_642
timestamp 1677677812
transform 1 0 2848 0 -1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_9
timestamp 1677677812
transform 1 0 2856 0 -1 4370
box -8 -3 32 105
use FILL  FILL_643
timestamp 1677677812
transform 1 0 2880 0 -1 4370
box -8 -3 16 105
use FILL  FILL_644
timestamp 1677677812
transform 1 0 2888 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_20
timestamp 1677677812
transform 1 0 2896 0 -1 4370
box -8 -3 34 105
use FILL  FILL_645
timestamp 1677677812
transform 1 0 2928 0 -1 4370
box -8 -3 16 105
use FILL  FILL_646
timestamp 1677677812
transform 1 0 2936 0 -1 4370
box -8 -3 16 105
use NOR2X1  NOR2X1_10
timestamp 1677677812
transform 1 0 2944 0 -1 4370
box -8 -3 32 105
use FILL  FILL_651
timestamp 1677677812
transform 1 0 2968 0 -1 4370
box -8 -3 16 105
use FILL  FILL_652
timestamp 1677677812
transform 1 0 2976 0 -1 4370
box -8 -3 16 105
use FILL  FILL_653
timestamp 1677677812
transform 1 0 2984 0 -1 4370
box -8 -3 16 105
use FILL  FILL_654
timestamp 1677677812
transform 1 0 2992 0 -1 4370
box -8 -3 16 105
use FILL  FILL_655
timestamp 1677677812
transform 1 0 3000 0 -1 4370
box -8 -3 16 105
use OAI21X1  OAI21X1_23
timestamp 1677677812
transform -1 0 3040 0 -1 4370
box -8 -3 34 105
use FILL  FILL_657
timestamp 1677677812
transform 1 0 3040 0 -1 4370
box -8 -3 16 105
use FILL  FILL_659
timestamp 1677677812
transform 1 0 3048 0 -1 4370
box -8 -3 16 105
use FILL  FILL_661
timestamp 1677677812
transform 1 0 3056 0 -1 4370
box -8 -3 16 105
use FILL  FILL_669
timestamp 1677677812
transform 1 0 3064 0 -1 4370
box -8 -3 16 105
use FILL  FILL_670
timestamp 1677677812
transform 1 0 3072 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_56
timestamp 1677677812
transform 1 0 3080 0 -1 4370
box -8 -3 104 105
use INVX2  INVX2_65
timestamp 1677677812
transform 1 0 3176 0 -1 4370
box -9 -3 26 105
use FILL  FILL_671
timestamp 1677677812
transform 1 0 3192 0 -1 4370
box -8 -3 16 105
use FILL  FILL_672
timestamp 1677677812
transform 1 0 3200 0 -1 4370
box -8 -3 16 105
use FILL  FILL_673
timestamp 1677677812
transform 1 0 3208 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_32
timestamp 1677677812
transform 1 0 3216 0 -1 4370
box -8 -3 46 105
use FILL  FILL_674
timestamp 1677677812
transform 1 0 3256 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_742
timestamp 1677677812
transform 1 0 3276 0 1 4275
box -3 -3 3 3
use FILL  FILL_675
timestamp 1677677812
transform 1 0 3264 0 -1 4370
box -8 -3 16 105
use FILL  FILL_679
timestamp 1677677812
transform 1 0 3272 0 -1 4370
box -8 -3 16 105
use FILL  FILL_680
timestamp 1677677812
transform 1 0 3280 0 -1 4370
box -8 -3 16 105
use FILL  FILL_681
timestamp 1677677812
transform 1 0 3288 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_58
timestamp 1677677812
transform 1 0 3296 0 -1 4370
box -8 -3 104 105
use FILL  FILL_682
timestamp 1677677812
transform 1 0 3392 0 -1 4370
box -8 -3 16 105
use FILL  FILL_683
timestamp 1677677812
transform 1 0 3400 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_60
timestamp 1677677812
transform 1 0 3408 0 -1 4370
box -8 -3 104 105
use FILL  FILL_690
timestamp 1677677812
transform 1 0 3504 0 -1 4370
box -8 -3 16 105
use FILL  FILL_691
timestamp 1677677812
transform 1 0 3512 0 -1 4370
box -8 -3 16 105
use FILL  FILL_692
timestamp 1677677812
transform 1 0 3520 0 -1 4370
box -8 -3 16 105
use FILL  FILL_693
timestamp 1677677812
transform 1 0 3528 0 -1 4370
box -8 -3 16 105
use FILL  FILL_694
timestamp 1677677812
transform 1 0 3536 0 -1 4370
box -8 -3 16 105
use FILL  FILL_695
timestamp 1677677812
transform 1 0 3544 0 -1 4370
box -8 -3 16 105
use FILL  FILL_696
timestamp 1677677812
transform 1 0 3552 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_743
timestamp 1677677812
transform 1 0 3588 0 1 4275
box -3 -3 3 3
use INVX2  INVX2_67
timestamp 1677677812
transform 1 0 3560 0 -1 4370
box -9 -3 26 105
use FILL  FILL_697
timestamp 1677677812
transform 1 0 3576 0 -1 4370
box -8 -3 16 105
use FILL  FILL_698
timestamp 1677677812
transform 1 0 3584 0 -1 4370
box -8 -3 16 105
use FILL  FILL_699
timestamp 1677677812
transform 1 0 3592 0 -1 4370
box -8 -3 16 105
use FILL  FILL_700
timestamp 1677677812
transform 1 0 3600 0 -1 4370
box -8 -3 16 105
use FILL  FILL_701
timestamp 1677677812
transform 1 0 3608 0 -1 4370
box -8 -3 16 105
use FILL  FILL_703
timestamp 1677677812
transform 1 0 3616 0 -1 4370
box -8 -3 16 105
use FILL  FILL_705
timestamp 1677677812
transform 1 0 3624 0 -1 4370
box -8 -3 16 105
use FILL  FILL_707
timestamp 1677677812
transform 1 0 3632 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_33
timestamp 1677677812
transform 1 0 3640 0 -1 4370
box -8 -3 46 105
use FILL  FILL_714
timestamp 1677677812
transform 1 0 3680 0 -1 4370
box -8 -3 16 105
use FILL  FILL_716
timestamp 1677677812
transform 1 0 3688 0 -1 4370
box -8 -3 16 105
use FILL  FILL_718
timestamp 1677677812
transform 1 0 3696 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_61
timestamp 1677677812
transform 1 0 3704 0 -1 4370
box -8 -3 104 105
use FILL  FILL_729
timestamp 1677677812
transform 1 0 3800 0 -1 4370
box -8 -3 16 105
use FILL  FILL_730
timestamp 1677677812
transform 1 0 3808 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_69
timestamp 1677677812
transform 1 0 3816 0 -1 4370
box -9 -3 26 105
use FILL  FILL_731
timestamp 1677677812
transform 1 0 3832 0 -1 4370
box -8 -3 16 105
use FILL  FILL_736
timestamp 1677677812
transform 1 0 3840 0 -1 4370
box -8 -3 16 105
use FILL  FILL_737
timestamp 1677677812
transform 1 0 3848 0 -1 4370
box -8 -3 16 105
use FILL  FILL_738
timestamp 1677677812
transform 1 0 3856 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_34
timestamp 1677677812
transform -1 0 3904 0 -1 4370
box -8 -3 46 105
use FILL  FILL_739
timestamp 1677677812
transform 1 0 3904 0 -1 4370
box -8 -3 16 105
use FILL  FILL_741
timestamp 1677677812
transform 1 0 3912 0 -1 4370
box -8 -3 16 105
use FILL  FILL_744
timestamp 1677677812
transform 1 0 3920 0 -1 4370
box -8 -3 16 105
use FILL  FILL_745
timestamp 1677677812
transform 1 0 3928 0 -1 4370
box -8 -3 16 105
use FILL  FILL_746
timestamp 1677677812
transform 1 0 3936 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_70
timestamp 1677677812
transform -1 0 3960 0 -1 4370
box -9 -3 26 105
use FILL  FILL_747
timestamp 1677677812
transform 1 0 3960 0 -1 4370
box -8 -3 16 105
use FILL  FILL_749
timestamp 1677677812
transform 1 0 3968 0 -1 4370
box -8 -3 16 105
use FILL  FILL_769
timestamp 1677677812
transform 1 0 3976 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_35
timestamp 1677677812
transform -1 0 4024 0 -1 4370
box -8 -3 46 105
use FILL  FILL_770
timestamp 1677677812
transform 1 0 4024 0 -1 4370
box -8 -3 16 105
use M3_M2  M3_M2_744
timestamp 1677677812
transform 1 0 4132 0 1 4275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_63
timestamp 1677677812
transform -1 0 4128 0 -1 4370
box -8 -3 104 105
use FILL  FILL_771
timestamp 1677677812
transform 1 0 4128 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_36
timestamp 1677677812
transform 1 0 4136 0 -1 4370
box -8 -3 46 105
use FILL  FILL_772
timestamp 1677677812
transform 1 0 4176 0 -1 4370
box -8 -3 16 105
use FILL  FILL_773
timestamp 1677677812
transform 1 0 4184 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_64
timestamp 1677677812
transform 1 0 4192 0 -1 4370
box -8 -3 104 105
use FILL  FILL_774
timestamp 1677677812
transform 1 0 4288 0 -1 4370
box -8 -3 16 105
use FILL  FILL_775
timestamp 1677677812
transform 1 0 4296 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_75
timestamp 1677677812
transform 1 0 4304 0 -1 4370
box -9 -3 26 105
use FILL  FILL_776
timestamp 1677677812
transform 1 0 4320 0 -1 4370
box -8 -3 16 105
use FILL  FILL_787
timestamp 1677677812
transform 1 0 4328 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_65
timestamp 1677677812
transform -1 0 4432 0 -1 4370
box -8 -3 104 105
use FILL  FILL_788
timestamp 1677677812
transform 1 0 4432 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_66
timestamp 1677677812
transform 1 0 4440 0 -1 4370
box -8 -3 104 105
use FILL  FILL_789
timestamp 1677677812
transform 1 0 4536 0 -1 4370
box -8 -3 16 105
use FILL  FILL_796
timestamp 1677677812
transform 1 0 4544 0 -1 4370
box -8 -3 16 105
use OAI22X1  OAI22X1_40
timestamp 1677677812
transform 1 0 4552 0 -1 4370
box -8 -3 46 105
use FILL  FILL_797
timestamp 1677677812
transform 1 0 4592 0 -1 4370
box -8 -3 16 105
use FILL  FILL_798
timestamp 1677677812
transform 1 0 4600 0 -1 4370
box -8 -3 16 105
use FILL  FILL_799
timestamp 1677677812
transform 1 0 4608 0 -1 4370
box -8 -3 16 105
use FILL  FILL_800
timestamp 1677677812
transform 1 0 4616 0 -1 4370
box -8 -3 16 105
use INVX2  INVX2_78
timestamp 1677677812
transform -1 0 4640 0 -1 4370
box -9 -3 26 105
use FILL  FILL_801
timestamp 1677677812
transform 1 0 4640 0 -1 4370
box -8 -3 16 105
use FILL  FILL_803
timestamp 1677677812
transform 1 0 4648 0 -1 4370
box -8 -3 16 105
use FILL  FILL_807
timestamp 1677677812
transform 1 0 4656 0 -1 4370
box -8 -3 16 105
use FILL  FILL_808
timestamp 1677677812
transform 1 0 4664 0 -1 4370
box -8 -3 16 105
use FILL  FILL_809
timestamp 1677677812
transform 1 0 4672 0 -1 4370
box -8 -3 16 105
use FILL  FILL_810
timestamp 1677677812
transform 1 0 4680 0 -1 4370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_68
timestamp 1677677812
transform 1 0 4688 0 -1 4370
box -8 -3 104 105
use FILL  FILL_811
timestamp 1677677812
transform 1 0 4784 0 -1 4370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_9
timestamp 1677677812
transform 1 0 4843 0 1 4270
box -10 -3 10 3
use M3_M2  M3_M2_788
timestamp 1677677812
transform 1 0 132 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1677677812
transform 1 0 172 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1677677812
transform 1 0 132 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_926
timestamp 1677677812
transform 1 0 164 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1677677812
transform 1 0 172 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1677677812
transform 1 0 84 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_878
timestamp 1677677812
transform 1 0 164 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1677677812
transform 1 0 204 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_791
timestamp 1677677812
transform 1 0 220 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_928
timestamp 1677677812
transform 1 0 212 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_792
timestamp 1677677812
transform 1 0 260 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_832
timestamp 1677677812
transform 1 0 236 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_929
timestamp 1677677812
transform 1 0 244 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_930
timestamp 1677677812
transform 1 0 260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1044
timestamp 1677677812
transform 1 0 228 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1677677812
transform 1 0 236 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1046
timestamp 1677677812
transform 1 0 252 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_863
timestamp 1677677812
transform 1 0 260 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1677677812
transform 1 0 252 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1677677812
transform 1 0 284 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1677677812
transform 1 0 308 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_795
timestamp 1677677812
transform 1 0 332 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_796
timestamp 1677677812
transform 1 0 372 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_833
timestamp 1677677812
transform 1 0 284 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_834
timestamp 1677677812
transform 1 0 324 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_931
timestamp 1677677812
transform 1 0 332 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_932
timestamp 1677677812
transform 1 0 364 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1677677812
transform 1 0 372 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1677677812
transform 1 0 284 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_880
timestamp 1677677812
transform 1 0 284 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1677677812
transform 1 0 364 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_934
timestamp 1677677812
transform 1 0 404 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_797
timestamp 1677677812
transform 1 0 420 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_935
timestamp 1677677812
transform 1 0 420 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_835
timestamp 1677677812
transform 1 0 428 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_936
timestamp 1677677812
transform 1 0 436 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1677677812
transform 1 0 420 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1677677812
transform 1 0 428 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1677677812
transform 1 0 444 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1677677812
transform 1 0 452 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_882
timestamp 1677677812
transform 1 0 444 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_836
timestamp 1677677812
transform 1 0 468 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_837
timestamp 1677677812
transform 1 0 484 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_937
timestamp 1677677812
transform 1 0 508 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1677677812
transform 1 0 484 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1053
timestamp 1677677812
transform 1 0 572 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1677677812
transform 1 0 588 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_864
timestamp 1677677812
transform 1 0 588 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_918
timestamp 1677677812
transform 1 0 580 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_798
timestamp 1677677812
transform 1 0 604 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_939
timestamp 1677677812
transform 1 0 604 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_940
timestamp 1677677812
transform 1 0 620 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1677677812
transform 1 0 636 0 1 4214
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1677677812
transform 1 0 644 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1677677812
transform 1 0 604 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_865
timestamp 1677677812
transform 1 0 620 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1677677812
transform 1 0 644 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1055
timestamp 1677677812
transform 1 0 668 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_884
timestamp 1677677812
transform 1 0 668 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_942
timestamp 1677677812
transform 1 0 684 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1677677812
transform 1 0 700 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1677677812
transform 1 0 692 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_866
timestamp 1677677812
transform 1 0 700 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_766
timestamp 1677677812
transform 1 0 716 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_1057
timestamp 1677677812
transform 1 0 708 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_885
timestamp 1677677812
transform 1 0 708 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1677677812
transform 1 0 780 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_944
timestamp 1677677812
transform 1 0 788 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_839
timestamp 1677677812
transform 1 0 820 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1058
timestamp 1677677812
transform 1 0 820 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_799
timestamp 1677677812
transform 1 0 908 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_800
timestamp 1677677812
transform 1 0 948 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_945
timestamp 1677677812
transform 1 0 908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_946
timestamp 1677677812
transform 1 0 940 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_947
timestamp 1677677812
transform 1 0 948 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1677677812
transform 1 0 860 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_886
timestamp 1677677812
transform 1 0 924 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1060
timestamp 1677677812
transform 1 0 948 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_887
timestamp 1677677812
transform 1 0 948 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_774
timestamp 1677677812
transform 1 0 972 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_867
timestamp 1677677812
transform 1 0 972 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1152
timestamp 1677677812
transform 1 0 972 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1677677812
transform 1 0 988 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1677677812
transform 1 0 1028 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_840
timestamp 1677677812
transform 1 0 1036 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1062
timestamp 1677677812
transform 1 0 1036 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_949
timestamp 1677677812
transform 1 0 1060 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_775
timestamp 1677677812
transform 1 0 1132 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_917
timestamp 1677677812
transform 1 0 1100 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_950
timestamp 1677677812
transform 1 0 1092 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1677677812
transform 1 0 1084 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_801
timestamp 1677677812
transform 1 0 1108 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_951
timestamp 1677677812
transform 1 0 1108 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1677677812
transform 1 0 1124 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_888
timestamp 1677677812
transform 1 0 1100 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_919
timestamp 1677677812
transform 1 0 1092 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_841
timestamp 1677677812
transform 1 0 1132 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_953
timestamp 1677677812
transform 1 0 1140 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1064
timestamp 1677677812
transform 1 0 1116 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1677677812
transform 1 0 1132 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1677677812
transform 1 0 1140 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_954
timestamp 1677677812
transform 1 0 1156 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_776
timestamp 1677677812
transform 1 0 1180 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_918
timestamp 1677677812
transform 1 0 1276 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1677677812
transform 1 0 1172 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1677677812
transform 1 0 1180 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1677677812
transform 1 0 1212 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_842
timestamp 1677677812
transform 1 0 1276 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_958
timestamp 1677677812
transform 1 0 1292 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_868
timestamp 1677677812
transform 1 0 1172 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_869
timestamp 1677677812
transform 1 0 1212 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1067
timestamp 1677677812
transform 1 0 1260 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1068
timestamp 1677677812
transform 1 0 1276 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_889
timestamp 1677677812
transform 1 0 1276 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1677677812
transform 1 0 1308 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_959
timestamp 1677677812
transform 1 0 1348 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_960
timestamp 1677677812
transform 1 0 1404 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1069
timestamp 1677677812
transform 1 0 1340 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_890
timestamp 1677677812
transform 1 0 1340 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1070
timestamp 1677677812
transform 1 0 1428 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_961
timestamp 1677677812
transform 1 0 1444 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_891
timestamp 1677677812
transform 1 0 1444 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_920
timestamp 1677677812
transform 1 0 1404 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_921
timestamp 1677677812
transform 1 0 1436 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_753
timestamp 1677677812
transform 1 0 1476 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_922
timestamp 1677677812
transform 1 0 1484 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1677677812
transform 1 0 1508 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1677677812
transform 1 0 1508 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_870
timestamp 1677677812
transform 1 0 1500 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_754
timestamp 1677677812
transform 1 0 1524 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1677677812
transform 1 0 1540 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1677677812
transform 1 0 1516 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_755
timestamp 1677677812
transform 1 0 1556 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_962
timestamp 1677677812
transform 1 0 1524 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_963
timestamp 1677677812
transform 1 0 1540 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_845
timestamp 1677677812
transform 1 0 1548 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1071
timestamp 1677677812
transform 1 0 1508 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1072
timestamp 1677677812
transform 1 0 1516 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1677677812
transform 1 0 1532 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_892
timestamp 1677677812
transform 1 0 1524 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1074
timestamp 1677677812
transform 1 0 1556 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1677677812
transform 1 0 1564 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1075
timestamp 1677677812
transform 1 0 1580 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1076
timestamp 1677677812
transform 1 0 1588 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1677677812
transform 1 0 1612 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1677677812
transform 1 0 1636 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_746
timestamp 1677677812
transform 1 0 1652 0 1 4265
box -3 -3 3 3
use M2_M1  M2_M1_967
timestamp 1677677812
transform 1 0 1652 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1077
timestamp 1677677812
transform 1 0 1652 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1677677812
transform 1 0 1660 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1677677812
transform 1 0 1668 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1677677812
transform 1 0 1676 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_893
timestamp 1677677812
transform 1 0 1668 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_923
timestamp 1677677812
transform 1 0 1676 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1079
timestamp 1677677812
transform 1 0 1684 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_779
timestamp 1677677812
transform 1 0 1780 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_970
timestamp 1677677812
transform 1 0 1780 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_846
timestamp 1677677812
transform 1 0 1804 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_971
timestamp 1677677812
transform 1 0 1812 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1677677812
transform 1 0 1732 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_924
timestamp 1677677812
transform 1 0 1748 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_972
timestamp 1677677812
transform 1 0 1828 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1677677812
transform 1 0 1820 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1677677812
transform 1 0 1860 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_847
timestamp 1677677812
transform 1 0 1868 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_780
timestamp 1677677812
transform 1 0 1884 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_974
timestamp 1677677812
transform 1 0 1876 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_975
timestamp 1677677812
transform 1 0 1884 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1677677812
transform 1 0 1868 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_894
timestamp 1677677812
transform 1 0 1860 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1083
timestamp 1677677812
transform 1 0 1892 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_756
timestamp 1677677812
transform 1 0 1924 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1677677812
transform 1 0 1932 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_976
timestamp 1677677812
transform 1 0 1924 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1677677812
transform 1 0 1924 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1677677812
transform 1 0 1932 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_895
timestamp 1677677812
transform 1 0 1924 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_977
timestamp 1677677812
transform 1 0 1948 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1677677812
transform 1 0 1988 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1677677812
transform 1 0 2004 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1677677812
transform 1 0 1980 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_896
timestamp 1677677812
transform 1 0 1980 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1087
timestamp 1677677812
transform 1 0 2020 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_897
timestamp 1677677812
transform 1 0 2036 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1088
timestamp 1677677812
transform 1 0 2052 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_898
timestamp 1677677812
transform 1 0 2060 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1089
timestamp 1677677812
transform 1 0 2148 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1677677812
transform 1 0 2156 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1677677812
transform 1 0 2212 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_981
timestamp 1677677812
transform 1 0 2212 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_747
timestamp 1677677812
transform 1 0 2228 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_781
timestamp 1677677812
transform 1 0 2300 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_804
timestamp 1677677812
transform 1 0 2252 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_982
timestamp 1677677812
transform 1 0 2252 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_983
timestamp 1677677812
transform 1 0 2308 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1677677812
transform 1 0 2228 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_848
timestamp 1677677812
transform 1 0 2316 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1091
timestamp 1677677812
transform 1 0 2316 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_748
timestamp 1677677812
transform 1 0 2364 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_757
timestamp 1677677812
transform 1 0 2356 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_984
timestamp 1677677812
transform 1 0 2332 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_985
timestamp 1677677812
transform 1 0 2356 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1092
timestamp 1677677812
transform 1 0 2348 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1093
timestamp 1677677812
transform 1 0 2364 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_758
timestamp 1677677812
transform 1 0 2404 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_986
timestamp 1677677812
transform 1 0 2420 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_759
timestamp 1677677812
transform 1 0 2468 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_987
timestamp 1677677812
transform 1 0 2484 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_782
timestamp 1677677812
transform 1 0 2588 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_988
timestamp 1677677812
transform 1 0 2564 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1677677812
transform 1 0 2620 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1677677812
transform 1 0 2540 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_783
timestamp 1677677812
transform 1 0 2636 0 1 4235
box -3 -3 3 3
use M2_M1  M2_M1_990
timestamp 1677677812
transform 1 0 2636 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1677677812
transform 1 0 2628 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_899
timestamp 1677677812
transform 1 0 2620 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_991
timestamp 1677677812
transform 1 0 2660 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_849
timestamp 1677677812
transform 1 0 2668 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_992
timestamp 1677677812
transform 1 0 2676 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1096
timestamp 1677677812
transform 1 0 2668 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1097
timestamp 1677677812
transform 1 0 2676 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_805
timestamp 1677677812
transform 1 0 2740 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_993
timestamp 1677677812
transform 1 0 2740 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_760
timestamp 1677677812
transform 1 0 2828 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_761
timestamp 1677677812
transform 1 0 2852 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1677677812
transform 1 0 2860 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_806
timestamp 1677677812
transform 1 0 2780 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_807
timestamp 1677677812
transform 1 0 2844 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_994
timestamp 1677677812
transform 1 0 2780 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_995
timestamp 1677677812
transform 1 0 2844 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_996
timestamp 1677677812
transform 1 0 2852 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1677677812
transform 1 0 2756 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1099
timestamp 1677677812
transform 1 0 2844 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_900
timestamp 1677677812
transform 1 0 2844 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_850
timestamp 1677677812
transform 1 0 2876 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_919
timestamp 1677677812
transform 1 0 2892 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_997
timestamp 1677677812
transform 1 0 2884 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1677677812
transform 1 0 2868 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1101
timestamp 1677677812
transform 1 0 2876 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_901
timestamp 1677677812
transform 1 0 2892 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_998
timestamp 1677677812
transform 1 0 2908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1677677812
transform 1 0 2932 0 1 4195
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1677677812
transform 1 0 2948 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_851
timestamp 1677677812
transform 1 0 2948 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1102
timestamp 1677677812
transform 1 0 2956 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1677677812
transform 1 0 2988 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1677677812
transform 1 0 2972 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_852
timestamp 1677677812
transform 1 0 2980 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1103
timestamp 1677677812
transform 1 0 2972 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1104
timestamp 1677677812
transform 1 0 2980 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_902
timestamp 1677677812
transform 1 0 2996 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_922
timestamp 1677677812
transform 1 0 3012 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_853
timestamp 1677677812
transform 1 0 3052 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1000
timestamp 1677677812
transform 1 0 3068 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1677677812
transform 1 0 3108 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1677677812
transform 1 0 3124 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1677677812
transform 1 0 3108 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1677677812
transform 1 0 3116 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1107
timestamp 1677677812
transform 1 0 3132 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1108
timestamp 1677677812
transform 1 0 3148 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1109
timestamp 1677677812
transform 1 0 3156 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_903
timestamp 1677677812
transform 1 0 3116 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_925
timestamp 1677677812
transform 1 0 3116 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_904
timestamp 1677677812
transform 1 0 3156 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_926
timestamp 1677677812
transform 1 0 3148 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1002
timestamp 1677677812
transform 1 0 3188 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_905
timestamp 1677677812
transform 1 0 3188 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1110
timestamp 1677677812
transform 1 0 3196 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_809
timestamp 1677677812
transform 1 0 3236 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_810
timestamp 1677677812
transform 1 0 3260 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1003
timestamp 1677677812
transform 1 0 3236 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1004
timestamp 1677677812
transform 1 0 3252 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1005
timestamp 1677677812
transform 1 0 3260 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1677677812
transform 1 0 3244 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_906
timestamp 1677677812
transform 1 0 3252 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_927
timestamp 1677677812
transform 1 0 3228 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_928
timestamp 1677677812
transform 1 0 3244 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1112
timestamp 1677677812
transform 1 0 3276 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_907
timestamp 1677677812
transform 1 0 3276 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_929
timestamp 1677677812
transform 1 0 3308 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_854
timestamp 1677677812
transform 1 0 3348 0 1 4215
box -3 -3 3 3
use M3_M2  M3_M2_908
timestamp 1677677812
transform 1 0 3348 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_811
timestamp 1677677812
transform 1 0 3364 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_812
timestamp 1677677812
transform 1 0 3388 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_855
timestamp 1677677812
transform 1 0 3372 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1006
timestamp 1677677812
transform 1 0 3388 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1677677812
transform 1 0 3364 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1114
timestamp 1677677812
transform 1 0 3372 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1677677812
transform 1 0 3420 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_767
timestamp 1677677812
transform 1 0 3452 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_1007
timestamp 1677677812
transform 1 0 3452 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1677677812
transform 1 0 3468 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_813
timestamp 1677677812
transform 1 0 3484 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1009
timestamp 1677677812
transform 1 0 3484 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1116
timestamp 1677677812
transform 1 0 3436 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1677677812
transform 1 0 3444 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1677677812
transform 1 0 3460 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1677677812
transform 1 0 3476 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_909
timestamp 1677677812
transform 1 0 3444 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_910
timestamp 1677677812
transform 1 0 3476 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1120
timestamp 1677677812
transform 1 0 3500 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_814
timestamp 1677677812
transform 1 0 3516 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1677677812
transform 1 0 3540 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_1121
timestamp 1677677812
transform 1 0 3532 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_930
timestamp 1677677812
transform 1 0 3532 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_931
timestamp 1677677812
transform 1 0 3548 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_762
timestamp 1677677812
transform 1 0 3596 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_769
timestamp 1677677812
transform 1 0 3628 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_815
timestamp 1677677812
transform 1 0 3620 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1010
timestamp 1677677812
transform 1 0 3588 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_856
timestamp 1677677812
transform 1 0 3596 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1677677812
transform 1 0 3620 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1122
timestamp 1677677812
transform 1 0 3596 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1677677812
transform 1 0 3612 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1677677812
transform 1 0 3636 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1154
timestamp 1677677812
transform 1 0 3636 0 1 4185
box -2 -2 2 2
use M3_M2  M3_M2_816
timestamp 1677677812
transform 1 0 3644 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_817
timestamp 1677677812
transform 1 0 3660 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1124
timestamp 1677677812
transform 1 0 3652 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1013
timestamp 1677677812
transform 1 0 3668 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_911
timestamp 1677677812
transform 1 0 3676 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_749
timestamp 1677677812
transform 1 0 3740 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1677677812
transform 1 0 3732 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1014
timestamp 1677677812
transform 1 0 3732 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_871
timestamp 1677677812
transform 1 0 3716 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1125
timestamp 1677677812
transform 1 0 3780 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_770
timestamp 1677677812
transform 1 0 3868 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_819
timestamp 1677677812
transform 1 0 3836 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_820
timestamp 1677677812
transform 1 0 3860 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1015
timestamp 1677677812
transform 1 0 3828 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1016
timestamp 1677677812
transform 1 0 3844 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1126
timestamp 1677677812
transform 1 0 3836 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_912
timestamp 1677677812
transform 1 0 3828 0 1 4195
box -3 -3 3 3
use M2_M1  M2_M1_1127
timestamp 1677677812
transform 1 0 3868 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_913
timestamp 1677677812
transform 1 0 3868 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_932
timestamp 1677677812
transform 1 0 3868 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1017
timestamp 1677677812
transform 1 0 3884 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_872
timestamp 1677677812
transform 1 0 3884 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1677677812
transform 1 0 3908 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_771
timestamp 1677677812
transform 1 0 3924 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_821
timestamp 1677677812
transform 1 0 3916 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1018
timestamp 1677677812
transform 1 0 3908 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1019
timestamp 1677677812
transform 1 0 3924 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1677677812
transform 1 0 3900 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1129
timestamp 1677677812
transform 1 0 3916 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_873
timestamp 1677677812
transform 1 0 3924 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1020
timestamp 1677677812
transform 1 0 3956 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1677677812
transform 1 0 3956 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_822
timestamp 1677677812
transform 1 0 3996 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1021
timestamp 1677677812
transform 1 0 3996 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_857
timestamp 1677677812
transform 1 0 4044 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1131
timestamp 1677677812
transform 1 0 4044 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_751
timestamp 1677677812
transform 1 0 4116 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_823
timestamp 1677677812
transform 1 0 4124 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_858
timestamp 1677677812
transform 1 0 4116 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1022
timestamp 1677677812
transform 1 0 4124 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_859
timestamp 1677677812
transform 1 0 4148 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1677677812
transform 1 0 4084 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_763
timestamp 1677677812
transform 1 0 4204 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_824
timestamp 1677677812
transform 1 0 4220 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1023
timestamp 1677677812
transform 1 0 4196 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_860
timestamp 1677677812
transform 1 0 4204 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1024
timestamp 1677677812
transform 1 0 4212 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1025
timestamp 1677677812
transform 1 0 4228 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_874
timestamp 1677677812
transform 1 0 4196 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1133
timestamp 1677677812
transform 1 0 4204 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1677677812
transform 1 0 4220 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_875
timestamp 1677677812
transform 1 0 4228 0 1 4205
box -3 -3 3 3
use M2_M1  M2_M1_1135
timestamp 1677677812
transform 1 0 4236 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1677677812
transform 1 0 4252 0 1 4225
box -2 -2 2 2
use M3_M2  M3_M2_772
timestamp 1677677812
transform 1 0 4276 0 1 4245
box -3 -3 3 3
use M2_M1  M2_M1_916
timestamp 1677677812
transform 1 0 4268 0 1 4235
box -2 -2 2 2
use M3_M2  M3_M2_825
timestamp 1677677812
transform 1 0 4268 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1026
timestamp 1677677812
transform 1 0 4276 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1677677812
transform 1 0 4292 0 1 4225
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1677677812
transform 1 0 4316 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1028
timestamp 1677677812
transform 1 0 4332 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1136
timestamp 1677677812
transform 1 0 4300 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1137
timestamp 1677677812
transform 1 0 4308 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_876
timestamp 1677677812
transform 1 0 4316 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_933
timestamp 1677677812
transform 1 0 4300 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1677677812
transform 1 0 4372 0 1 4255
box -3 -3 3 3
use M3_M2  M3_M2_785
timestamp 1677677812
transform 1 0 4364 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_826
timestamp 1677677812
transform 1 0 4356 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1029
timestamp 1677677812
transform 1 0 4348 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_827
timestamp 1677677812
transform 1 0 4388 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_861
timestamp 1677677812
transform 1 0 4364 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1030
timestamp 1677677812
transform 1 0 4388 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1138
timestamp 1677677812
transform 1 0 4356 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1139
timestamp 1677677812
transform 1 0 4364 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1140
timestamp 1677677812
transform 1 0 4380 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1141
timestamp 1677677812
transform 1 0 4396 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_914
timestamp 1677677812
transform 1 0 4380 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_752
timestamp 1677677812
transform 1 0 4428 0 1 4265
box -3 -3 3 3
use M3_M2  M3_M2_765
timestamp 1677677812
transform 1 0 4420 0 1 4255
box -3 -3 3 3
use M2_M1  M2_M1_1031
timestamp 1677677812
transform 1 0 4452 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1677677812
transform 1 0 4428 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_915
timestamp 1677677812
transform 1 0 4452 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_934
timestamp 1677677812
transform 1 0 4468 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_828
timestamp 1677677812
transform 1 0 4524 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1032
timestamp 1677677812
transform 1 0 4524 0 1 4215
box -2 -2 2 2
use M3_M2  M3_M2_786
timestamp 1677677812
transform 1 0 4540 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1677677812
transform 1 0 4564 0 1 4245
box -3 -3 3 3
use M3_M2  M3_M2_829
timestamp 1677677812
transform 1 0 4572 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1033
timestamp 1677677812
transform 1 0 4556 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1677677812
transform 1 0 4572 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1035
timestamp 1677677812
transform 1 0 4596 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1143
timestamp 1677677812
transform 1 0 4564 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1144
timestamp 1677677812
transform 1 0 4580 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1145
timestamp 1677677812
transform 1 0 4588 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_916
timestamp 1677677812
transform 1 0 4564 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1677677812
transform 1 0 4708 0 1 4235
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1677677812
transform 1 0 4644 0 1 4225
box -3 -3 3 3
use M3_M2  M3_M2_831
timestamp 1677677812
transform 1 0 4700 0 1 4225
box -3 -3 3 3
use M2_M1  M2_M1_1036
timestamp 1677677812
transform 1 0 4644 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1677677812
transform 1 0 4700 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1677677812
transform 1 0 4716 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1677677812
transform 1 0 4732 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1146
timestamp 1677677812
transform 1 0 4620 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_877
timestamp 1677677812
transform 1 0 4700 0 1 4205
box -3 -3 3 3
use M3_M2  M3_M2_862
timestamp 1677677812
transform 1 0 4740 0 1 4215
box -3 -3 3 3
use M2_M1  M2_M1_1040
timestamp 1677677812
transform 1 0 4748 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1041
timestamp 1677677812
transform 1 0 4764 0 1 4215
box -2 -2 2 2
use M2_M1  M2_M1_1147
timestamp 1677677812
transform 1 0 4708 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1677677812
transform 1 0 4724 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1149
timestamp 1677677812
transform 1 0 4740 0 1 4205
box -2 -2 2 2
use M2_M1  M2_M1_1150
timestamp 1677677812
transform 1 0 4756 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_935
timestamp 1677677812
transform 1 0 4620 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_936
timestamp 1677677812
transform 1 0 4668 0 1 4185
box -3 -3 3 3
use M3_M2  M3_M2_917
timestamp 1677677812
transform 1 0 4764 0 1 4195
box -3 -3 3 3
use M3_M2  M3_M2_937
timestamp 1677677812
transform 1 0 4740 0 1 4185
box -3 -3 3 3
use M2_M1  M2_M1_1151
timestamp 1677677812
transform 1 0 4780 0 1 4205
box -2 -2 2 2
use M3_M2  M3_M2_938
timestamp 1677677812
transform 1 0 4772 0 1 4185
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_10
timestamp 1677677812
transform 1 0 48 0 1 4170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_69
timestamp 1677677812
transform 1 0 72 0 1 4170
box -8 -3 104 105
use FILL  FILL_812
timestamp 1677677812
transform 1 0 168 0 1 4170
box -8 -3 16 105
use FILL  FILL_813
timestamp 1677677812
transform 1 0 176 0 1 4170
box -8 -3 16 105
use FILL  FILL_814
timestamp 1677677812
transform 1 0 184 0 1 4170
box -8 -3 16 105
use FILL  FILL_815
timestamp 1677677812
transform 1 0 192 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_939
timestamp 1677677812
transform 1 0 212 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_80
timestamp 1677677812
transform -1 0 216 0 1 4170
box -9 -3 26 105
use FILL  FILL_816
timestamp 1677677812
transform 1 0 216 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_43
timestamp 1677677812
transform 1 0 224 0 1 4170
box -8 -3 46 105
use FILL  FILL_827
timestamp 1677677812
transform 1 0 264 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_70
timestamp 1677677812
transform 1 0 272 0 1 4170
box -8 -3 104 105
use M3_M2  M3_M2_940
timestamp 1677677812
transform 1 0 388 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_83
timestamp 1677677812
transform -1 0 384 0 1 4170
box -9 -3 26 105
use FILL  FILL_828
timestamp 1677677812
transform 1 0 384 0 1 4170
box -8 -3 16 105
use FILL  FILL_829
timestamp 1677677812
transform 1 0 392 0 1 4170
box -8 -3 16 105
use FILL  FILL_830
timestamp 1677677812
transform 1 0 400 0 1 4170
box -8 -3 16 105
use FILL  FILL_831
timestamp 1677677812
transform 1 0 408 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_44
timestamp 1677677812
transform 1 0 416 0 1 4170
box -8 -3 46 105
use FILL  FILL_832
timestamp 1677677812
transform 1 0 456 0 1 4170
box -8 -3 16 105
use FILL  FILL_833
timestamp 1677677812
transform 1 0 464 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_71
timestamp 1677677812
transform 1 0 472 0 1 4170
box -8 -3 104 105
use FILL  FILL_834
timestamp 1677677812
transform 1 0 568 0 1 4170
box -8 -3 16 105
use FILL  FILL_847
timestamp 1677677812
transform 1 0 576 0 1 4170
box -8 -3 16 105
use FILL  FILL_849
timestamp 1677677812
transform 1 0 584 0 1 4170
box -8 -3 16 105
use FILL  FILL_851
timestamp 1677677812
transform 1 0 592 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_46
timestamp 1677677812
transform 1 0 600 0 1 4170
box -8 -3 46 105
use FILL  FILL_852
timestamp 1677677812
transform 1 0 640 0 1 4170
box -8 -3 16 105
use FILL  FILL_855
timestamp 1677677812
transform 1 0 648 0 1 4170
box -8 -3 16 105
use FILL  FILL_857
timestamp 1677677812
transform 1 0 656 0 1 4170
box -8 -3 16 105
use FILL  FILL_859
timestamp 1677677812
transform 1 0 664 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_42
timestamp 1677677812
transform 1 0 672 0 1 4170
box -8 -3 46 105
use FILL  FILL_860
timestamp 1677677812
transform 1 0 712 0 1 4170
box -8 -3 16 105
use FILL  FILL_863
timestamp 1677677812
transform 1 0 720 0 1 4170
box -8 -3 16 105
use FILL  FILL_865
timestamp 1677677812
transform 1 0 728 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_73
timestamp 1677677812
transform -1 0 832 0 1 4170
box -8 -3 104 105
use FILL  FILL_867
timestamp 1677677812
transform 1 0 832 0 1 4170
box -8 -3 16 105
use FILL  FILL_869
timestamp 1677677812
transform 1 0 840 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_941
timestamp 1677677812
transform 1 0 900 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_75
timestamp 1677677812
transform 1 0 848 0 1 4170
box -8 -3 104 105
use FILL  FILL_871
timestamp 1677677812
transform 1 0 944 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_89
timestamp 1677677812
transform 1 0 952 0 1 4170
box -9 -3 26 105
use FILL  FILL_877
timestamp 1677677812
transform 1 0 968 0 1 4170
box -8 -3 16 105
use FILL  FILL_881
timestamp 1677677812
transform 1 0 976 0 1 4170
box -8 -3 16 105
use FILL  FILL_883
timestamp 1677677812
transform 1 0 984 0 1 4170
box -8 -3 16 105
use FILL  FILL_884
timestamp 1677677812
transform 1 0 992 0 1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_12
timestamp 1677677812
transform 1 0 1000 0 1 4170
box -8 -3 32 105
use FILL  FILL_885
timestamp 1677677812
transform 1 0 1024 0 1 4170
box -8 -3 16 105
use FILL  FILL_888
timestamp 1677677812
transform 1 0 1032 0 1 4170
box -8 -3 16 105
use FILL  FILL_890
timestamp 1677677812
transform 1 0 1040 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_25
timestamp 1677677812
transform 1 0 1048 0 1 4170
box -8 -3 34 105
use FILL  FILL_892
timestamp 1677677812
transform 1 0 1080 0 1 4170
box -8 -3 16 105
use FILL  FILL_895
timestamp 1677677812
transform 1 0 1088 0 1 4170
box -8 -3 16 105
use FILL  FILL_897
timestamp 1677677812
transform 1 0 1096 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_49
timestamp 1677677812
transform 1 0 1104 0 1 4170
box -8 -3 46 105
use FILL  FILL_899
timestamp 1677677812
transform 1 0 1144 0 1 4170
box -8 -3 16 105
use FILL  FILL_902
timestamp 1677677812
transform 1 0 1152 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_90
timestamp 1677677812
transform 1 0 1160 0 1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_76
timestamp 1677677812
transform -1 0 1272 0 1 4170
box -8 -3 104 105
use OAI21X1  OAI21X1_27
timestamp 1677677812
transform -1 0 1304 0 1 4170
box -8 -3 34 105
use FILL  FILL_904
timestamp 1677677812
transform 1 0 1304 0 1 4170
box -8 -3 16 105
use FILL  FILL_905
timestamp 1677677812
transform 1 0 1312 0 1 4170
box -8 -3 16 105
use FILL  FILL_906
timestamp 1677677812
transform 1 0 1320 0 1 4170
box -8 -3 16 105
use FILL  FILL_907
timestamp 1677677812
transform 1 0 1328 0 1 4170
box -8 -3 16 105
use FILL  FILL_908
timestamp 1677677812
transform 1 0 1336 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_77
timestamp 1677677812
transform -1 0 1440 0 1 4170
box -8 -3 104 105
use FILL  FILL_909
timestamp 1677677812
transform 1 0 1440 0 1 4170
box -8 -3 16 105
use FILL  FILL_910
timestamp 1677677812
transform 1 0 1448 0 1 4170
box -8 -3 16 105
use FILL  FILL_911
timestamp 1677677812
transform 1 0 1456 0 1 4170
box -8 -3 16 105
use FILL  FILL_925
timestamp 1677677812
transform 1 0 1464 0 1 4170
box -8 -3 16 105
use FILL  FILL_927
timestamp 1677677812
transform 1 0 1472 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_93
timestamp 1677677812
transform -1 0 1496 0 1 4170
box -9 -3 26 105
use FILL  FILL_928
timestamp 1677677812
transform 1 0 1496 0 1 4170
box -8 -3 16 105
use FILL  FILL_929
timestamp 1677677812
transform 1 0 1504 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_45
timestamp 1677677812
transform -1 0 1552 0 1 4170
box -8 -3 46 105
use FILL  FILL_930
timestamp 1677677812
transform 1 0 1552 0 1 4170
box -8 -3 16 105
use FILL  FILL_931
timestamp 1677677812
transform 1 0 1560 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_94
timestamp 1677677812
transform -1 0 1584 0 1 4170
box -9 -3 26 105
use FILL  FILL_932
timestamp 1677677812
transform 1 0 1584 0 1 4170
box -8 -3 16 105
use FILL  FILL_936
timestamp 1677677812
transform 1 0 1592 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_95
timestamp 1677677812
transform 1 0 1600 0 1 4170
box -9 -3 26 105
use FILL  FILL_938
timestamp 1677677812
transform 1 0 1616 0 1 4170
box -8 -3 16 105
use FILL  FILL_939
timestamp 1677677812
transform 1 0 1624 0 1 4170
box -8 -3 16 105
use FILL  FILL_940
timestamp 1677677812
transform 1 0 1632 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_96
timestamp 1677677812
transform -1 0 1656 0 1 4170
box -9 -3 26 105
use M3_M2  M3_M2_942
timestamp 1677677812
transform 1 0 1684 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_97
timestamp 1677677812
transform 1 0 1656 0 1 4170
box -9 -3 26 105
use FILL  FILL_941
timestamp 1677677812
transform 1 0 1672 0 1 4170
box -8 -3 16 105
use FILL  FILL_947
timestamp 1677677812
transform 1 0 1680 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_98
timestamp 1677677812
transform 1 0 1688 0 1 4170
box -9 -3 26 105
use FILL  FILL_949
timestamp 1677677812
transform 1 0 1704 0 1 4170
box -8 -3 16 105
use FILL  FILL_950
timestamp 1677677812
transform 1 0 1712 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_943
timestamp 1677677812
transform 1 0 1812 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_80
timestamp 1677677812
transform 1 0 1720 0 1 4170
box -8 -3 104 105
use FILL  FILL_951
timestamp 1677677812
transform 1 0 1816 0 1 4170
box -8 -3 16 105
use FILL  FILL_955
timestamp 1677677812
transform 1 0 1824 0 1 4170
box -8 -3 16 105
use FILL  FILL_957
timestamp 1677677812
transform 1 0 1832 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_50
timestamp 1677677812
transform 1 0 1840 0 1 4170
box -8 -3 46 105
use FILL  FILL_959
timestamp 1677677812
transform 1 0 1880 0 1 4170
box -8 -3 16 105
use FILL  FILL_960
timestamp 1677677812
transform 1 0 1888 0 1 4170
box -8 -3 16 105
use FILL  FILL_961
timestamp 1677677812
transform 1 0 1896 0 1 4170
box -8 -3 16 105
use FILL  FILL_965
timestamp 1677677812
transform 1 0 1904 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_100
timestamp 1677677812
transform -1 0 1928 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_101
timestamp 1677677812
transform 1 0 1928 0 1 4170
box -9 -3 26 105
use FILL  FILL_966
timestamp 1677677812
transform 1 0 1944 0 1 4170
box -8 -3 16 105
use FILL  FILL_973
timestamp 1677677812
transform 1 0 1952 0 1 4170
box -8 -3 16 105
use FILL  FILL_975
timestamp 1677677812
transform 1 0 1960 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_52
timestamp 1677677812
transform 1 0 1968 0 1 4170
box -8 -3 46 105
use FILL  FILL_976
timestamp 1677677812
transform 1 0 2008 0 1 4170
box -8 -3 16 105
use FILL  FILL_979
timestamp 1677677812
transform 1 0 2016 0 1 4170
box -8 -3 16 105
use FILL  FILL_981
timestamp 1677677812
transform 1 0 2024 0 1 4170
box -8 -3 16 105
use FILL  FILL_982
timestamp 1677677812
transform 1 0 2032 0 1 4170
box -8 -3 16 105
use FILL  FILL_983
timestamp 1677677812
transform 1 0 2040 0 1 4170
box -8 -3 16 105
use FILL  FILL_984
timestamp 1677677812
transform 1 0 2048 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_944
timestamp 1677677812
transform 1 0 2068 0 1 4175
box -3 -3 3 3
use FILL  FILL_985
timestamp 1677677812
transform 1 0 2056 0 1 4170
box -8 -3 16 105
use FILL  FILL_986
timestamp 1677677812
transform 1 0 2064 0 1 4170
box -8 -3 16 105
use FILL  FILL_987
timestamp 1677677812
transform 1 0 2072 0 1 4170
box -8 -3 16 105
use FILL  FILL_990
timestamp 1677677812
transform 1 0 2080 0 1 4170
box -8 -3 16 105
use FILL  FILL_992
timestamp 1677677812
transform 1 0 2088 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_102
timestamp 1677677812
transform 1 0 2096 0 1 4170
box -9 -3 26 105
use FILL  FILL_994
timestamp 1677677812
transform 1 0 2112 0 1 4170
box -8 -3 16 105
use FILL  FILL_998
timestamp 1677677812
transform 1 0 2120 0 1 4170
box -8 -3 16 105
use FILL  FILL_999
timestamp 1677677812
transform 1 0 2128 0 1 4170
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1677677812
transform 1 0 2136 0 1 4170
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1677677812
transform 1 0 2144 0 1 4170
box -8 -3 16 105
use FILL  FILL_1002
timestamp 1677677812
transform 1 0 2152 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_103
timestamp 1677677812
transform 1 0 2160 0 1 4170
box -9 -3 26 105
use FILL  FILL_1003
timestamp 1677677812
transform 1 0 2176 0 1 4170
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1677677812
transform 1 0 2184 0 1 4170
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1677677812
transform 1 0 2192 0 1 4170
box -8 -3 16 105
use FILL  FILL_1006
timestamp 1677677812
transform 1 0 2200 0 1 4170
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1677677812
transform 1 0 2208 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_82
timestamp 1677677812
transform 1 0 2216 0 1 4170
box -8 -3 104 105
use FILL  FILL_1008
timestamp 1677677812
transform 1 0 2312 0 1 4170
box -8 -3 16 105
use FILL  FILL_1022
timestamp 1677677812
transform 1 0 2320 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_48
timestamp 1677677812
transform 1 0 2328 0 1 4170
box -8 -3 46 105
use FILL  FILL_1024
timestamp 1677677812
transform 1 0 2368 0 1 4170
box -8 -3 16 105
use FILL  FILL_1031
timestamp 1677677812
transform 1 0 2376 0 1 4170
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1677677812
transform 1 0 2384 0 1 4170
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1677677812
transform 1 0 2392 0 1 4170
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1677677812
transform 1 0 2400 0 1 4170
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1677677812
transform 1 0 2408 0 1 4170
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1677677812
transform 1 0 2416 0 1 4170
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1677677812
transform 1 0 2424 0 1 4170
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1677677812
transform 1 0 2432 0 1 4170
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1677677812
transform 1 0 2440 0 1 4170
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1677677812
transform 1 0 2448 0 1 4170
box -8 -3 16 105
use FILL  FILL_1046
timestamp 1677677812
transform 1 0 2456 0 1 4170
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1677677812
transform 1 0 2464 0 1 4170
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1677677812
transform 1 0 2472 0 1 4170
box -8 -3 16 105
use FILL  FILL_1051
timestamp 1677677812
transform 1 0 2480 0 1 4170
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1677677812
transform 1 0 2488 0 1 4170
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1677677812
transform 1 0 2496 0 1 4170
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1677677812
transform 1 0 2504 0 1 4170
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1677677812
transform 1 0 2512 0 1 4170
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1677677812
transform 1 0 2520 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_945
timestamp 1677677812
transform 1 0 2540 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_946
timestamp 1677677812
transform 1 0 2580 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_947
timestamp 1677677812
transform 1 0 2612 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_84
timestamp 1677677812
transform 1 0 2528 0 1 4170
box -8 -3 104 105
use M3_M2  M3_M2_948
timestamp 1677677812
transform 1 0 2636 0 1 4175
box -3 -3 3 3
use FILL  FILL_1061
timestamp 1677677812
transform 1 0 2624 0 1 4170
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1677677812
transform 1 0 2632 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_54
timestamp 1677677812
transform 1 0 2640 0 1 4170
box -8 -3 46 105
use FILL  FILL_1063
timestamp 1677677812
transform 1 0 2680 0 1 4170
box -8 -3 16 105
use FILL  FILL_1064
timestamp 1677677812
transform 1 0 2688 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_105
timestamp 1677677812
transform 1 0 2696 0 1 4170
box -9 -3 26 105
use FILL  FILL_1065
timestamp 1677677812
transform 1 0 2712 0 1 4170
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1677677812
transform 1 0 2720 0 1 4170
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1677677812
transform 1 0 2728 0 1 4170
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1677677812
transform 1 0 2736 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_86
timestamp 1677677812
transform 1 0 2744 0 1 4170
box -8 -3 104 105
use OAI21X1  OAI21X1_29
timestamp 1677677812
transform 1 0 2840 0 1 4170
box -8 -3 34 105
use FILL  FILL_1078
timestamp 1677677812
transform 1 0 2872 0 1 4170
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1677677812
transform 1 0 2880 0 1 4170
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1677677812
transform 1 0 2888 0 1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_30
timestamp 1677677812
transform 1 0 2896 0 1 4170
box -8 -3 34 105
use FILL  FILL_1094
timestamp 1677677812
transform 1 0 2928 0 1 4170
box -8 -3 16 105
use FILL  FILL_1095
timestamp 1677677812
transform 1 0 2936 0 1 4170
box -8 -3 16 105
use FILL  FILL_1096
timestamp 1677677812
transform 1 0 2944 0 1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_16
timestamp 1677677812
transform 1 0 2952 0 1 4170
box -8 -3 32 105
use FILL  FILL_1097
timestamp 1677677812
transform 1 0 2976 0 1 4170
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1677677812
transform 1 0 2984 0 1 4170
box -8 -3 16 105
use FILL  FILL_1106
timestamp 1677677812
transform 1 0 2992 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_949
timestamp 1677677812
transform 1 0 3012 0 1 4175
box -3 -3 3 3
use FILL  FILL_1107
timestamp 1677677812
transform 1 0 3000 0 1 4170
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1677677812
transform 1 0 3008 0 1 4170
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1677677812
transform 1 0 3016 0 1 4170
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1677677812
transform 1 0 3024 0 1 4170
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1677677812
transform 1 0 3032 0 1 4170
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1677677812
transform 1 0 3040 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_950
timestamp 1677677812
transform 1 0 3068 0 1 4175
box -3 -3 3 3
use OAI21X1  OAI21X1_33
timestamp 1677677812
transform -1 0 3080 0 1 4170
box -8 -3 34 105
use FILL  FILL_1116
timestamp 1677677812
transform 1 0 3080 0 1 4170
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1677677812
transform 1 0 3088 0 1 4170
box -8 -3 16 105
use FILL  FILL_1120
timestamp 1677677812
transform 1 0 3096 0 1 4170
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1677677812
transform 1 0 3104 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_951
timestamp 1677677812
transform 1 0 3156 0 1 4175
box -3 -3 3 3
use OAI22X1  OAI22X1_51
timestamp 1677677812
transform -1 0 3152 0 1 4170
box -8 -3 46 105
use FILL  FILL_1123
timestamp 1677677812
transform 1 0 3152 0 1 4170
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1677677812
transform 1 0 3160 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_952
timestamp 1677677812
transform 1 0 3196 0 1 4175
box -3 -3 3 3
use INVX2  INVX2_107
timestamp 1677677812
transform 1 0 3168 0 1 4170
box -9 -3 26 105
use FILL  FILL_1125
timestamp 1677677812
transform 1 0 3184 0 1 4170
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1677677812
transform 1 0 3192 0 1 4170
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1677677812
transform 1 0 3200 0 1 4170
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1677677812
transform 1 0 3208 0 1 4170
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1677677812
transform 1 0 3216 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_53
timestamp 1677677812
transform -1 0 3264 0 1 4170
box -8 -3 46 105
use FILL  FILL_1137
timestamp 1677677812
transform 1 0 3264 0 1 4170
box -8 -3 16 105
use FILL  FILL_1138
timestamp 1677677812
transform 1 0 3272 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_109
timestamp 1677677812
transform -1 0 3296 0 1 4170
box -9 -3 26 105
use FILL  FILL_1139
timestamp 1677677812
transform 1 0 3296 0 1 4170
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1677677812
transform 1 0 3304 0 1 4170
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1677677812
transform 1 0 3312 0 1 4170
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1677677812
transform 1 0 3320 0 1 4170
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1677677812
transform 1 0 3328 0 1 4170
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1677677812
transform 1 0 3336 0 1 4170
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1677677812
transform 1 0 3344 0 1 4170
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1677677812
transform 1 0 3352 0 1 4170
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1677677812
transform 1 0 3360 0 1 4170
box -8 -3 16 105
use BUFX2  BUFX2_0
timestamp 1677677812
transform -1 0 3392 0 1 4170
box -5 -3 28 105
use BUFX2  BUFX2_1
timestamp 1677677812
transform 1 0 3392 0 1 4170
box -5 -3 28 105
use FILL  FILL_1152
timestamp 1677677812
transform 1 0 3416 0 1 4170
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1677677812
transform 1 0 3424 0 1 4170
box -8 -3 16 105
use FILL  FILL_1160
timestamp 1677677812
transform 1 0 3432 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_54
timestamp 1677677812
transform 1 0 3440 0 1 4170
box -8 -3 46 105
use FILL  FILL_1162
timestamp 1677677812
transform 1 0 3480 0 1 4170
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1677677812
transform 1 0 3488 0 1 4170
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1677677812
transform 1 0 3496 0 1 4170
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1677677812
transform 1 0 3504 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_111
timestamp 1677677812
transform 1 0 3512 0 1 4170
box -9 -3 26 105
use FILL  FILL_1170
timestamp 1677677812
transform 1 0 3528 0 1 4170
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1677677812
transform 1 0 3536 0 1 4170
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1677677812
transform 1 0 3544 0 1 4170
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1677677812
transform 1 0 3552 0 1 4170
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1677677812
transform 1 0 3560 0 1 4170
box -8 -3 16 105
use FILL  FILL_1179
timestamp 1677677812
transform 1 0 3568 0 1 4170
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1677677812
transform 1 0 3576 0 1 4170
box -8 -3 16 105
use FILL  FILL_1181
timestamp 1677677812
transform 1 0 3584 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_55
timestamp 1677677812
transform 1 0 3592 0 1 4170
box -8 -3 46 105
use FILL  FILL_1184
timestamp 1677677812
transform 1 0 3632 0 1 4170
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1677677812
transform 1 0 3640 0 1 4170
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1677677812
transform 1 0 3648 0 1 4170
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1677677812
transform 1 0 3656 0 1 4170
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1677677812
transform 1 0 3664 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_112
timestamp 1677677812
transform -1 0 3688 0 1 4170
box -9 -3 26 105
use FILL  FILL_1192
timestamp 1677677812
transform 1 0 3688 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_88
timestamp 1677677812
transform -1 0 3792 0 1 4170
box -8 -3 104 105
use FILL  FILL_1193
timestamp 1677677812
transform 1 0 3792 0 1 4170
box -8 -3 16 105
use FILL  FILL_1198
timestamp 1677677812
transform 1 0 3800 0 1 4170
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1677677812
transform 1 0 3808 0 1 4170
box -8 -3 16 105
use FILL  FILL_1201
timestamp 1677677812
transform 1 0 3816 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_58
timestamp 1677677812
transform -1 0 3864 0 1 4170
box -8 -3 46 105
use FILL  FILL_1202
timestamp 1677677812
transform 1 0 3864 0 1 4170
box -8 -3 16 105
use FILL  FILL_1206
timestamp 1677677812
transform 1 0 3872 0 1 4170
box -8 -3 16 105
use FILL  FILL_1208
timestamp 1677677812
transform 1 0 3880 0 1 4170
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1677677812
transform 1 0 3888 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_57
timestamp 1677677812
transform 1 0 3896 0 1 4170
box -8 -3 46 105
use FILL  FILL_1210
timestamp 1677677812
transform 1 0 3936 0 1 4170
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1677677812
transform 1 0 3944 0 1 4170
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1677677812
transform 1 0 3952 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_90
timestamp 1677677812
transform -1 0 4056 0 1 4170
box -8 -3 104 105
use FILL  FILL_1217
timestamp 1677677812
transform 1 0 4056 0 1 4170
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1677677812
transform 1 0 4064 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_91
timestamp 1677677812
transform 1 0 4072 0 1 4170
box -8 -3 104 105
use FILL  FILL_1219
timestamp 1677677812
transform 1 0 4168 0 1 4170
box -8 -3 16 105
use INVX2  INVX2_114
timestamp 1677677812
transform 1 0 4176 0 1 4170
box -9 -3 26 105
use FILL  FILL_1220
timestamp 1677677812
transform 1 0 4192 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_58
timestamp 1677677812
transform 1 0 4200 0 1 4170
box -8 -3 46 105
use FILL  FILL_1221
timestamp 1677677812
transform 1 0 4240 0 1 4170
box -8 -3 16 105
use FILL  FILL_1233
timestamp 1677677812
transform 1 0 4248 0 1 4170
box -8 -3 16 105
use NAND3X1  NAND3X1_5
timestamp 1677677812
transform -1 0 4288 0 1 4170
box -8 -3 40 105
use FILL  FILL_1235
timestamp 1677677812
transform 1 0 4288 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_60
timestamp 1677677812
transform -1 0 4336 0 1 4170
box -8 -3 46 105
use FILL  FILL_1237
timestamp 1677677812
transform 1 0 4336 0 1 4170
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1677677812
transform 1 0 4344 0 1 4170
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1677677812
transform 1 0 4352 0 1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_61
timestamp 1677677812
transform 1 0 4360 0 1 4170
box -8 -3 46 105
use FILL  FILL_1243
timestamp 1677677812
transform 1 0 4400 0 1 4170
box -8 -3 16 105
use FILL  FILL_1244
timestamp 1677677812
transform 1 0 4408 0 1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_93
timestamp 1677677812
transform 1 0 4416 0 1 4170
box -8 -3 104 105
use INVX2  INVX2_117
timestamp 1677677812
transform 1 0 4512 0 1 4170
box -9 -3 26 105
use FILL  FILL_1247
timestamp 1677677812
transform 1 0 4528 0 1 4170
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1677677812
transform 1 0 4536 0 1 4170
box -8 -3 16 105
use FILL  FILL_1253
timestamp 1677677812
transform 1 0 4544 0 1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_62
timestamp 1677677812
transform 1 0 4552 0 1 4170
box -8 -3 46 105
use FILL  FILL_1255
timestamp 1677677812
transform 1 0 4592 0 1 4170
box -8 -3 16 105
use FILL  FILL_1257
timestamp 1677677812
transform 1 0 4600 0 1 4170
box -8 -3 16 105
use M3_M2  M3_M2_953
timestamp 1677677812
transform 1 0 4708 0 1 4175
box -3 -3 3 3
use M3_M2  M3_M2_954
timestamp 1677677812
transform 1 0 4732 0 1 4175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_95
timestamp 1677677812
transform 1 0 4608 0 1 4170
box -8 -3 104 105
use OAI22X1  OAI22X1_63
timestamp 1677677812
transform 1 0 4704 0 1 4170
box -8 -3 46 105
use INVX2  INVX2_118
timestamp 1677677812
transform -1 0 4760 0 1 4170
box -9 -3 26 105
use INVX2  INVX2_119
timestamp 1677677812
transform -1 0 4776 0 1 4170
box -9 -3 26 105
use FILL  FILL_1259
timestamp 1677677812
transform 1 0 4776 0 1 4170
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1677677812
transform 1 0 4784 0 1 4170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_11
timestamp 1677677812
transform 1 0 4819 0 1 4170
box -10 -3 10 3
use M3_M2  M3_M2_1108
timestamp 1677677812
transform 1 0 84 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1271
timestamp 1677677812
transform 1 0 116 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1161
timestamp 1677677812
transform 1 0 164 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1677677812
transform 1 0 172 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1677677812
transform 1 0 188 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1272
timestamp 1677677812
transform 1 0 164 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1061
timestamp 1677677812
transform 1 0 172 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1273
timestamp 1677677812
transform 1 0 180 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1274
timestamp 1677677812
transform 1 0 196 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1275
timestamp 1677677812
transform 1 0 204 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1073
timestamp 1677677812
transform 1 0 164 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1074
timestamp 1677677812
transform 1 0 204 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1109
timestamp 1677677812
transform 1 0 180 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1164
timestamp 1677677812
transform 1 0 220 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1027
timestamp 1677677812
transform 1 0 228 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1276
timestamp 1677677812
transform 1 0 228 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_955
timestamp 1677677812
transform 1 0 284 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_981
timestamp 1677677812
transform 1 0 276 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1165
timestamp 1677677812
transform 1 0 252 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1166
timestamp 1677677812
transform 1 0 260 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1167
timestamp 1677677812
transform 1 0 276 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1168
timestamp 1677677812
transform 1 0 292 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1169
timestamp 1677677812
transform 1 0 300 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1277
timestamp 1677677812
transform 1 0 244 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1134
timestamp 1677677812
transform 1 0 236 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1062
timestamp 1677677812
transform 1 0 260 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1278
timestamp 1677677812
transform 1 0 268 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1279
timestamp 1677677812
transform 1 0 284 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1135
timestamp 1677677812
transform 1 0 284 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_956
timestamp 1677677812
transform 1 0 308 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1004
timestamp 1677677812
transform 1 0 404 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1170
timestamp 1677677812
transform 1 0 324 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1280
timestamp 1677677812
transform 1 0 308 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1281
timestamp 1677677812
transform 1 0 372 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1282
timestamp 1677677812
transform 1 0 404 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1283
timestamp 1677677812
transform 1 0 412 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1075
timestamp 1677677812
transform 1 0 372 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1076
timestamp 1677677812
transform 1 0 412 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1110
timestamp 1677677812
transform 1 0 404 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1005
timestamp 1677677812
transform 1 0 428 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1028
timestamp 1677677812
transform 1 0 436 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1284
timestamp 1677677812
transform 1 0 436 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1029
timestamp 1677677812
transform 1 0 452 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1171
timestamp 1677677812
transform 1 0 460 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1677677812
transform 1 0 468 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1173
timestamp 1677677812
transform 1 0 484 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1285
timestamp 1677677812
transform 1 0 476 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1063
timestamp 1677677812
transform 1 0 484 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_1111
timestamp 1677677812
transform 1 0 468 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1286
timestamp 1677677812
transform 1 0 500 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1287
timestamp 1677677812
transform 1 0 508 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1077
timestamp 1677677812
transform 1 0 500 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1174
timestamp 1677677812
transform 1 0 548 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1030
timestamp 1677677812
transform 1 0 556 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1136
timestamp 1677677812
transform 1 0 556 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1175
timestamp 1677677812
transform 1 0 572 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1288
timestamp 1677677812
transform 1 0 564 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1176
timestamp 1677677812
transform 1 0 588 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1289
timestamp 1677677812
transform 1 0 580 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1078
timestamp 1677677812
transform 1 0 580 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1006
timestamp 1677677812
transform 1 0 620 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1177
timestamp 1677677812
transform 1 0 604 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1031
timestamp 1677677812
transform 1 0 612 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1178
timestamp 1677677812
transform 1 0 620 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1064
timestamp 1677677812
transform 1 0 604 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1290
timestamp 1677677812
transform 1 0 612 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1291
timestamp 1677677812
transform 1 0 636 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1137
timestamp 1677677812
transform 1 0 636 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1179
timestamp 1677677812
transform 1 0 660 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1112
timestamp 1677677812
transform 1 0 660 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1007
timestamp 1677677812
transform 1 0 700 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1180
timestamp 1677677812
transform 1 0 684 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1032
timestamp 1677677812
transform 1 0 692 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1181
timestamp 1677677812
transform 1 0 700 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1292
timestamp 1677677812
transform 1 0 676 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1293
timestamp 1677677812
transform 1 0 692 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1079
timestamp 1677677812
transform 1 0 676 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1294
timestamp 1677677812
transform 1 0 732 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_957
timestamp 1677677812
transform 1 0 820 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1182
timestamp 1677677812
transform 1 0 820 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1295
timestamp 1677677812
transform 1 0 772 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1080
timestamp 1677677812
transform 1 0 748 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1138
timestamp 1677677812
transform 1 0 780 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_982
timestamp 1677677812
transform 1 0 836 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1157
timestamp 1677677812
transform 1 0 836 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1677677812
transform 1 0 868 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1139
timestamp 1677677812
transform 1 0 860 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1008
timestamp 1677677812
transform 1 0 892 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1296
timestamp 1677677812
transform 1 0 892 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1297
timestamp 1677677812
transform 1 0 900 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1677677812
transform 1 0 916 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1185
timestamp 1677677812
transform 1 0 932 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1298
timestamp 1677677812
transform 1 0 924 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_983
timestamp 1677677812
transform 1 0 964 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1299
timestamp 1677677812
transform 1 0 964 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1300
timestamp 1677677812
transform 1 0 972 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1009
timestamp 1677677812
transform 1 0 1020 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1158
timestamp 1677677812
transform 1 0 1028 0 1 4145
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1677677812
transform 1 0 1020 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1033
timestamp 1677677812
transform 1 0 1028 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1385
timestamp 1677677812
transform 1 0 1036 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1187
timestamp 1677677812
transform 1 0 1052 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_984
timestamp 1677677812
transform 1 0 1100 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1188
timestamp 1677677812
transform 1 0 1084 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1189
timestamp 1677677812
transform 1 0 1092 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1301
timestamp 1677677812
transform 1 0 1076 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1148
timestamp 1677677812
transform 1 0 1076 0 1 4085
box -3 -3 3 3
use M2_M1  M2_M1_1190
timestamp 1677677812
transform 1 0 1132 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1677677812
transform 1 0 1148 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1010
timestamp 1677677812
transform 1 0 1164 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1386
timestamp 1677677812
transform 1 0 1164 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1034
timestamp 1677677812
transform 1 0 1180 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1035
timestamp 1677677812
transform 1 0 1220 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1192
timestamp 1677677812
transform 1 0 1268 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1302
timestamp 1677677812
transform 1 0 1180 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1303
timestamp 1677677812
transform 1 0 1188 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1304
timestamp 1677677812
transform 1 0 1220 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1011
timestamp 1677677812
transform 1 0 1284 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1193
timestamp 1677677812
transform 1 0 1284 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1036
timestamp 1677677812
transform 1 0 1292 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1387
timestamp 1677677812
transform 1 0 1292 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1388
timestamp 1677677812
transform 1 0 1308 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_985
timestamp 1677677812
transform 1 0 1340 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1037
timestamp 1677677812
transform 1 0 1332 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1194
timestamp 1677677812
transform 1 0 1340 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1677677812
transform 1 0 1348 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1305
timestamp 1677677812
transform 1 0 1332 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1306
timestamp 1677677812
transform 1 0 1340 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_958
timestamp 1677677812
transform 1 0 1380 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_959
timestamp 1677677812
transform 1 0 1404 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1038
timestamp 1677677812
transform 1 0 1396 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1196
timestamp 1677677812
transform 1 0 1404 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1307
timestamp 1677677812
transform 1 0 1412 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1039
timestamp 1677677812
transform 1 0 1428 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1197
timestamp 1677677812
transform 1 0 1436 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_960
timestamp 1677677812
transform 1 0 1460 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1040
timestamp 1677677812
transform 1 0 1460 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1198
timestamp 1677677812
transform 1 0 1468 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1308
timestamp 1677677812
transform 1 0 1428 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1309
timestamp 1677677812
transform 1 0 1452 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1677677812
transform 1 0 1484 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_961
timestamp 1677677812
transform 1 0 1516 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_986
timestamp 1677677812
transform 1 0 1564 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1012
timestamp 1677677812
transform 1 0 1548 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1677677812
transform 1 0 1500 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1041
timestamp 1677677812
transform 1 0 1540 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_962
timestamp 1677677812
transform 1 0 1588 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1201
timestamp 1677677812
transform 1 0 1588 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1310
timestamp 1677677812
transform 1 0 1548 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1311
timestamp 1677677812
transform 1 0 1580 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1042
timestamp 1677677812
transform 1 0 1612 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_963
timestamp 1677677812
transform 1 0 1636 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_987
timestamp 1677677812
transform 1 0 1628 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1013
timestamp 1677677812
transform 1 0 1636 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1202
timestamp 1677677812
transform 1 0 1620 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1203
timestamp 1677677812
transform 1 0 1636 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1043
timestamp 1677677812
transform 1 0 1644 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1312
timestamp 1677677812
transform 1 0 1628 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1313
timestamp 1677677812
transform 1 0 1644 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1204
timestamp 1677677812
transform 1 0 1692 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1314
timestamp 1677677812
transform 1 0 1684 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_964
timestamp 1677677812
transform 1 0 1772 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1014
timestamp 1677677812
transform 1 0 1788 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1205
timestamp 1677677812
transform 1 0 1708 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1044
timestamp 1677677812
transform 1 0 1756 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1045
timestamp 1677677812
transform 1 0 1796 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1315
timestamp 1677677812
transform 1 0 1756 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1316
timestamp 1677677812
transform 1 0 1788 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1317
timestamp 1677677812
transform 1 0 1796 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_988
timestamp 1677677812
transform 1 0 1820 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1318
timestamp 1677677812
transform 1 0 1812 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_989
timestamp 1677677812
transform 1 0 1868 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1015
timestamp 1677677812
transform 1 0 1884 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1206
timestamp 1677677812
transform 1 0 1860 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1207
timestamp 1677677812
transform 1 0 1868 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1208
timestamp 1677677812
transform 1 0 1884 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1319
timestamp 1677677812
transform 1 0 1876 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1320
timestamp 1677677812
transform 1 0 1892 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1321
timestamp 1677677812
transform 1 0 1900 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1155
timestamp 1677677812
transform 1 0 1908 0 1 4155
box -2 -2 2 2
use M3_M2  M3_M2_1016
timestamp 1677677812
transform 1 0 1908 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_965
timestamp 1677677812
transform 1 0 1940 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1156
timestamp 1677677812
transform 1 0 1956 0 1 4155
box -2 -2 2 2
use M2_M1  M2_M1_1322
timestamp 1677677812
transform 1 0 1956 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_966
timestamp 1677677812
transform 1 0 1988 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1017
timestamp 1677677812
transform 1 0 1980 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1209
timestamp 1677677812
transform 1 0 1980 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1323
timestamp 1677677812
transform 1 0 1988 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1324
timestamp 1677677812
transform 1 0 2004 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_990
timestamp 1677677812
transform 1 0 2044 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_991
timestamp 1677677812
transform 1 0 2076 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1210
timestamp 1677677812
transform 1 0 2044 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1211
timestamp 1677677812
transform 1 0 2060 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1212
timestamp 1677677812
transform 1 0 2068 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1325
timestamp 1677677812
transform 1 0 2052 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1326
timestamp 1677677812
transform 1 0 2076 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1213
timestamp 1677677812
transform 1 0 2116 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1046
timestamp 1677677812
transform 1 0 2124 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1214
timestamp 1677677812
transform 1 0 2212 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1327
timestamp 1677677812
transform 1 0 2164 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_967
timestamp 1677677812
transform 1 0 2228 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1215
timestamp 1677677812
transform 1 0 2308 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1081
timestamp 1677677812
transform 1 0 2332 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1216
timestamp 1677677812
transform 1 0 2412 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1217
timestamp 1677677812
transform 1 0 2428 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1328
timestamp 1677677812
transform 1 0 2404 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1065
timestamp 1677677812
transform 1 0 2412 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1329
timestamp 1677677812
transform 1 0 2420 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1082
timestamp 1677677812
transform 1 0 2420 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1113
timestamp 1677677812
transform 1 0 2412 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1114
timestamp 1677677812
transform 1 0 2436 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1218
timestamp 1677677812
transform 1 0 2476 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1047
timestamp 1677677812
transform 1 0 2484 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1219
timestamp 1677677812
transform 1 0 2492 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1083
timestamp 1677677812
transform 1 0 2476 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1048
timestamp 1677677812
transform 1 0 2516 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1330
timestamp 1677677812
transform 1 0 2516 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1140
timestamp 1677677812
transform 1 0 2516 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1220
timestamp 1677677812
transform 1 0 2532 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1331
timestamp 1677677812
transform 1 0 2540 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1084
timestamp 1677677812
transform 1 0 2540 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1049
timestamp 1677677812
transform 1 0 2564 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1332
timestamp 1677677812
transform 1 0 2572 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1115
timestamp 1677677812
transform 1 0 2572 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_992
timestamp 1677677812
transform 1 0 2596 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1221
timestamp 1677677812
transform 1 0 2596 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1222
timestamp 1677677812
transform 1 0 2604 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_993
timestamp 1677677812
transform 1 0 2620 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1333
timestamp 1677677812
transform 1 0 2620 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1085
timestamp 1677677812
transform 1 0 2620 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1116
timestamp 1677677812
transform 1 0 2620 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1223
timestamp 1677677812
transform 1 0 2636 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1159
timestamp 1677677812
transform 1 0 2724 0 1 4145
box -2 -2 2 2
use M3_M2  M3_M2_1050
timestamp 1677677812
transform 1 0 2724 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1334
timestamp 1677677812
transform 1 0 2660 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1335
timestamp 1677677812
transform 1 0 2716 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1086
timestamp 1677677812
transform 1 0 2660 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1160
timestamp 1677677812
transform 1 0 2772 0 1 4145
box -2 -2 2 2
use M3_M2  M3_M2_1066
timestamp 1677677812
transform 1 0 2772 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1224
timestamp 1677677812
transform 1 0 2868 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1336
timestamp 1677677812
transform 1 0 2860 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1225
timestamp 1677677812
transform 1 0 2900 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1226
timestamp 1677677812
transform 1 0 2908 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1337
timestamp 1677677812
transform 1 0 2892 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1149
timestamp 1677677812
transform 1 0 2884 0 1 4085
box -3 -3 3 3
use M3_M2  M3_M2_1067
timestamp 1677677812
transform 1 0 2900 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1389
timestamp 1677677812
transform 1 0 2940 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1117
timestamp 1677677812
transform 1 0 2940 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_994
timestamp 1677677812
transform 1 0 2972 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1227
timestamp 1677677812
transform 1 0 2988 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1228
timestamp 1677677812
transform 1 0 2996 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1338
timestamp 1677677812
transform 1 0 2996 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1339
timestamp 1677677812
transform 1 0 3012 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1390
timestamp 1677677812
transform 1 0 2972 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1391
timestamp 1677677812
transform 1 0 2980 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1118
timestamp 1677677812
transform 1 0 2972 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1087
timestamp 1677677812
transform 1 0 2988 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1018
timestamp 1677677812
transform 1 0 3036 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1229
timestamp 1677677812
transform 1 0 3036 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1230
timestamp 1677677812
transform 1 0 3052 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1231
timestamp 1677677812
transform 1 0 3068 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1340
timestamp 1677677812
transform 1 0 3060 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1341
timestamp 1677677812
transform 1 0 3076 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1088
timestamp 1677677812
transform 1 0 3076 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1119
timestamp 1677677812
transform 1 0 3060 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1342
timestamp 1677677812
transform 1 0 3092 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1089
timestamp 1677677812
transform 1 0 3092 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1232
timestamp 1677677812
transform 1 0 3108 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1233
timestamp 1677677812
transform 1 0 3124 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1234
timestamp 1677677812
transform 1 0 3156 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1019
timestamp 1677677812
transform 1 0 3172 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1051
timestamp 1677677812
transform 1 0 3172 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1235
timestamp 1677677812
transform 1 0 3180 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1343
timestamp 1677677812
transform 1 0 3172 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1344
timestamp 1677677812
transform 1 0 3188 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1090
timestamp 1677677812
transform 1 0 3180 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1120
timestamp 1677677812
transform 1 0 3172 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1121
timestamp 1677677812
transform 1 0 3188 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1122
timestamp 1677677812
transform 1 0 3204 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1020
timestamp 1677677812
transform 1 0 3220 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1236
timestamp 1677677812
transform 1 0 3228 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1123
timestamp 1677677812
transform 1 0 3228 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1021
timestamp 1677677812
transform 1 0 3292 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1237
timestamp 1677677812
transform 1 0 3244 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1345
timestamp 1677677812
transform 1 0 3268 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1091
timestamp 1677677812
transform 1 0 3268 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_968
timestamp 1677677812
transform 1 0 3372 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1052
timestamp 1677677812
transform 1 0 3364 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1346
timestamp 1677677812
transform 1 0 3364 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1347
timestamp 1677677812
transform 1 0 3388 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1238
timestamp 1677677812
transform 1 0 3404 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1141
timestamp 1677677812
transform 1 0 3404 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1068
timestamp 1677677812
transform 1 0 3420 0 1 4125
box -3 -3 3 3
use M3_M2  M3_M2_969
timestamp 1677677812
transform 1 0 3444 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1239
timestamp 1677677812
transform 1 0 3452 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1053
timestamp 1677677812
transform 1 0 3460 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1240
timestamp 1677677812
transform 1 0 3484 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1348
timestamp 1677677812
transform 1 0 3460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1349
timestamp 1677677812
transform 1 0 3476 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1350
timestamp 1677677812
transform 1 0 3492 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1124
timestamp 1677677812
transform 1 0 3500 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1142
timestamp 1677677812
transform 1 0 3492 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1392
timestamp 1677677812
transform 1 0 3524 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_995
timestamp 1677677812
transform 1 0 3564 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1351
timestamp 1677677812
transform 1 0 3572 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1092
timestamp 1677677812
transform 1 0 3572 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1396
timestamp 1677677812
transform 1 0 3564 0 1 4105
box -2 -2 2 2
use M3_M2  M3_M2_996
timestamp 1677677812
transform 1 0 3604 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1352
timestamp 1677677812
transform 1 0 3596 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1125
timestamp 1677677812
transform 1 0 3588 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1393
timestamp 1677677812
transform 1 0 3604 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1143
timestamp 1677677812
transform 1 0 3596 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_970
timestamp 1677677812
transform 1 0 3692 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1241
timestamp 1677677812
transform 1 0 3620 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1242
timestamp 1677677812
transform 1 0 3644 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1353
timestamp 1677677812
transform 1 0 3628 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1093
timestamp 1677677812
transform 1 0 3628 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1054
timestamp 1677677812
transform 1 0 3652 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1243
timestamp 1677677812
transform 1 0 3668 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1055
timestamp 1677677812
transform 1 0 3700 0 1 4135
box -3 -3 3 3
use M3_M2  M3_M2_1056
timestamp 1677677812
transform 1 0 3716 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1354
timestamp 1677677812
transform 1 0 3652 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1355
timestamp 1677677812
transform 1 0 3716 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1126
timestamp 1677677812
transform 1 0 3660 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_971
timestamp 1677677812
transform 1 0 3772 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1244
timestamp 1677677812
transform 1 0 3772 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1356
timestamp 1677677812
transform 1 0 3788 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1357
timestamp 1677677812
transform 1 0 3796 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1094
timestamp 1677677812
transform 1 0 3788 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1127
timestamp 1677677812
transform 1 0 3780 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_997
timestamp 1677677812
transform 1 0 3844 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1057
timestamp 1677677812
transform 1 0 3820 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1245
timestamp 1677677812
transform 1 0 3828 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1358
timestamp 1677677812
transform 1 0 3820 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1359
timestamp 1677677812
transform 1 0 3836 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1095
timestamp 1677677812
transform 1 0 3836 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1246
timestamp 1677677812
transform 1 0 3852 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1360
timestamp 1677677812
transform 1 0 3868 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_998
timestamp 1677677812
transform 1 0 3908 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1247
timestamp 1677677812
transform 1 0 3884 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1248
timestamp 1677677812
transform 1 0 3892 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1361
timestamp 1677677812
transform 1 0 3908 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1362
timestamp 1677677812
transform 1 0 3924 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1096
timestamp 1677677812
transform 1 0 3892 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1128
timestamp 1677677812
transform 1 0 3916 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_972
timestamp 1677677812
transform 1 0 3940 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_973
timestamp 1677677812
transform 1 0 3956 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_974
timestamp 1677677812
transform 1 0 4004 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_999
timestamp 1677677812
transform 1 0 3980 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1000
timestamp 1677677812
transform 1 0 4012 0 1 4155
box -3 -3 3 3
use M2_M1  M2_M1_1249
timestamp 1677677812
transform 1 0 3964 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1250
timestamp 1677677812
transform 1 0 3972 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1251
timestamp 1677677812
transform 1 0 3988 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1252
timestamp 1677677812
transform 1 0 4004 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1097
timestamp 1677677812
transform 1 0 3964 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1363
timestamp 1677677812
transform 1 0 3980 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1364
timestamp 1677677812
transform 1 0 3996 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1098
timestamp 1677677812
transform 1 0 3996 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1365
timestamp 1677677812
transform 1 0 4012 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1099
timestamp 1677677812
transform 1 0 4012 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_975
timestamp 1677677812
transform 1 0 4084 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_976
timestamp 1677677812
transform 1 0 4132 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1253
timestamp 1677677812
transform 1 0 4052 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1254
timestamp 1677677812
transform 1 0 4068 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1366
timestamp 1677677812
transform 1 0 4116 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1100
timestamp 1677677812
transform 1 0 4116 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1129
timestamp 1677677812
transform 1 0 4068 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1130
timestamp 1677677812
transform 1 0 4108 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1022
timestamp 1677677812
transform 1 0 4196 0 1 4145
box -3 -3 3 3
use M3_M2  M3_M2_1058
timestamp 1677677812
transform 1 0 4188 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1255
timestamp 1677677812
transform 1 0 4196 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1256
timestamp 1677677812
transform 1 0 4212 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1059
timestamp 1677677812
transform 1 0 4220 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1367
timestamp 1677677812
transform 1 0 4188 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1069
timestamp 1677677812
transform 1 0 4196 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1368
timestamp 1677677812
transform 1 0 4204 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1369
timestamp 1677677812
transform 1 0 4220 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1101
timestamp 1677677812
transform 1 0 4212 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1144
timestamp 1677677812
transform 1 0 4204 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1257
timestamp 1677677812
transform 1 0 4236 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1145
timestamp 1677677812
transform 1 0 4236 0 1 4095
box -3 -3 3 3
use M2_M1  M2_M1_1370
timestamp 1677677812
transform 1 0 4276 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1394
timestamp 1677677812
transform 1 0 4260 0 1 4115
box -2 -2 2 2
use M3_M2  M3_M2_1102
timestamp 1677677812
transform 1 0 4276 0 1 4115
box -3 -3 3 3
use M2_M1  M2_M1_1395
timestamp 1677677812
transform 1 0 4284 0 1 4115
box -2 -2 2 2
use M2_M1  M2_M1_1397
timestamp 1677677812
transform 1 0 4268 0 1 4105
box -2 -2 2 2
use M3_M2  M3_M2_1131
timestamp 1677677812
transform 1 0 4284 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1258
timestamp 1677677812
transform 1 0 4308 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1060
timestamp 1677677812
transform 1 0 4316 0 1 4135
box -3 -3 3 3
use M2_M1  M2_M1_1371
timestamp 1677677812
transform 1 0 4300 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1372
timestamp 1677677812
transform 1 0 4316 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1373
timestamp 1677677812
transform 1 0 4332 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1132
timestamp 1677677812
transform 1 0 4316 0 1 4105
box -3 -3 3 3
use M2_M1  M2_M1_1374
timestamp 1677677812
transform 1 0 4348 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1023
timestamp 1677677812
transform 1 0 4388 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1259
timestamp 1677677812
transform 1 0 4364 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1260
timestamp 1677677812
transform 1 0 4372 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1261
timestamp 1677677812
transform 1 0 4388 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1262
timestamp 1677677812
transform 1 0 4404 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_1070
timestamp 1677677812
transform 1 0 4372 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1375
timestamp 1677677812
transform 1 0 4396 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1103
timestamp 1677677812
transform 1 0 4364 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1104
timestamp 1677677812
transform 1 0 4396 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1024
timestamp 1677677812
transform 1 0 4460 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1263
timestamp 1677677812
transform 1 0 4436 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1376
timestamp 1677677812
transform 1 0 4460 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1377
timestamp 1677677812
transform 1 0 4516 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1071
timestamp 1677677812
transform 1 0 4540 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1264
timestamp 1677677812
transform 1 0 4564 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1265
timestamp 1677677812
transform 1 0 4580 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1266
timestamp 1677677812
transform 1 0 4588 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1267
timestamp 1677677812
transform 1 0 4596 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1378
timestamp 1677677812
transform 1 0 4556 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1379
timestamp 1677677812
transform 1 0 4572 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1105
timestamp 1677677812
transform 1 0 4564 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1133
timestamp 1677677812
transform 1 0 4572 0 1 4105
box -3 -3 3 3
use M3_M2  M3_M2_1146
timestamp 1677677812
transform 1 0 4556 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_1072
timestamp 1677677812
transform 1 0 4596 0 1 4125
box -3 -3 3 3
use M2_M1  M2_M1_1380
timestamp 1677677812
transform 1 0 4612 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1001
timestamp 1677677812
transform 1 0 4636 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1002
timestamp 1677677812
transform 1 0 4652 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1025
timestamp 1677677812
transform 1 0 4644 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1268
timestamp 1677677812
transform 1 0 4644 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1381
timestamp 1677677812
transform 1 0 4628 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1382
timestamp 1677677812
transform 1 0 4652 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1106
timestamp 1677677812
transform 1 0 4652 0 1 4115
box -3 -3 3 3
use M3_M2  M3_M2_1147
timestamp 1677677812
transform 1 0 4652 0 1 4095
box -3 -3 3 3
use M3_M2  M3_M2_977
timestamp 1677677812
transform 1 0 4676 0 1 4165
box -3 -3 3 3
use M2_M1  M2_M1_1269
timestamp 1677677812
transform 1 0 4676 0 1 4135
box -2 -2 2 2
use M3_M2  M3_M2_978
timestamp 1677677812
transform 1 0 4740 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_979
timestamp 1677677812
transform 1 0 4756 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_980
timestamp 1677677812
transform 1 0 4780 0 1 4165
box -3 -3 3 3
use M3_M2  M3_M2_1003
timestamp 1677677812
transform 1 0 4716 0 1 4155
box -3 -3 3 3
use M3_M2  M3_M2_1026
timestamp 1677677812
transform 1 0 4724 0 1 4145
box -3 -3 3 3
use M2_M1  M2_M1_1270
timestamp 1677677812
transform 1 0 4700 0 1 4135
box -2 -2 2 2
use M2_M1  M2_M1_1383
timestamp 1677677812
transform 1 0 4724 0 1 4125
box -2 -2 2 2
use M2_M1  M2_M1_1384
timestamp 1677677812
transform 1 0 4780 0 1 4125
box -2 -2 2 2
use M3_M2  M3_M2_1107
timestamp 1677677812
transform 1 0 4748 0 1 4115
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_12
timestamp 1677677812
transform 1 0 24 0 1 4070
box -10 -3 10 3
use FILL  FILL_817
timestamp 1677677812
transform 1 0 72 0 -1 4170
box -8 -3 16 105
use FILL  FILL_818
timestamp 1677677812
transform 1 0 80 0 -1 4170
box -8 -3 16 105
use FILL  FILL_819
timestamp 1677677812
transform 1 0 88 0 -1 4170
box -8 -3 16 105
use FILL  FILL_820
timestamp 1677677812
transform 1 0 96 0 -1 4170
box -8 -3 16 105
use FILL  FILL_821
timestamp 1677677812
transform 1 0 104 0 -1 4170
box -8 -3 16 105
use FILL  FILL_822
timestamp 1677677812
transform 1 0 112 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_81
timestamp 1677677812
transform -1 0 136 0 -1 4170
box -9 -3 26 105
use FILL  FILL_823
timestamp 1677677812
transform 1 0 136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_824
timestamp 1677677812
transform 1 0 144 0 -1 4170
box -8 -3 16 105
use FILL  FILL_825
timestamp 1677677812
transform 1 0 152 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_42
timestamp 1677677812
transform -1 0 200 0 -1 4170
box -8 -3 46 105
use INVX2  INVX2_82
timestamp 1677677812
transform 1 0 200 0 -1 4170
box -9 -3 26 105
use FILL  FILL_826
timestamp 1677677812
transform 1 0 216 0 -1 4170
box -8 -3 16 105
use FILL  FILL_835
timestamp 1677677812
transform 1 0 224 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1150
timestamp 1677677812
transform 1 0 244 0 1 4075
box -3 -3 3 3
use FILL  FILL_836
timestamp 1677677812
transform 1 0 232 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_84
timestamp 1677677812
transform -1 0 256 0 -1 4170
box -9 -3 26 105
use M3_M2  M3_M2_1151
timestamp 1677677812
transform 1 0 300 0 1 4075
box -3 -3 3 3
use OAI22X1  OAI22X1_41
timestamp 1677677812
transform 1 0 256 0 -1 4170
box -8 -3 46 105
use INVX2  INVX2_85
timestamp 1677677812
transform 1 0 296 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_72
timestamp 1677677812
transform 1 0 312 0 -1 4170
box -8 -3 104 105
use INVX2  INVX2_86
timestamp 1677677812
transform -1 0 424 0 -1 4170
box -9 -3 26 105
use FILL  FILL_837
timestamp 1677677812
transform 1 0 424 0 -1 4170
box -8 -3 16 105
use FILL  FILL_838
timestamp 1677677812
transform 1 0 432 0 -1 4170
box -8 -3 16 105
use FILL  FILL_839
timestamp 1677677812
transform 1 0 440 0 -1 4170
box -8 -3 16 105
use FILL  FILL_840
timestamp 1677677812
transform 1 0 448 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_45
timestamp 1677677812
transform -1 0 496 0 -1 4170
box -8 -3 46 105
use FILL  FILL_841
timestamp 1677677812
transform 1 0 496 0 -1 4170
box -8 -3 16 105
use FILL  FILL_842
timestamp 1677677812
transform 1 0 504 0 -1 4170
box -8 -3 16 105
use FILL  FILL_843
timestamp 1677677812
transform 1 0 512 0 -1 4170
box -8 -3 16 105
use FILL  FILL_844
timestamp 1677677812
transform 1 0 520 0 -1 4170
box -8 -3 16 105
use FILL  FILL_845
timestamp 1677677812
transform 1 0 528 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_87
timestamp 1677677812
transform -1 0 552 0 -1 4170
box -9 -3 26 105
use INVX2  INVX2_88
timestamp 1677677812
transform -1 0 568 0 -1 4170
box -9 -3 26 105
use FILL  FILL_846
timestamp 1677677812
transform 1 0 568 0 -1 4170
box -8 -3 16 105
use FILL  FILL_848
timestamp 1677677812
transform 1 0 576 0 -1 4170
box -8 -3 16 105
use FILL  FILL_850
timestamp 1677677812
transform 1 0 584 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_47
timestamp 1677677812
transform 1 0 592 0 -1 4170
box -8 -3 46 105
use FILL  FILL_853
timestamp 1677677812
transform 1 0 632 0 -1 4170
box -8 -3 16 105
use FILL  FILL_854
timestamp 1677677812
transform 1 0 640 0 -1 4170
box -8 -3 16 105
use FILL  FILL_856
timestamp 1677677812
transform 1 0 648 0 -1 4170
box -8 -3 16 105
use FILL  FILL_858
timestamp 1677677812
transform 1 0 656 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_43
timestamp 1677677812
transform 1 0 664 0 -1 4170
box -8 -3 46 105
use FILL  FILL_861
timestamp 1677677812
transform 1 0 704 0 -1 4170
box -8 -3 16 105
use FILL  FILL_862
timestamp 1677677812
transform 1 0 712 0 -1 4170
box -8 -3 16 105
use FILL  FILL_864
timestamp 1677677812
transform 1 0 720 0 -1 4170
box -8 -3 16 105
use FILL  FILL_866
timestamp 1677677812
transform 1 0 728 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_74
timestamp 1677677812
transform -1 0 832 0 -1 4170
box -8 -3 104 105
use FILL  FILL_868
timestamp 1677677812
transform 1 0 832 0 -1 4170
box -8 -3 16 105
use FILL  FILL_870
timestamp 1677677812
transform 1 0 840 0 -1 4170
box -8 -3 16 105
use FILL  FILL_872
timestamp 1677677812
transform 1 0 848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_873
timestamp 1677677812
transform 1 0 856 0 -1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_11
timestamp 1677677812
transform 1 0 864 0 -1 4170
box -8 -3 32 105
use FILL  FILL_874
timestamp 1677677812
transform 1 0 888 0 -1 4170
box -8 -3 16 105
use FILL  FILL_875
timestamp 1677677812
transform 1 0 896 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_48
timestamp 1677677812
transform 1 0 904 0 -1 4170
box -8 -3 46 105
use FILL  FILL_876
timestamp 1677677812
transform 1 0 944 0 -1 4170
box -8 -3 16 105
use FILL  FILL_878
timestamp 1677677812
transform 1 0 952 0 -1 4170
box -8 -3 16 105
use FILL  FILL_879
timestamp 1677677812
transform 1 0 960 0 -1 4170
box -8 -3 16 105
use FILL  FILL_880
timestamp 1677677812
transform 1 0 968 0 -1 4170
box -8 -3 16 105
use FILL  FILL_882
timestamp 1677677812
transform 1 0 976 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_24
timestamp 1677677812
transform 1 0 984 0 -1 4170
box -8 -3 34 105
use FILL  FILL_886
timestamp 1677677812
transform 1 0 1016 0 -1 4170
box -8 -3 16 105
use FILL  FILL_887
timestamp 1677677812
transform 1 0 1024 0 -1 4170
box -8 -3 16 105
use FILL  FILL_889
timestamp 1677677812
transform 1 0 1032 0 -1 4170
box -8 -3 16 105
use FILL  FILL_891
timestamp 1677677812
transform 1 0 1040 0 -1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_13
timestamp 1677677812
transform 1 0 1048 0 -1 4170
box -8 -3 32 105
use FILL  FILL_893
timestamp 1677677812
transform 1 0 1072 0 -1 4170
box -8 -3 16 105
use FILL  FILL_894
timestamp 1677677812
transform 1 0 1080 0 -1 4170
box -8 -3 16 105
use FILL  FILL_896
timestamp 1677677812
transform 1 0 1088 0 -1 4170
box -8 -3 16 105
use FILL  FILL_898
timestamp 1677677812
transform 1 0 1096 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_26
timestamp 1677677812
transform 1 0 1104 0 -1 4170
box -8 -3 34 105
use FILL  FILL_900
timestamp 1677677812
transform 1 0 1136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_901
timestamp 1677677812
transform 1 0 1144 0 -1 4170
box -8 -3 16 105
use FILL  FILL_903
timestamp 1677677812
transform 1 0 1152 0 -1 4170
box -8 -3 16 105
use FILL  FILL_912
timestamp 1677677812
transform 1 0 1160 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_91
timestamp 1677677812
transform 1 0 1168 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_78
timestamp 1677677812
transform -1 0 1280 0 -1 4170
box -8 -3 104 105
use FILL  FILL_913
timestamp 1677677812
transform 1 0 1280 0 -1 4170
box -8 -3 16 105
use FILL  FILL_914
timestamp 1677677812
transform 1 0 1288 0 -1 4170
box -8 -3 16 105
use FILL  FILL_915
timestamp 1677677812
transform 1 0 1296 0 -1 4170
box -8 -3 16 105
use FILL  FILL_916
timestamp 1677677812
transform 1 0 1304 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_28
timestamp 1677677812
transform -1 0 1344 0 -1 4170
box -8 -3 34 105
use FILL  FILL_917
timestamp 1677677812
transform 1 0 1344 0 -1 4170
box -8 -3 16 105
use FILL  FILL_918
timestamp 1677677812
transform 1 0 1352 0 -1 4170
box -8 -3 16 105
use FILL  FILL_919
timestamp 1677677812
transform 1 0 1360 0 -1 4170
box -8 -3 16 105
use FILL  FILL_920
timestamp 1677677812
transform 1 0 1368 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_92
timestamp 1677677812
transform 1 0 1376 0 -1 4170
box -9 -3 26 105
use FILL  FILL_921
timestamp 1677677812
transform 1 0 1392 0 -1 4170
box -8 -3 16 105
use FILL  FILL_922
timestamp 1677677812
transform 1 0 1400 0 -1 4170
box -8 -3 16 105
use FILL  FILL_923
timestamp 1677677812
transform 1 0 1408 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_44
timestamp 1677677812
transform -1 0 1456 0 -1 4170
box -8 -3 46 105
use FILL  FILL_924
timestamp 1677677812
transform 1 0 1456 0 -1 4170
box -8 -3 16 105
use FILL  FILL_926
timestamp 1677677812
transform 1 0 1464 0 -1 4170
box -8 -3 16 105
use FILL  FILL_933
timestamp 1677677812
transform 1 0 1472 0 -1 4170
box -8 -3 16 105
use FILL  FILL_934
timestamp 1677677812
transform 1 0 1480 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_79
timestamp 1677677812
transform 1 0 1488 0 -1 4170
box -8 -3 104 105
use FILL  FILL_935
timestamp 1677677812
transform 1 0 1584 0 -1 4170
box -8 -3 16 105
use FILL  FILL_937
timestamp 1677677812
transform 1 0 1592 0 -1 4170
box -8 -3 16 105
use FILL  FILL_942
timestamp 1677677812
transform 1 0 1600 0 -1 4170
box -8 -3 16 105
use FILL  FILL_943
timestamp 1677677812
transform 1 0 1608 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_46
timestamp 1677677812
transform -1 0 1656 0 -1 4170
box -8 -3 46 105
use FILL  FILL_944
timestamp 1677677812
transform 1 0 1656 0 -1 4170
box -8 -3 16 105
use FILL  FILL_945
timestamp 1677677812
transform 1 0 1664 0 -1 4170
box -8 -3 16 105
use FILL  FILL_946
timestamp 1677677812
transform 1 0 1672 0 -1 4170
box -8 -3 16 105
use FILL  FILL_948
timestamp 1677677812
transform 1 0 1680 0 -1 4170
box -8 -3 16 105
use FILL  FILL_952
timestamp 1677677812
transform 1 0 1688 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_81
timestamp 1677677812
transform 1 0 1696 0 -1 4170
box -8 -3 104 105
use FILL  FILL_953
timestamp 1677677812
transform 1 0 1792 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_99
timestamp 1677677812
transform -1 0 1816 0 -1 4170
box -9 -3 26 105
use FILL  FILL_954
timestamp 1677677812
transform 1 0 1816 0 -1 4170
box -8 -3 16 105
use FILL  FILL_956
timestamp 1677677812
transform 1 0 1824 0 -1 4170
box -8 -3 16 105
use FILL  FILL_958
timestamp 1677677812
transform 1 0 1832 0 -1 4170
box -8 -3 16 105
use FILL  FILL_962
timestamp 1677677812
transform 1 0 1840 0 -1 4170
box -8 -3 16 105
use FILL  FILL_963
timestamp 1677677812
transform 1 0 1848 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_51
timestamp 1677677812
transform 1 0 1856 0 -1 4170
box -8 -3 46 105
use FILL  FILL_964
timestamp 1677677812
transform 1 0 1896 0 -1 4170
box -8 -3 16 105
use FILL  FILL_967
timestamp 1677677812
transform 1 0 1904 0 -1 4170
box -8 -3 16 105
use FILL  FILL_968
timestamp 1677677812
transform 1 0 1912 0 -1 4170
box -8 -3 16 105
use FILL  FILL_969
timestamp 1677677812
transform 1 0 1920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_970
timestamp 1677677812
transform 1 0 1928 0 -1 4170
box -8 -3 16 105
use FILL  FILL_971
timestamp 1677677812
transform 1 0 1936 0 -1 4170
box -8 -3 16 105
use FILL  FILL_972
timestamp 1677677812
transform 1 0 1944 0 -1 4170
box -8 -3 16 105
use FILL  FILL_974
timestamp 1677677812
transform 1 0 1952 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_47
timestamp 1677677812
transform 1 0 1960 0 -1 4170
box -8 -3 46 105
use FILL  FILL_977
timestamp 1677677812
transform 1 0 2000 0 -1 4170
box -8 -3 16 105
use FILL  FILL_978
timestamp 1677677812
transform 1 0 2008 0 -1 4170
box -8 -3 16 105
use FILL  FILL_980
timestamp 1677677812
transform 1 0 2016 0 -1 4170
box -8 -3 16 105
use FILL  FILL_988
timestamp 1677677812
transform 1 0 2024 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_53
timestamp 1677677812
transform -1 0 2072 0 -1 4170
box -8 -3 46 105
use FILL  FILL_989
timestamp 1677677812
transform 1 0 2072 0 -1 4170
box -8 -3 16 105
use FILL  FILL_991
timestamp 1677677812
transform 1 0 2080 0 -1 4170
box -8 -3 16 105
use FILL  FILL_993
timestamp 1677677812
transform 1 0 2088 0 -1 4170
box -8 -3 16 105
use FILL  FILL_995
timestamp 1677677812
transform 1 0 2096 0 -1 4170
box -8 -3 16 105
use FILL  FILL_996
timestamp 1677677812
transform 1 0 2104 0 -1 4170
box -8 -3 16 105
use FILL  FILL_997
timestamp 1677677812
transform 1 0 2112 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1677677812
transform 1 0 2120 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_83
timestamp 1677677812
transform -1 0 2224 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1010
timestamp 1677677812
transform 1 0 2224 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1011
timestamp 1677677812
transform 1 0 2232 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1677677812
transform 1 0 2240 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1677677812
transform 1 0 2248 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1677677812
transform 1 0 2256 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1677677812
transform 1 0 2264 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1677677812
transform 1 0 2272 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1677677812
transform 1 0 2280 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1677677812
transform 1 0 2288 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1677677812
transform 1 0 2296 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1677677812
transform 1 0 2304 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1677677812
transform 1 0 2312 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1677677812
transform 1 0 2320 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1677677812
transform 1 0 2328 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1677677812
transform 1 0 2336 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1677677812
transform 1 0 2344 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1677677812
transform 1 0 2352 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1029
timestamp 1677677812
transform 1 0 2360 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1677677812
transform 1 0 2368 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1677677812
transform 1 0 2376 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1677677812
transform 1 0 2384 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_49
timestamp 1677677812
transform -1 0 2432 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1041
timestamp 1677677812
transform 1 0 2432 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1043
timestamp 1677677812
transform 1 0 2440 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1677677812
transform 1 0 2448 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1677677812
transform 1 0 2456 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1677677812
transform 1 0 2464 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_104
timestamp 1677677812
transform 1 0 2472 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1053
timestamp 1677677812
transform 1 0 2488 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1677677812
transform 1 0 2496 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1677677812
transform 1 0 2504 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1677677812
transform 1 0 2512 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_55
timestamp 1677677812
transform 1 0 2520 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1067
timestamp 1677677812
transform 1 0 2560 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1677677812
transform 1 0 2568 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1677677812
transform 1 0 2576 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1070
timestamp 1677677812
transform 1 0 2584 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1071
timestamp 1677677812
transform 1 0 2592 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_106
timestamp 1677677812
transform 1 0 2600 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1072
timestamp 1677677812
transform 1 0 2616 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_85
timestamp 1677677812
transform 1 0 2624 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1073
timestamp 1677677812
transform 1 0 2720 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1677677812
transform 1 0 2728 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1677677812
transform 1 0 2736 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1152
timestamp 1677677812
transform 1 0 2756 0 1 4075
box -3 -3 3 3
use FILL  FILL_1081
timestamp 1677677812
transform 1 0 2744 0 -1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1677677812
transform 1 0 2752 0 -1 4170
box -8 -3 32 105
use FILL  FILL_1082
timestamp 1677677812
transform 1 0 2776 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1083
timestamp 1677677812
transform 1 0 2784 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1084
timestamp 1677677812
transform 1 0 2792 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1677677812
transform 1 0 2800 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1677677812
transform 1 0 2808 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1677677812
transform 1 0 2816 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1088
timestamp 1677677812
transform 1 0 2824 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1677677812
transform 1 0 2832 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1090
timestamp 1677677812
transform 1 0 2840 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1677677812
transform 1 0 2848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1677677812
transform 1 0 2856 0 -1 4170
box -8 -3 16 105
use NOR2X1  NOR2X1_15
timestamp 1677677812
transform 1 0 2864 0 -1 4170
box -8 -3 32 105
use FILL  FILL_1093
timestamp 1677677812
transform 1 0 2888 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1677677812
transform 1 0 2896 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1677677812
transform 1 0 2904 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1677677812
transform 1 0 2912 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1677677812
transform 1 0 2920 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1677677812
transform 1 0 2928 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_31
timestamp 1677677812
transform -1 0 2968 0 -1 4170
box -8 -3 34 105
use FILL  FILL_1103
timestamp 1677677812
transform 1 0 2968 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1104
timestamp 1677677812
transform 1 0 2976 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1677677812
transform 1 0 2984 0 -1 4170
box -8 -3 16 105
use OAI21X1  OAI21X1_32
timestamp 1677677812
transform -1 0 3024 0 -1 4170
box -8 -3 34 105
use FILL  FILL_1112
timestamp 1677677812
transform 1 0 3024 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1677677812
transform 1 0 3032 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1677677812
transform 1 0 3040 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_50
timestamp 1677677812
transform 1 0 3048 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1119
timestamp 1677677812
transform 1 0 3088 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1677677812
transform 1 0 3096 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1128
timestamp 1677677812
transform 1 0 3104 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_108
timestamp 1677677812
transform -1 0 3128 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1129
timestamp 1677677812
transform 1 0 3128 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1677677812
transform 1 0 3136 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1677677812
transform 1 0 3144 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1132
timestamp 1677677812
transform 1 0 3152 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_52
timestamp 1677677812
transform -1 0 3200 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1133
timestamp 1677677812
transform 1 0 3200 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1677677812
transform 1 0 3208 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1144
timestamp 1677677812
transform 1 0 3216 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1145
timestamp 1677677812
transform 1 0 3224 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_87
timestamp 1677677812
transform 1 0 3232 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1146
timestamp 1677677812
transform 1 0 3328 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1677677812
transform 1 0 3336 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_110
timestamp 1677677812
transform 1 0 3344 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1153
timestamp 1677677812
transform 1 0 3360 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1677677812
transform 1 0 3368 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1155
timestamp 1677677812
transform 1 0 3376 0 -1 4170
box -8 -3 16 105
use BUFX2  BUFX2_2
timestamp 1677677812
transform 1 0 3384 0 -1 4170
box -5 -3 28 105
use FILL  FILL_1156
timestamp 1677677812
transform 1 0 3408 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1677677812
transform 1 0 3416 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1159
timestamp 1677677812
transform 1 0 3424 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1161
timestamp 1677677812
transform 1 0 3432 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1677677812
transform 1 0 3440 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1677677812
transform 1 0 3448 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_56
timestamp 1677677812
transform -1 0 3496 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1167
timestamp 1677677812
transform 1 0 3496 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1677677812
transform 1 0 3504 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1677677812
transform 1 0 3512 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1677677812
transform 1 0 3520 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1173
timestamp 1677677812
transform 1 0 3528 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1677677812
transform 1 0 3536 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1182
timestamp 1677677812
transform 1 0 3544 0 -1 4170
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1677677812
transform -1 0 3584 0 -1 4170
box -8 -3 40 105
use FILL  FILL_1183
timestamp 1677677812
transform 1 0 3584 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1677677812
transform 1 0 3592 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1677677812
transform 1 0 3600 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_57
timestamp 1677677812
transform 1 0 3608 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1189
timestamp 1677677812
transform 1 0 3648 0 -1 4170
box -8 -3 16 105
use M3_M2  M3_M2_1153
timestamp 1677677812
transform 1 0 3668 0 1 4075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_89
timestamp 1677677812
transform 1 0 3656 0 -1 4170
box -8 -3 104 105
use M3_M2  M3_M2_1154
timestamp 1677677812
transform 1 0 3764 0 1 4075
box -3 -3 3 3
use INVX2  INVX2_113
timestamp 1677677812
transform 1 0 3752 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1194
timestamp 1677677812
transform 1 0 3768 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1677677812
transform 1 0 3776 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1677677812
transform 1 0 3784 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1677677812
transform 1 0 3792 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1677677812
transform 1 0 3800 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_56
timestamp 1677677812
transform 1 0 3808 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1203
timestamp 1677677812
transform 1 0 3848 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1677677812
transform 1 0 3856 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1677677812
transform 1 0 3864 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1677677812
transform 1 0 3872 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1211
timestamp 1677677812
transform 1 0 3880 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_59
timestamp 1677677812
transform -1 0 3928 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1212
timestamp 1677677812
transform 1 0 3928 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1677677812
transform 1 0 3936 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1215
timestamp 1677677812
transform 1 0 3944 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1677677812
transform 1 0 3952 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1677677812
transform 1 0 3960 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_59
timestamp 1677677812
transform 1 0 3968 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1224
timestamp 1677677812
transform 1 0 4008 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1677677812
transform 1 0 4016 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1226
timestamp 1677677812
transform 1 0 4024 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1677677812
transform 1 0 4032 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_115
timestamp 1677677812
transform -1 0 4056 0 -1 4170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_92
timestamp 1677677812
transform 1 0 4056 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1228
timestamp 1677677812
transform 1 0 4152 0 -1 4170
box -8 -3 16 105
use INVX2  INVX2_116
timestamp 1677677812
transform 1 0 4160 0 -1 4170
box -9 -3 26 105
use FILL  FILL_1229
timestamp 1677677812
transform 1 0 4176 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1677677812
transform 1 0 4184 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_60
timestamp 1677677812
transform 1 0 4192 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1231
timestamp 1677677812
transform 1 0 4232 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1232
timestamp 1677677812
transform 1 0 4240 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1234
timestamp 1677677812
transform 1 0 4248 0 -1 4170
box -8 -3 16 105
use NAND3X1  NAND3X1_6
timestamp 1677677812
transform -1 0 4288 0 -1 4170
box -8 -3 40 105
use FILL  FILL_1236
timestamp 1677677812
transform 1 0 4288 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_61
timestamp 1677677812
transform -1 0 4336 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1238
timestamp 1677677812
transform 1 0 4336 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1677677812
transform 1 0 4344 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1677677812
transform 1 0 4352 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1245
timestamp 1677677812
transform 1 0 4360 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_62
timestamp 1677677812
transform 1 0 4368 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1246
timestamp 1677677812
transform 1 0 4408 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1677677812
transform 1 0 4416 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_94
timestamp 1677677812
transform 1 0 4424 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1249
timestamp 1677677812
transform 1 0 4520 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1677677812
transform 1 0 4528 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1677677812
transform 1 0 4536 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1677677812
transform 1 0 4544 0 -1 4170
box -8 -3 16 105
use AOI22X1  AOI22X1_63
timestamp 1677677812
transform 1 0 4552 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1256
timestamp 1677677812
transform 1 0 4592 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1677677812
transform 1 0 4600 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1677677812
transform 1 0 4608 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1262
timestamp 1677677812
transform 1 0 4616 0 -1 4170
box -8 -3 16 105
use OAI22X1  OAI22X1_64
timestamp 1677677812
transform 1 0 4624 0 -1 4170
box -8 -3 46 105
use FILL  FILL_1263
timestamp 1677677812
transform 1 0 4664 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1677677812
transform 1 0 4672 0 -1 4170
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1677677812
transform 1 0 4680 0 -1 4170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_96
timestamp 1677677812
transform 1 0 4688 0 -1 4170
box -8 -3 104 105
use FILL  FILL_1266
timestamp 1677677812
transform 1 0 4784 0 -1 4170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_13
timestamp 1677677812
transform 1 0 4843 0 1 4070
box -10 -3 10 3
use M3_M2  M3_M2_1185
timestamp 1677677812
transform 1 0 84 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1202
timestamp 1677677812
transform 1 0 156 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1411
timestamp 1677677812
transform 1 0 116 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1523
timestamp 1677677812
transform 1 0 84 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1412
timestamp 1677677812
transform 1 0 172 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1203
timestamp 1677677812
transform 1 0 196 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1413
timestamp 1677677812
transform 1 0 196 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1414
timestamp 1677677812
transform 1 0 212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1415
timestamp 1677677812
transform 1 0 228 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1524
timestamp 1677677812
transform 1 0 188 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1525
timestamp 1677677812
transform 1 0 220 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1167
timestamp 1677677812
transform 1 0 244 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1204
timestamp 1677677812
transform 1 0 244 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1416
timestamp 1677677812
transform 1 0 244 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1526
timestamp 1677677812
transform 1 0 252 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1205
timestamp 1677677812
transform 1 0 308 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1417
timestamp 1677677812
transform 1 0 284 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1418
timestamp 1677677812
transform 1 0 300 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1186
timestamp 1677677812
transform 1 0 324 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1206
timestamp 1677677812
transform 1 0 356 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1419
timestamp 1677677812
transform 1 0 324 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1420
timestamp 1677677812
transform 1 0 356 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1527
timestamp 1677677812
transform 1 0 404 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1207
timestamp 1677677812
transform 1 0 492 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1421
timestamp 1677677812
transform 1 0 492 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1528
timestamp 1677677812
transform 1 0 444 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1208
timestamp 1677677812
transform 1 0 564 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1422
timestamp 1677677812
transform 1 0 556 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1423
timestamp 1677677812
transform 1 0 572 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1529
timestamp 1677677812
transform 1 0 564 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1530
timestamp 1677677812
transform 1 0 588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1278
timestamp 1677677812
transform 1 0 564 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1531
timestamp 1677677812
transform 1 0 604 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1209
timestamp 1677677812
transform 1 0 620 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1424
timestamp 1677677812
transform 1 0 620 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1425
timestamp 1677677812
transform 1 0 636 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1240
timestamp 1677677812
transform 1 0 644 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1532
timestamp 1677677812
transform 1 0 620 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1259
timestamp 1677677812
transform 1 0 636 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1533
timestamp 1677677812
transform 1 0 644 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1308
timestamp 1677677812
transform 1 0 620 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1309
timestamp 1677677812
transform 1 0 644 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1534
timestamp 1677677812
transform 1 0 660 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1279
timestamp 1677677812
transform 1 0 660 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1426
timestamp 1677677812
transform 1 0 684 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1427
timestamp 1677677812
transform 1 0 708 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1241
timestamp 1677677812
transform 1 0 732 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1535
timestamp 1677677812
transform 1 0 716 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1536
timestamp 1677677812
transform 1 0 732 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1310
timestamp 1677677812
transform 1 0 716 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1428
timestamp 1677677812
transform 1 0 748 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1429
timestamp 1677677812
transform 1 0 764 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1430
timestamp 1677677812
transform 1 0 812 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1537
timestamp 1677677812
transform 1 0 756 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1260
timestamp 1677677812
transform 1 0 764 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1538
timestamp 1677677812
transform 1 0 780 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1431
timestamp 1677677812
transform 1 0 876 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1261
timestamp 1677677812
transform 1 0 876 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1614
timestamp 1677677812
transform 1 0 868 0 1 3995
box -2 -2 2 2
use M3_M2  M3_M2_1311
timestamp 1677677812
transform 1 0 868 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1398
timestamp 1677677812
transform 1 0 900 0 1 4045
box -2 -2 2 2
use M2_M1  M2_M1_1539
timestamp 1677677812
transform 1 0 916 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1312
timestamp 1677677812
transform 1 0 924 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1262
timestamp 1677677812
transform 1 0 956 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1280
timestamp 1677677812
transform 1 0 964 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1399
timestamp 1677677812
transform 1 0 972 0 1 4045
box -2 -2 2 2
use M3_M2  M3_M2_1187
timestamp 1677677812
transform 1 0 972 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1210
timestamp 1677677812
transform 1 0 980 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1432
timestamp 1677677812
transform 1 0 972 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1540
timestamp 1677677812
transform 1 0 980 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1155
timestamp 1677677812
transform 1 0 1036 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1242
timestamp 1677677812
transform 1 0 1036 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1211
timestamp 1677677812
transform 1 0 1060 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1168
timestamp 1677677812
transform 1 0 1084 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1433
timestamp 1677677812
transform 1 0 1044 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1434
timestamp 1677677812
transform 1 0 1060 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1435
timestamp 1677677812
transform 1 0 1076 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1436
timestamp 1677677812
transform 1 0 1084 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1541
timestamp 1677677812
transform 1 0 1036 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1542
timestamp 1677677812
transform 1 0 1044 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1313
timestamp 1677677812
transform 1 0 1044 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1281
timestamp 1677677812
transform 1 0 1076 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1314
timestamp 1677677812
transform 1 0 1076 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1543
timestamp 1677677812
transform 1 0 1092 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1544
timestamp 1677677812
transform 1 0 1108 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1545
timestamp 1677677812
transform 1 0 1116 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1315
timestamp 1677677812
transform 1 0 1108 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1188
timestamp 1677677812
transform 1 0 1132 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1212
timestamp 1677677812
transform 1 0 1140 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1437
timestamp 1677677812
transform 1 0 1132 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1438
timestamp 1677677812
transform 1 0 1148 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1439
timestamp 1677677812
transform 1 0 1164 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1440
timestamp 1677677812
transform 1 0 1172 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1263
timestamp 1677677812
transform 1 0 1132 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1282
timestamp 1677677812
transform 1 0 1164 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1213
timestamp 1677677812
transform 1 0 1188 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1546
timestamp 1677677812
transform 1 0 1196 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1547
timestamp 1677677812
transform 1 0 1236 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1156
timestamp 1677677812
transform 1 0 1252 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1402
timestamp 1677677812
transform 1 0 1244 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1548
timestamp 1677677812
transform 1 0 1252 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1283
timestamp 1677677812
transform 1 0 1244 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1157
timestamp 1677677812
transform 1 0 1284 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1189
timestamp 1677677812
transform 1 0 1260 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1403
timestamp 1677677812
transform 1 0 1260 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1190
timestamp 1677677812
transform 1 0 1292 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1404
timestamp 1677677812
transform 1 0 1292 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1441
timestamp 1677677812
transform 1 0 1276 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1442
timestamp 1677677812
transform 1 0 1292 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1443
timestamp 1677677812
transform 1 0 1308 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1549
timestamp 1677677812
transform 1 0 1284 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1550
timestamp 1677677812
transform 1 0 1292 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1284
timestamp 1677677812
transform 1 0 1292 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1551
timestamp 1677677812
transform 1 0 1332 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1158
timestamp 1677677812
transform 1 0 1340 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1552
timestamp 1677677812
transform 1 0 1404 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1444
timestamp 1677677812
transform 1 0 1420 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1445
timestamp 1677677812
transform 1 0 1436 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1446
timestamp 1677677812
transform 1 0 1452 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1264
timestamp 1677677812
transform 1 0 1428 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1553
timestamp 1677677812
transform 1 0 1444 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1554
timestamp 1677677812
transform 1 0 1460 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1159
timestamp 1677677812
transform 1 0 1500 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1447
timestamp 1677677812
transform 1 0 1524 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1160
timestamp 1677677812
transform 1 0 1548 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1448
timestamp 1677677812
transform 1 0 1596 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1555
timestamp 1677677812
transform 1 0 1548 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1285
timestamp 1677677812
transform 1 0 1596 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1556
timestamp 1677677812
transform 1 0 1636 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1449
timestamp 1677677812
transform 1 0 1652 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1169
timestamp 1677677812
transform 1 0 1708 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1178
timestamp 1677677812
transform 1 0 1708 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1450
timestamp 1677677812
transform 1 0 1668 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1451
timestamp 1677677812
transform 1 0 1684 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1452
timestamp 1677677812
transform 1 0 1692 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1243
timestamp 1677677812
transform 1 0 1708 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1557
timestamp 1677677812
transform 1 0 1676 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1558
timestamp 1677677812
transform 1 0 1692 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1559
timestamp 1677677812
transform 1 0 1708 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1286
timestamp 1677677812
transform 1 0 1676 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1170
timestamp 1677677812
transform 1 0 1764 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1453
timestamp 1677677812
transform 1 0 1788 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1560
timestamp 1677677812
transform 1 0 1796 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1287
timestamp 1677677812
transform 1 0 1796 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1214
timestamp 1677677812
transform 1 0 1820 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1454
timestamp 1677677812
transform 1 0 1820 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1288
timestamp 1677677812
transform 1 0 1820 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1161
timestamp 1677677812
transform 1 0 1868 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1171
timestamp 1677677812
transform 1 0 1836 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1191
timestamp 1677677812
transform 1 0 1884 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1215
timestamp 1677677812
transform 1 0 1860 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1455
timestamp 1677677812
transform 1 0 1860 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1456
timestamp 1677677812
transform 1 0 1916 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1561
timestamp 1677677812
transform 1 0 1836 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1162
timestamp 1677677812
transform 1 0 1956 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1163
timestamp 1677677812
transform 1 0 2028 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1216
timestamp 1677677812
transform 1 0 2004 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1457
timestamp 1677677812
transform 1 0 1948 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1458
timestamp 1677677812
transform 1 0 2004 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1562
timestamp 1677677812
transform 1 0 2028 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1217
timestamp 1677677812
transform 1 0 2044 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1459
timestamp 1677677812
transform 1 0 2044 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1563
timestamp 1677677812
transform 1 0 2044 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1218
timestamp 1677677812
transform 1 0 2148 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1244
timestamp 1677677812
transform 1 0 2084 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1460
timestamp 1677677812
transform 1 0 2108 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1245
timestamp 1677677812
transform 1 0 2132 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1461
timestamp 1677677812
transform 1 0 2164 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1564
timestamp 1677677812
transform 1 0 2084 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1265
timestamp 1677677812
transform 1 0 2124 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1289
timestamp 1677677812
transform 1 0 2084 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1565
timestamp 1677677812
transform 1 0 2180 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1290
timestamp 1677677812
transform 1 0 2180 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1316
timestamp 1677677812
transform 1 0 2180 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1164
timestamp 1677677812
transform 1 0 2212 0 1 4065
box -3 -3 3 3
use M3_M2  M3_M2_1192
timestamp 1677677812
transform 1 0 2220 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1462
timestamp 1677677812
transform 1 0 2212 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1463
timestamp 1677677812
transform 1 0 2220 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1266
timestamp 1677677812
transform 1 0 2228 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1179
timestamp 1677677812
transform 1 0 2244 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1219
timestamp 1677677812
transform 1 0 2268 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1220
timestamp 1677677812
transform 1 0 2284 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1464
timestamp 1677677812
transform 1 0 2244 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1465
timestamp 1677677812
transform 1 0 2268 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1466
timestamp 1677677812
transform 1 0 2284 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1467
timestamp 1677677812
transform 1 0 2292 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1566
timestamp 1677677812
transform 1 0 2236 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1567
timestamp 1677677812
transform 1 0 2252 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1180
timestamp 1677677812
transform 1 0 2300 0 1 4045
box -3 -3 3 3
use M3_M2  M3_M2_1267
timestamp 1677677812
transform 1 0 2292 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1317
timestamp 1677677812
transform 1 0 2284 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1568
timestamp 1677677812
transform 1 0 2308 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1291
timestamp 1677677812
transform 1 0 2316 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1318
timestamp 1677677812
transform 1 0 2316 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1221
timestamp 1677677812
transform 1 0 2340 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1268
timestamp 1677677812
transform 1 0 2356 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1181
timestamp 1677677812
transform 1 0 2372 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1468
timestamp 1677677812
transform 1 0 2372 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1469
timestamp 1677677812
transform 1 0 2396 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1470
timestamp 1677677812
transform 1 0 2412 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1569
timestamp 1677677812
transform 1 0 2372 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1570
timestamp 1677677812
transform 1 0 2380 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1292
timestamp 1677677812
transform 1 0 2372 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1269
timestamp 1677677812
transform 1 0 2412 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1471
timestamp 1677677812
transform 1 0 2428 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1472
timestamp 1677677812
transform 1 0 2484 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1571
timestamp 1677677812
transform 1 0 2532 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1293
timestamp 1677677812
transform 1 0 2532 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1182
timestamp 1677677812
transform 1 0 2548 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1473
timestamp 1677677812
transform 1 0 2548 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1572
timestamp 1677677812
transform 1 0 2556 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1270
timestamp 1677677812
transform 1 0 2580 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1246
timestamp 1677677812
transform 1 0 2596 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1474
timestamp 1677677812
transform 1 0 2604 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1475
timestamp 1677677812
transform 1 0 2620 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1476
timestamp 1677677812
transform 1 0 2628 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1573
timestamp 1677677812
transform 1 0 2596 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1271
timestamp 1677677812
transform 1 0 2620 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1319
timestamp 1677677812
transform 1 0 2628 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1222
timestamp 1677677812
transform 1 0 2668 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1247
timestamp 1677677812
transform 1 0 2676 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1477
timestamp 1677677812
transform 1 0 2692 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1248
timestamp 1677677812
transform 1 0 2700 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1223
timestamp 1677677812
transform 1 0 2716 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1478
timestamp 1677677812
transform 1 0 2716 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1574
timestamp 1677677812
transform 1 0 2668 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1575
timestamp 1677677812
transform 1 0 2676 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1576
timestamp 1677677812
transform 1 0 2700 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1577
timestamp 1677677812
transform 1 0 2708 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1272
timestamp 1677677812
transform 1 0 2716 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1320
timestamp 1677677812
transform 1 0 2732 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1479
timestamp 1677677812
transform 1 0 2764 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1321
timestamp 1677677812
transform 1 0 2756 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1249
timestamp 1677677812
transform 1 0 2812 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1480
timestamp 1677677812
transform 1 0 2820 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1224
timestamp 1677677812
transform 1 0 2844 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1578
timestamp 1677677812
transform 1 0 2844 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1165
timestamp 1677677812
transform 1 0 2868 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1481
timestamp 1677677812
transform 1 0 2868 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1405
timestamp 1677677812
transform 1 0 2908 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1579
timestamp 1677677812
transform 1 0 2892 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1580
timestamp 1677677812
transform 1 0 2900 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1406
timestamp 1677677812
transform 1 0 2940 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1172
timestamp 1677677812
transform 1 0 2996 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1482
timestamp 1677677812
transform 1 0 2988 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1483
timestamp 1677677812
transform 1 0 3004 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1581
timestamp 1677677812
transform 1 0 3028 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1322
timestamp 1677677812
transform 1 0 3028 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1173
timestamp 1677677812
transform 1 0 3052 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1484
timestamp 1677677812
transform 1 0 3068 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1250
timestamp 1677677812
transform 1 0 3108 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1485
timestamp 1677677812
transform 1 0 3124 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1582
timestamp 1677677812
transform 1 0 3044 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1583
timestamp 1677677812
transform 1 0 3132 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1225
timestamp 1677677812
transform 1 0 3180 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1486
timestamp 1677677812
transform 1 0 3172 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1487
timestamp 1677677812
transform 1 0 3188 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1251
timestamp 1677677812
transform 1 0 3196 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1584
timestamp 1677677812
transform 1 0 3180 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1585
timestamp 1677677812
transform 1 0 3196 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1294
timestamp 1677677812
transform 1 0 3164 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1323
timestamp 1677677812
transform 1 0 3188 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1295
timestamp 1677677812
transform 1 0 3220 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1226
timestamp 1677677812
transform 1 0 3268 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1488
timestamp 1677677812
transform 1 0 3268 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1586
timestamp 1677677812
transform 1 0 3244 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1296
timestamp 1677677812
transform 1 0 3244 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1489
timestamp 1677677812
transform 1 0 3348 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1324
timestamp 1677677812
transform 1 0 3348 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1193
timestamp 1677677812
transform 1 0 3380 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1490
timestamp 1677677812
transform 1 0 3380 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1252
timestamp 1677677812
transform 1 0 3388 0 1 4015
box -3 -3 3 3
use M3_M2  M3_M2_1273
timestamp 1677677812
transform 1 0 3380 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1174
timestamp 1677677812
transform 1 0 3404 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1400
timestamp 1677677812
transform 1 0 3420 0 1 4035
box -2 -2 2 2
use M2_M1  M2_M1_1407
timestamp 1677677812
transform 1 0 3412 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1227
timestamp 1677677812
transform 1 0 3428 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1253
timestamp 1677677812
transform 1 0 3404 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1491
timestamp 1677677812
transform 1 0 3428 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1587
timestamp 1677677812
transform 1 0 3404 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1183
timestamp 1677677812
transform 1 0 3444 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1408
timestamp 1677677812
transform 1 0 3444 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1194
timestamp 1677677812
transform 1 0 3452 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1492
timestamp 1677677812
transform 1 0 3452 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1228
timestamp 1677677812
transform 1 0 3476 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1229
timestamp 1677677812
transform 1 0 3500 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1175
timestamp 1677677812
transform 1 0 3588 0 1 4055
box -3 -3 3 3
use M2_M1  M2_M1_1493
timestamp 1677677812
transform 1 0 3564 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1588
timestamp 1677677812
transform 1 0 3588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1297
timestamp 1677677812
transform 1 0 3564 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1325
timestamp 1677677812
transform 1 0 3588 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1589
timestamp 1677677812
transform 1 0 3604 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1195
timestamp 1677677812
transform 1 0 3644 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1494
timestamp 1677677812
transform 1 0 3644 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1495
timestamp 1677677812
transform 1 0 3660 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1590
timestamp 1677677812
transform 1 0 3636 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1591
timestamp 1677677812
transform 1 0 3652 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1298
timestamp 1677677812
transform 1 0 3652 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1496
timestamp 1677677812
transform 1 0 3676 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1274
timestamp 1677677812
transform 1 0 3676 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1592
timestamp 1677677812
transform 1 0 3692 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1326
timestamp 1677677812
transform 1 0 3700 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1593
timestamp 1677677812
transform 1 0 3740 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1299
timestamp 1677677812
transform 1 0 3740 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1497
timestamp 1677677812
transform 1 0 3788 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1594
timestamp 1677677812
transform 1 0 3764 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1498
timestamp 1677677812
transform 1 0 3868 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1499
timestamp 1677677812
transform 1 0 3876 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1300
timestamp 1677677812
transform 1 0 3876 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1184
timestamp 1677677812
transform 1 0 3908 0 1 4045
box -3 -3 3 3
use M2_M1  M2_M1_1500
timestamp 1677677812
transform 1 0 3924 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1595
timestamp 1677677812
transform 1 0 3916 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1301
timestamp 1677677812
transform 1 0 3924 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1327
timestamp 1677677812
transform 1 0 3916 0 1 3985
box -3 -3 3 3
use M3_M2  M3_M2_1254
timestamp 1677677812
transform 1 0 3972 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1596
timestamp 1677677812
transform 1 0 3972 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1176
timestamp 1677677812
transform 1 0 4052 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1177
timestamp 1677677812
transform 1 0 4076 0 1 4055
box -3 -3 3 3
use M3_M2  M3_M2_1196
timestamp 1677677812
transform 1 0 3988 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1197
timestamp 1677677812
transform 1 0 4020 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1501
timestamp 1677677812
transform 1 0 4020 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1255
timestamp 1677677812
transform 1 0 4044 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1502
timestamp 1677677812
transform 1 0 4076 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1597
timestamp 1677677812
transform 1 0 3996 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1328
timestamp 1677677812
transform 1 0 3996 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1503
timestamp 1677677812
transform 1 0 4156 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1230
timestamp 1677677812
transform 1 0 4212 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1256
timestamp 1677677812
transform 1 0 4204 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1598
timestamp 1677677812
transform 1 0 4108 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1275
timestamp 1677677812
transform 1 0 4196 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1302
timestamp 1677677812
transform 1 0 4156 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1599
timestamp 1677677812
transform 1 0 4212 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1231
timestamp 1677677812
transform 1 0 4228 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1232
timestamp 1677677812
transform 1 0 4260 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1504
timestamp 1677677812
transform 1 0 4228 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1505
timestamp 1677677812
transform 1 0 4236 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1506
timestamp 1677677812
transform 1 0 4244 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1257
timestamp 1677677812
transform 1 0 4252 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1507
timestamp 1677677812
transform 1 0 4260 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1600
timestamp 1677677812
transform 1 0 4252 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1601
timestamp 1677677812
transform 1 0 4268 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1303
timestamp 1677677812
transform 1 0 4252 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1233
timestamp 1677677812
transform 1 0 4284 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1602
timestamp 1677677812
transform 1 0 4284 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1198
timestamp 1677677812
transform 1 0 4316 0 1 4035
box -3 -3 3 3
use M2_M1  M2_M1_1508
timestamp 1677677812
transform 1 0 4300 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1509
timestamp 1677677812
transform 1 0 4316 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1510
timestamp 1677677812
transform 1 0 4332 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1409
timestamp 1677677812
transform 1 0 4356 0 1 4025
box -2 -2 2 2
use M3_M2  M3_M2_1258
timestamp 1677677812
transform 1 0 4356 0 1 4015
box -3 -3 3 3
use M2_M1  M2_M1_1603
timestamp 1677677812
transform 1 0 4356 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1166
timestamp 1677677812
transform 1 0 4372 0 1 4065
box -3 -3 3 3
use M2_M1  M2_M1_1401
timestamp 1677677812
transform 1 0 4372 0 1 4035
box -2 -2 2 2
use M3_M2  M3_M2_1199
timestamp 1677677812
transform 1 0 4380 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1234
timestamp 1677677812
transform 1 0 4372 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1410
timestamp 1677677812
transform 1 0 4380 0 1 4025
box -2 -2 2 2
use M2_M1  M2_M1_1511
timestamp 1677677812
transform 1 0 4380 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1276
timestamp 1677677812
transform 1 0 4380 0 1 4005
box -3 -3 3 3
use M3_M2  M3_M2_1235
timestamp 1677677812
transform 1 0 4404 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1512
timestamp 1677677812
transform 1 0 4396 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1236
timestamp 1677677812
transform 1 0 4452 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1604
timestamp 1677677812
transform 1 0 4452 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1200
timestamp 1677677812
transform 1 0 4580 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1237
timestamp 1677677812
transform 1 0 4516 0 1 4025
box -3 -3 3 3
use M3_M2  M3_M2_1238
timestamp 1677677812
transform 1 0 4556 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1513
timestamp 1677677812
transform 1 0 4516 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1514
timestamp 1677677812
transform 1 0 4556 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1515
timestamp 1677677812
transform 1 0 4564 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1516
timestamp 1677677812
transform 1 0 4580 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1517
timestamp 1677677812
transform 1 0 4596 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1605
timestamp 1677677812
transform 1 0 4468 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1606
timestamp 1677677812
transform 1 0 4556 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1607
timestamp 1677677812
transform 1 0 4572 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1608
timestamp 1677677812
transform 1 0 4588 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1304
timestamp 1677677812
transform 1 0 4516 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1305
timestamp 1677677812
transform 1 0 4572 0 1 3995
box -3 -3 3 3
use M2_M1  M2_M1_1609
timestamp 1677677812
transform 1 0 4604 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1518
timestamp 1677677812
transform 1 0 4612 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1610
timestamp 1677677812
transform 1 0 4612 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1201
timestamp 1677677812
transform 1 0 4668 0 1 4035
box -3 -3 3 3
use M3_M2  M3_M2_1239
timestamp 1677677812
transform 1 0 4660 0 1 4025
box -3 -3 3 3
use M2_M1  M2_M1_1519
timestamp 1677677812
transform 1 0 4636 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1520
timestamp 1677677812
transform 1 0 4652 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1521
timestamp 1677677812
transform 1 0 4668 0 1 4015
box -2 -2 2 2
use M2_M1  M2_M1_1522
timestamp 1677677812
transform 1 0 4676 0 1 4015
box -2 -2 2 2
use M3_M2  M3_M2_1277
timestamp 1677677812
transform 1 0 4636 0 1 4005
box -3 -3 3 3
use M2_M1  M2_M1_1611
timestamp 1677677812
transform 1 0 4652 0 1 4005
box -2 -2 2 2
use M2_M1  M2_M1_1612
timestamp 1677677812
transform 1 0 4660 0 1 4005
box -2 -2 2 2
use M3_M2  M3_M2_1306
timestamp 1677677812
transform 1 0 4652 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1307
timestamp 1677677812
transform 1 0 4676 0 1 3995
box -3 -3 3 3
use M3_M2  M3_M2_1329
timestamp 1677677812
transform 1 0 4700 0 1 3985
box -3 -3 3 3
use M2_M1  M2_M1_1613
timestamp 1677677812
transform 1 0 4780 0 1 4005
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_14
timestamp 1677677812
transform 1 0 48 0 1 3970
box -10 -3 10 3
use M3_M2  M3_M2_1330
timestamp 1677677812
transform 1 0 148 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_97
timestamp 1677677812
transform 1 0 72 0 1 3970
box -8 -3 104 105
use FILL  FILL_1267
timestamp 1677677812
transform 1 0 168 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1331
timestamp 1677677812
transform 1 0 188 0 1 3975
box -3 -3 3 3
use FILL  FILL_1268
timestamp 1677677812
transform 1 0 176 0 1 3970
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1677677812
transform 1 0 184 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_64
timestamp 1677677812
transform 1 0 192 0 1 3970
box -8 -3 46 105
use FILL  FILL_1270
timestamp 1677677812
transform 1 0 232 0 1 3970
box -8 -3 16 105
use FILL  FILL_1271
timestamp 1677677812
transform 1 0 240 0 1 3970
box -8 -3 16 105
use FILL  FILL_1272
timestamp 1677677812
transform 1 0 248 0 1 3970
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1677677812
transform 1 0 256 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_65
timestamp 1677677812
transform 1 0 264 0 1 3970
box -8 -3 46 105
use FILL  FILL_1274
timestamp 1677677812
transform 1 0 304 0 1 3970
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1677677812
transform 1 0 312 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_98
timestamp 1677677812
transform -1 0 416 0 1 3970
box -8 -3 104 105
use FILL  FILL_1276
timestamp 1677677812
transform 1 0 416 0 1 3970
box -8 -3 16 105
use FILL  FILL_1277
timestamp 1677677812
transform 1 0 424 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_99
timestamp 1677677812
transform 1 0 432 0 1 3970
box -8 -3 104 105
use FILL  FILL_1278
timestamp 1677677812
transform 1 0 528 0 1 3970
box -8 -3 16 105
use FILL  FILL_1287
timestamp 1677677812
transform 1 0 536 0 1 3970
box -8 -3 16 105
use FILL  FILL_1289
timestamp 1677677812
transform 1 0 544 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_67
timestamp 1677677812
transform -1 0 592 0 1 3970
box -8 -3 46 105
use FILL  FILL_1290
timestamp 1677677812
transform 1 0 592 0 1 3970
box -8 -3 16 105
use FILL  FILL_1291
timestamp 1677677812
transform 1 0 600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1295
timestamp 1677677812
transform 1 0 608 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_68
timestamp 1677677812
transform 1 0 616 0 1 3970
box -8 -3 46 105
use FILL  FILL_1297
timestamp 1677677812
transform 1 0 656 0 1 3970
box -8 -3 16 105
use FILL  FILL_1298
timestamp 1677677812
transform 1 0 664 0 1 3970
box -8 -3 16 105
use FILL  FILL_1299
timestamp 1677677812
transform 1 0 672 0 1 3970
box -8 -3 16 105
use FILL  FILL_1300
timestamp 1677677812
transform 1 0 680 0 1 3970
box -8 -3 16 105
use FILL  FILL_1305
timestamp 1677677812
transform 1 0 688 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_67
timestamp 1677677812
transform -1 0 736 0 1 3970
box -8 -3 46 105
use FILL  FILL_1306
timestamp 1677677812
transform 1 0 736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1312
timestamp 1677677812
transform 1 0 744 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_123
timestamp 1677677812
transform 1 0 752 0 1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_103
timestamp 1677677812
transform 1 0 768 0 1 3970
box -8 -3 104 105
use FILL  FILL_1313
timestamp 1677677812
transform 1 0 864 0 1 3970
box -8 -3 16 105
use NOR2X1  NOR2X1_17
timestamp 1677677812
transform 1 0 872 0 1 3970
box -8 -3 32 105
use FILL  FILL_1314
timestamp 1677677812
transform 1 0 896 0 1 3970
box -8 -3 16 105
use FILL  FILL_1321
timestamp 1677677812
transform 1 0 904 0 1 3970
box -8 -3 16 105
use FILL  FILL_1323
timestamp 1677677812
transform 1 0 912 0 1 3970
box -8 -3 16 105
use FILL  FILL_1325
timestamp 1677677812
transform 1 0 920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1327
timestamp 1677677812
transform 1 0 928 0 1 3970
box -8 -3 16 105
use FILL  FILL_1328
timestamp 1677677812
transform 1 0 936 0 1 3970
box -8 -3 16 105
use FILL  FILL_1329
timestamp 1677677812
transform 1 0 944 0 1 3970
box -8 -3 16 105
use FILL  FILL_1330
timestamp 1677677812
transform 1 0 952 0 1 3970
box -8 -3 16 105
use FILL  FILL_1331
timestamp 1677677812
transform 1 0 960 0 1 3970
box -8 -3 16 105
use FILL  FILL_1332
timestamp 1677677812
transform 1 0 968 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_125
timestamp 1677677812
transform 1 0 976 0 1 3970
box -9 -3 26 105
use FILL  FILL_1334
timestamp 1677677812
transform 1 0 992 0 1 3970
box -8 -3 16 105
use FILL  FILL_1338
timestamp 1677677812
transform 1 0 1000 0 1 3970
box -8 -3 16 105
use FILL  FILL_1339
timestamp 1677677812
transform 1 0 1008 0 1 3970
box -8 -3 16 105
use FILL  FILL_1340
timestamp 1677677812
transform 1 0 1016 0 1 3970
box -8 -3 16 105
use FILL  FILL_1341
timestamp 1677677812
transform 1 0 1024 0 1 3970
box -8 -3 16 105
use FILL  FILL_1342
timestamp 1677677812
transform 1 0 1032 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_71
timestamp 1677677812
transform 1 0 1040 0 1 3970
box -8 -3 46 105
use FILL  FILL_1343
timestamp 1677677812
transform 1 0 1080 0 1 3970
box -8 -3 16 105
use FILL  FILL_1344
timestamp 1677677812
transform 1 0 1088 0 1 3970
box -8 -3 16 105
use FILL  FILL_1345
timestamp 1677677812
transform 1 0 1096 0 1 3970
box -8 -3 16 105
use FILL  FILL_1347
timestamp 1677677812
transform 1 0 1104 0 1 3970
box -8 -3 16 105
use FILL  FILL_1349
timestamp 1677677812
transform 1 0 1112 0 1 3970
box -8 -3 16 105
use FILL  FILL_1351
timestamp 1677677812
transform 1 0 1120 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_72
timestamp 1677677812
transform 1 0 1128 0 1 3970
box -8 -3 46 105
use FILL  FILL_1353
timestamp 1677677812
transform 1 0 1168 0 1 3970
box -8 -3 16 105
use FILL  FILL_1354
timestamp 1677677812
transform 1 0 1176 0 1 3970
box -8 -3 16 105
use FILL  FILL_1355
timestamp 1677677812
transform 1 0 1184 0 1 3970
box -8 -3 16 105
use FILL  FILL_1356
timestamp 1677677812
transform 1 0 1192 0 1 3970
box -8 -3 16 105
use FILL  FILL_1357
timestamp 1677677812
transform 1 0 1200 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_34
timestamp 1677677812
transform 1 0 1208 0 1 3970
box -8 -3 34 105
use FILL  FILL_1358
timestamp 1677677812
transform 1 0 1240 0 1 3970
box -8 -3 16 105
use FILL  FILL_1362
timestamp 1677677812
transform 1 0 1248 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_35
timestamp 1677677812
transform -1 0 1288 0 1 3970
box -8 -3 34 105
use OAI21X1  OAI21X1_36
timestamp 1677677812
transform -1 0 1320 0 1 3970
box -8 -3 34 105
use FILL  FILL_1364
timestamp 1677677812
transform 1 0 1320 0 1 3970
box -8 -3 16 105
use FILL  FILL_1365
timestamp 1677677812
transform 1 0 1328 0 1 3970
box -8 -3 16 105
use FILL  FILL_1366
timestamp 1677677812
transform 1 0 1336 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_126
timestamp 1677677812
transform 1 0 1344 0 1 3970
box -9 -3 26 105
use FILL  FILL_1367
timestamp 1677677812
transform 1 0 1360 0 1 3970
box -8 -3 16 105
use FILL  FILL_1368
timestamp 1677677812
transform 1 0 1368 0 1 3970
box -8 -3 16 105
use FILL  FILL_1369
timestamp 1677677812
transform 1 0 1376 0 1 3970
box -8 -3 16 105
use FILL  FILL_1370
timestamp 1677677812
transform 1 0 1384 0 1 3970
box -8 -3 16 105
use FILL  FILL_1371
timestamp 1677677812
transform 1 0 1392 0 1 3970
box -8 -3 16 105
use FILL  FILL_1372
timestamp 1677677812
transform 1 0 1400 0 1 3970
box -8 -3 16 105
use FILL  FILL_1373
timestamp 1677677812
transform 1 0 1408 0 1 3970
box -8 -3 16 105
use FILL  FILL_1374
timestamp 1677677812
transform 1 0 1416 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1332
timestamp 1677677812
transform 1 0 1460 0 1 3975
box -3 -3 3 3
use OAI22X1  OAI22X1_68
timestamp 1677677812
transform -1 0 1464 0 1 3970
box -8 -3 46 105
use FILL  FILL_1375
timestamp 1677677812
transform 1 0 1464 0 1 3970
box -8 -3 16 105
use FILL  FILL_1387
timestamp 1677677812
transform 1 0 1472 0 1 3970
box -8 -3 16 105
use FILL  FILL_1388
timestamp 1677677812
transform 1 0 1480 0 1 3970
box -8 -3 16 105
use FILL  FILL_1389
timestamp 1677677812
transform 1 0 1488 0 1 3970
box -8 -3 16 105
use FILL  FILL_1391
timestamp 1677677812
transform 1 0 1496 0 1 3970
box -8 -3 16 105
use FILL  FILL_1393
timestamp 1677677812
transform 1 0 1504 0 1 3970
box -8 -3 16 105
use FILL  FILL_1395
timestamp 1677677812
transform 1 0 1512 0 1 3970
box -8 -3 16 105
use FILL  FILL_1397
timestamp 1677677812
transform 1 0 1520 0 1 3970
box -8 -3 16 105
use FILL  FILL_1399
timestamp 1677677812
transform 1 0 1528 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_108
timestamp 1677677812
transform 1 0 1536 0 1 3970
box -8 -3 104 105
use FILL  FILL_1401
timestamp 1677677812
transform 1 0 1632 0 1 3970
box -8 -3 16 105
use FILL  FILL_1403
timestamp 1677677812
transform 1 0 1640 0 1 3970
box -8 -3 16 105
use FILL  FILL_1405
timestamp 1677677812
transform 1 0 1648 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_69
timestamp 1677677812
transform -1 0 1696 0 1 3970
box -8 -3 46 105
use INVX2  INVX2_128
timestamp 1677677812
transform -1 0 1712 0 1 3970
box -9 -3 26 105
use FILL  FILL_1406
timestamp 1677677812
transform 1 0 1712 0 1 3970
box -8 -3 16 105
use FILL  FILL_1412
timestamp 1677677812
transform 1 0 1720 0 1 3970
box -8 -3 16 105
use FILL  FILL_1414
timestamp 1677677812
transform 1 0 1728 0 1 3970
box -8 -3 16 105
use FILL  FILL_1416
timestamp 1677677812
transform 1 0 1736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1418
timestamp 1677677812
transform 1 0 1744 0 1 3970
box -8 -3 16 105
use FILL  FILL_1420
timestamp 1677677812
transform 1 0 1752 0 1 3970
box -8 -3 16 105
use FILL  FILL_1422
timestamp 1677677812
transform 1 0 1760 0 1 3970
box -8 -3 16 105
use FILL  FILL_1424
timestamp 1677677812
transform 1 0 1768 0 1 3970
box -8 -3 16 105
use FILL  FILL_1426
timestamp 1677677812
transform 1 0 1776 0 1 3970
box -8 -3 16 105
use FILL  FILL_1428
timestamp 1677677812
transform 1 0 1784 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_131
timestamp 1677677812
transform 1 0 1792 0 1 3970
box -9 -3 26 105
use FILL  FILL_1430
timestamp 1677677812
transform 1 0 1808 0 1 3970
box -8 -3 16 105
use FILL  FILL_1431
timestamp 1677677812
transform 1 0 1816 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_110
timestamp 1677677812
transform 1 0 1824 0 1 3970
box -8 -3 104 105
use FILL  FILL_1432
timestamp 1677677812
transform 1 0 1920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1433
timestamp 1677677812
transform 1 0 1928 0 1 3970
box -8 -3 16 105
use FILL  FILL_1434
timestamp 1677677812
transform 1 0 1936 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_111
timestamp 1677677812
transform -1 0 2040 0 1 3970
box -8 -3 104 105
use FILL  FILL_1435
timestamp 1677677812
transform 1 0 2040 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_132
timestamp 1677677812
transform 1 0 2048 0 1 3970
box -9 -3 26 105
use FILL  FILL_1453
timestamp 1677677812
transform 1 0 2064 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_112
timestamp 1677677812
transform 1 0 2072 0 1 3970
box -8 -3 104 105
use FILL  FILL_1457
timestamp 1677677812
transform 1 0 2168 0 1 3970
box -8 -3 16 105
use FILL  FILL_1458
timestamp 1677677812
transform 1 0 2176 0 1 3970
box -8 -3 16 105
use FILL  FILL_1466
timestamp 1677677812
transform 1 0 2184 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_3
timestamp 1677677812
transform -1 0 2216 0 1 3970
box -5 -3 28 105
use BUFX2  BUFX2_4
timestamp 1677677812
transform 1 0 2216 0 1 3970
box -5 -3 28 105
use FILL  FILL_1467
timestamp 1677677812
transform 1 0 2240 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_76
timestamp 1677677812
transform 1 0 2248 0 1 3970
box -8 -3 46 105
use FILL  FILL_1473
timestamp 1677677812
transform 1 0 2288 0 1 3970
box -8 -3 16 105
use FILL  FILL_1474
timestamp 1677677812
transform 1 0 2296 0 1 3970
box -8 -3 16 105
use FILL  FILL_1477
timestamp 1677677812
transform 1 0 2304 0 1 3970
box -8 -3 16 105
use FILL  FILL_1479
timestamp 1677677812
transform 1 0 2312 0 1 3970
box -8 -3 16 105
use FILL  FILL_1480
timestamp 1677677812
transform 1 0 2320 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_6
timestamp 1677677812
transform 1 0 2328 0 1 3970
box -5 -3 28 105
use FILL  FILL_1481
timestamp 1677677812
transform 1 0 2352 0 1 3970
box -8 -3 16 105
use FILL  FILL_1483
timestamp 1677677812
transform 1 0 2360 0 1 3970
box -8 -3 16 105
use FILL  FILL_1485
timestamp 1677677812
transform 1 0 2368 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_78
timestamp 1677677812
transform 1 0 2376 0 1 3970
box -8 -3 46 105
use FILL  FILL_1487
timestamp 1677677812
transform 1 0 2416 0 1 3970
box -8 -3 16 105
use FILL  FILL_1492
timestamp 1677677812
transform 1 0 2424 0 1 3970
box -8 -3 16 105
use FILL  FILL_1494
timestamp 1677677812
transform 1 0 2432 0 1 3970
box -8 -3 16 105
use FILL  FILL_1496
timestamp 1677677812
transform 1 0 2440 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_113
timestamp 1677677812
transform -1 0 2544 0 1 3970
box -8 -3 104 105
use FILL  FILL_1497
timestamp 1677677812
transform 1 0 2544 0 1 3970
box -8 -3 16 105
use FILL  FILL_1498
timestamp 1677677812
transform 1 0 2552 0 1 3970
box -8 -3 16 105
use FILL  FILL_1499
timestamp 1677677812
transform 1 0 2560 0 1 3970
box -8 -3 16 105
use FILL  FILL_1500
timestamp 1677677812
transform 1 0 2568 0 1 3970
box -8 -3 16 105
use FILL  FILL_1501
timestamp 1677677812
transform 1 0 2576 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_79
timestamp 1677677812
transform 1 0 2584 0 1 3970
box -8 -3 46 105
use FILL  FILL_1502
timestamp 1677677812
transform 1 0 2624 0 1 3970
box -8 -3 16 105
use FILL  FILL_1503
timestamp 1677677812
transform 1 0 2632 0 1 3970
box -8 -3 16 105
use FILL  FILL_1504
timestamp 1677677812
transform 1 0 2640 0 1 3970
box -8 -3 16 105
use FILL  FILL_1505
timestamp 1677677812
transform 1 0 2648 0 1 3970
box -8 -3 16 105
use FILL  FILL_1506
timestamp 1677677812
transform 1 0 2656 0 1 3970
box -8 -3 16 105
use FILL  FILL_1507
timestamp 1677677812
transform 1 0 2664 0 1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_80
timestamp 1677677812
transform 1 0 2672 0 1 3970
box -8 -3 46 105
use FILL  FILL_1508
timestamp 1677677812
transform 1 0 2712 0 1 3970
box -8 -3 16 105
use FILL  FILL_1523
timestamp 1677677812
transform 1 0 2720 0 1 3970
box -8 -3 16 105
use FILL  FILL_1524
timestamp 1677677812
transform 1 0 2728 0 1 3970
box -8 -3 16 105
use FILL  FILL_1525
timestamp 1677677812
transform 1 0 2736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1526
timestamp 1677677812
transform 1 0 2744 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_137
timestamp 1677677812
transform 1 0 2752 0 1 3970
box -9 -3 26 105
use FILL  FILL_1527
timestamp 1677677812
transform 1 0 2768 0 1 3970
box -8 -3 16 105
use FILL  FILL_1528
timestamp 1677677812
transform 1 0 2776 0 1 3970
box -8 -3 16 105
use FILL  FILL_1529
timestamp 1677677812
transform 1 0 2784 0 1 3970
box -8 -3 16 105
use FILL  FILL_1530
timestamp 1677677812
transform 1 0 2792 0 1 3970
box -8 -3 16 105
use FILL  FILL_1531
timestamp 1677677812
transform 1 0 2800 0 1 3970
box -8 -3 16 105
use FILL  FILL_1532
timestamp 1677677812
transform 1 0 2808 0 1 3970
box -8 -3 16 105
use FILL  FILL_1533
timestamp 1677677812
transform 1 0 2816 0 1 3970
box -8 -3 16 105
use FILL  FILL_1535
timestamp 1677677812
transform 1 0 2824 0 1 3970
box -8 -3 16 105
use FILL  FILL_1537
timestamp 1677677812
transform 1 0 2832 0 1 3970
box -8 -3 16 105
use FILL  FILL_1539
timestamp 1677677812
transform 1 0 2840 0 1 3970
box -8 -3 16 105
use FILL  FILL_1540
timestamp 1677677812
transform 1 0 2848 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_38
timestamp 1677677812
transform 1 0 2856 0 1 3970
box -8 -3 34 105
use FILL  FILL_1541
timestamp 1677677812
transform 1 0 2888 0 1 3970
box -8 -3 16 105
use FILL  FILL_1545
timestamp 1677677812
transform 1 0 2896 0 1 3970
box -8 -3 16 105
use FILL  FILL_1547
timestamp 1677677812
transform 1 0 2904 0 1 3970
box -8 -3 16 105
use FILL  FILL_1548
timestamp 1677677812
transform 1 0 2912 0 1 3970
box -8 -3 16 105
use FILL  FILL_1549
timestamp 1677677812
transform 1 0 2920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1550
timestamp 1677677812
transform 1 0 2928 0 1 3970
box -8 -3 16 105
use FILL  FILL_1552
timestamp 1677677812
transform 1 0 2936 0 1 3970
box -8 -3 16 105
use FILL  FILL_1554
timestamp 1677677812
transform 1 0 2944 0 1 3970
box -8 -3 16 105
use FILL  FILL_1556
timestamp 1677677812
transform 1 0 2952 0 1 3970
box -8 -3 16 105
use FILL  FILL_1557
timestamp 1677677812
transform 1 0 2960 0 1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_40
timestamp 1677677812
transform -1 0 3000 0 1 3970
box -8 -3 34 105
use FILL  FILL_1558
timestamp 1677677812
transform 1 0 3000 0 1 3970
box -8 -3 16 105
use FILL  FILL_1559
timestamp 1677677812
transform 1 0 3008 0 1 3970
box -8 -3 16 105
use FILL  FILL_1560
timestamp 1677677812
transform 1 0 3016 0 1 3970
box -8 -3 16 105
use FILL  FILL_1561
timestamp 1677677812
transform 1 0 3024 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1333
timestamp 1677677812
transform 1 0 3092 0 1 3975
box -3 -3 3 3
use M3_M2  M3_M2_1334
timestamp 1677677812
transform 1 0 3132 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_116
timestamp 1677677812
transform 1 0 3032 0 1 3970
box -8 -3 104 105
use FILL  FILL_1562
timestamp 1677677812
transform 1 0 3128 0 1 3970
box -8 -3 16 105
use FILL  FILL_1563
timestamp 1677677812
transform 1 0 3136 0 1 3970
box -8 -3 16 105
use FILL  FILL_1564
timestamp 1677677812
transform 1 0 3144 0 1 3970
box -8 -3 16 105
use FILL  FILL_1565
timestamp 1677677812
transform 1 0 3152 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_72
timestamp 1677677812
transform 1 0 3160 0 1 3970
box -8 -3 46 105
use FILL  FILL_1566
timestamp 1677677812
transform 1 0 3200 0 1 3970
box -8 -3 16 105
use FILL  FILL_1580
timestamp 1677677812
transform 1 0 3208 0 1 3970
box -8 -3 16 105
use FILL  FILL_1581
timestamp 1677677812
transform 1 0 3216 0 1 3970
box -8 -3 16 105
use FILL  FILL_1582
timestamp 1677677812
transform 1 0 3224 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_118
timestamp 1677677812
transform 1 0 3232 0 1 3970
box -8 -3 104 105
use FILL  FILL_1583
timestamp 1677677812
transform 1 0 3328 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_139
timestamp 1677677812
transform 1 0 3336 0 1 3970
box -9 -3 26 105
use FILL  FILL_1584
timestamp 1677677812
transform 1 0 3352 0 1 3970
box -8 -3 16 105
use FILL  FILL_1585
timestamp 1677677812
transform 1 0 3360 0 1 3970
box -8 -3 16 105
use FILL  FILL_1586
timestamp 1677677812
transform 1 0 3368 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_7
timestamp 1677677812
transform 1 0 3376 0 1 3970
box -5 -3 28 105
use FILL  FILL_1587
timestamp 1677677812
transform 1 0 3400 0 1 3970
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1677677812
transform -1 0 3440 0 1 3970
box -8 -3 40 105
use FILL  FILL_1588
timestamp 1677677812
transform 1 0 3440 0 1 3970
box -8 -3 16 105
use FILL  FILL_1595
timestamp 1677677812
transform 1 0 3448 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_140
timestamp 1677677812
transform -1 0 3472 0 1 3970
box -9 -3 26 105
use FILL  FILL_1596
timestamp 1677677812
transform 1 0 3472 0 1 3970
box -8 -3 16 105
use FILL  FILL_1597
timestamp 1677677812
transform 1 0 3480 0 1 3970
box -8 -3 16 105
use FILL  FILL_1598
timestamp 1677677812
transform 1 0 3488 0 1 3970
box -8 -3 16 105
use FILL  FILL_1599
timestamp 1677677812
transform 1 0 3496 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_121
timestamp 1677677812
transform -1 0 3600 0 1 3970
box -8 -3 104 105
use FILL  FILL_1600
timestamp 1677677812
transform 1 0 3600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1601
timestamp 1677677812
transform 1 0 3608 0 1 3970
box -8 -3 16 105
use FILL  FILL_1602
timestamp 1677677812
transform 1 0 3616 0 1 3970
box -8 -3 16 105
use FILL  FILL_1603
timestamp 1677677812
transform 1 0 3624 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_74
timestamp 1677677812
transform -1 0 3672 0 1 3970
box -8 -3 46 105
use FILL  FILL_1604
timestamp 1677677812
transform 1 0 3672 0 1 3970
box -8 -3 16 105
use FILL  FILL_1605
timestamp 1677677812
transform 1 0 3680 0 1 3970
box -8 -3 16 105
use FILL  FILL_1606
timestamp 1677677812
transform 1 0 3688 0 1 3970
box -8 -3 16 105
use FILL  FILL_1607
timestamp 1677677812
transform 1 0 3696 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_8
timestamp 1677677812
transform 1 0 3704 0 1 3970
box -5 -3 28 105
use FILL  FILL_1608
timestamp 1677677812
transform 1 0 3728 0 1 3970
box -8 -3 16 105
use FILL  FILL_1609
timestamp 1677677812
transform 1 0 3736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1622
timestamp 1677677812
transform 1 0 3744 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_123
timestamp 1677677812
transform 1 0 3752 0 1 3970
box -8 -3 104 105
use FILL  FILL_1624
timestamp 1677677812
transform 1 0 3848 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_141
timestamp 1677677812
transform 1 0 3856 0 1 3970
box -9 -3 26 105
use FILL  FILL_1625
timestamp 1677677812
transform 1 0 3872 0 1 3970
box -8 -3 16 105
use FILL  FILL_1626
timestamp 1677677812
transform 1 0 3880 0 1 3970
box -8 -3 16 105
use FILL  FILL_1639
timestamp 1677677812
transform 1 0 3888 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_10
timestamp 1677677812
transform 1 0 3896 0 1 3970
box -5 -3 28 105
use FILL  FILL_1641
timestamp 1677677812
transform 1 0 3920 0 1 3970
box -8 -3 16 105
use FILL  FILL_1642
timestamp 1677677812
transform 1 0 3928 0 1 3970
box -8 -3 16 105
use BUFX2  BUFX2_11
timestamp 1677677812
transform 1 0 3936 0 1 3970
box -5 -3 28 105
use FILL  FILL_1643
timestamp 1677677812
transform 1 0 3960 0 1 3970
box -8 -3 16 105
use FILL  FILL_1644
timestamp 1677677812
transform 1 0 3968 0 1 3970
box -8 -3 16 105
use FILL  FILL_1645
timestamp 1677677812
transform 1 0 3976 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1335
timestamp 1677677812
transform 1 0 4052 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_124
timestamp 1677677812
transform 1 0 3984 0 1 3970
box -8 -3 104 105
use FILL  FILL_1646
timestamp 1677677812
transform 1 0 4080 0 1 3970
box -8 -3 16 105
use FILL  FILL_1647
timestamp 1677677812
transform 1 0 4088 0 1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_125
timestamp 1677677812
transform 1 0 4096 0 1 3970
box -8 -3 104 105
use M3_M2  M3_M2_1336
timestamp 1677677812
transform 1 0 4212 0 1 3975
box -3 -3 3 3
use INVX2  INVX2_142
timestamp 1677677812
transform 1 0 4192 0 1 3970
box -9 -3 26 105
use FILL  FILL_1648
timestamp 1677677812
transform 1 0 4208 0 1 3970
box -8 -3 16 105
use FILL  FILL_1649
timestamp 1677677812
transform 1 0 4216 0 1 3970
box -8 -3 16 105
use FILL  FILL_1655
timestamp 1677677812
transform 1 0 4224 0 1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_78
timestamp 1677677812
transform 1 0 4232 0 1 3970
box -8 -3 46 105
use FILL  FILL_1657
timestamp 1677677812
transform 1 0 4272 0 1 3970
box -8 -3 16 105
use FILL  FILL_1659
timestamp 1677677812
transform 1 0 4280 0 1 3970
box -8 -3 16 105
use FILL  FILL_1660
timestamp 1677677812
transform 1 0 4288 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1337
timestamp 1677677812
transform 1 0 4316 0 1 3975
box -3 -3 3 3
use AOI22X1  AOI22X1_82
timestamp 1677677812
transform -1 0 4336 0 1 3970
box -8 -3 46 105
use FILL  FILL_1661
timestamp 1677677812
transform 1 0 4336 0 1 3970
box -8 -3 16 105
use FILL  FILL_1662
timestamp 1677677812
transform 1 0 4344 0 1 3970
box -8 -3 16 105
use FILL  FILL_1663
timestamp 1677677812
transform 1 0 4352 0 1 3970
box -8 -3 16 105
use NAND3X1  NAND3X1_8
timestamp 1677677812
transform -1 0 4392 0 1 3970
box -8 -3 40 105
use FILL  FILL_1664
timestamp 1677677812
transform 1 0 4392 0 1 3970
box -8 -3 16 105
use FILL  FILL_1665
timestamp 1677677812
transform 1 0 4400 0 1 3970
box -8 -3 16 105
use FILL  FILL_1666
timestamp 1677677812
transform 1 0 4408 0 1 3970
box -8 -3 16 105
use FILL  FILL_1667
timestamp 1677677812
transform 1 0 4416 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_143
timestamp 1677677812
transform -1 0 4440 0 1 3970
box -9 -3 26 105
use FILL  FILL_1668
timestamp 1677677812
transform 1 0 4440 0 1 3970
box -8 -3 16 105
use FILL  FILL_1669
timestamp 1677677812
transform 1 0 4448 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1338
timestamp 1677677812
transform 1 0 4500 0 1 3975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_129
timestamp 1677677812
transform 1 0 4456 0 1 3970
box -8 -3 104 105
use OAI22X1  OAI22X1_80
timestamp 1677677812
transform 1 0 4552 0 1 3970
box -8 -3 46 105
use FILL  FILL_1670
timestamp 1677677812
transform 1 0 4592 0 1 3970
box -8 -3 16 105
use FILL  FILL_1685
timestamp 1677677812
transform 1 0 4600 0 1 3970
box -8 -3 16 105
use FILL  FILL_1686
timestamp 1677677812
transform 1 0 4608 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1339
timestamp 1677677812
transform 1 0 4636 0 1 3975
box -3 -3 3 3
use AOI22X1  AOI22X1_83
timestamp 1677677812
transform -1 0 4656 0 1 3970
box -8 -3 46 105
use INVX2  INVX2_146
timestamp 1677677812
transform 1 0 4656 0 1 3970
box -9 -3 26 105
use FILL  FILL_1687
timestamp 1677677812
transform 1 0 4672 0 1 3970
box -8 -3 16 105
use FILL  FILL_1691
timestamp 1677677812
transform 1 0 4680 0 1 3970
box -8 -3 16 105
use FILL  FILL_1693
timestamp 1677677812
transform 1 0 4688 0 1 3970
box -8 -3 16 105
use FILL  FILL_1694
timestamp 1677677812
transform 1 0 4696 0 1 3970
box -8 -3 16 105
use FILL  FILL_1695
timestamp 1677677812
transform 1 0 4704 0 1 3970
box -8 -3 16 105
use INVX2  INVX2_148
timestamp 1677677812
transform -1 0 4728 0 1 3970
box -9 -3 26 105
use FILL  FILL_1696
timestamp 1677677812
transform 1 0 4728 0 1 3970
box -8 -3 16 105
use FILL  FILL_1697
timestamp 1677677812
transform 1 0 4736 0 1 3970
box -8 -3 16 105
use FILL  FILL_1698
timestamp 1677677812
transform 1 0 4744 0 1 3970
box -8 -3 16 105
use FILL  FILL_1699
timestamp 1677677812
transform 1 0 4752 0 1 3970
box -8 -3 16 105
use FILL  FILL_1700
timestamp 1677677812
transform 1 0 4760 0 1 3970
box -8 -3 16 105
use FILL  FILL_1701
timestamp 1677677812
transform 1 0 4768 0 1 3970
box -8 -3 16 105
use FILL  FILL_1702
timestamp 1677677812
transform 1 0 4776 0 1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1340
timestamp 1677677812
transform 1 0 4796 0 1 3975
box -3 -3 3 3
use FILL  FILL_1703
timestamp 1677677812
transform 1 0 4784 0 1 3970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_15
timestamp 1677677812
transform 1 0 4819 0 1 3970
box -10 -3 10 3
use M3_M2  M3_M2_1362
timestamp 1677677812
transform 1 0 196 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1383
timestamp 1677677812
transform 1 0 180 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1384
timestamp 1677677812
transform 1 0 212 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1616
timestamp 1677677812
transform 1 0 84 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1412
timestamp 1677677812
transform 1 0 164 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1617
timestamp 1677677812
transform 1 0 180 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1618
timestamp 1677677812
transform 1 0 196 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1709
timestamp 1677677812
transform 1 0 132 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1428
timestamp 1677677812
transform 1 0 148 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1413
timestamp 1677677812
transform 1 0 220 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1710
timestamp 1677677812
transform 1 0 164 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1711
timestamp 1677677812
transform 1 0 172 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1429
timestamp 1677677812
transform 1 0 180 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1712
timestamp 1677677812
transform 1 0 244 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1442
timestamp 1677677812
transform 1 0 132 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1443
timestamp 1677677812
transform 1 0 172 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1619
timestamp 1677677812
transform 1 0 300 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1414
timestamp 1677677812
transform 1 0 308 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1363
timestamp 1677677812
transform 1 0 340 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1620
timestamp 1677677812
transform 1 0 316 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1621
timestamp 1677677812
transform 1 0 332 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1713
timestamp 1677677812
transform 1 0 300 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1714
timestamp 1677677812
transform 1 0 308 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1715
timestamp 1677677812
transform 1 0 324 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1476
timestamp 1677677812
transform 1 0 292 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1364
timestamp 1677677812
transform 1 0 364 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1365
timestamp 1677677812
transform 1 0 444 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1385
timestamp 1677677812
transform 1 0 444 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1622
timestamp 1677677812
transform 1 0 364 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1716
timestamp 1677677812
transform 1 0 412 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1717
timestamp 1677677812
transform 1 0 444 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1718
timestamp 1677677812
transform 1 0 452 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1444
timestamp 1677677812
transform 1 0 412 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1445
timestamp 1677677812
transform 1 0 452 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1386
timestamp 1677677812
transform 1 0 516 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1623
timestamp 1677677812
transform 1 0 492 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1624
timestamp 1677677812
transform 1 0 500 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1625
timestamp 1677677812
transform 1 0 516 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1719
timestamp 1677677812
transform 1 0 492 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1430
timestamp 1677677812
transform 1 0 500 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1720
timestamp 1677677812
transform 1 0 508 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1721
timestamp 1677677812
transform 1 0 524 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1485
timestamp 1677677812
transform 1 0 492 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1477
timestamp 1677677812
transform 1 0 524 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1722
timestamp 1677677812
transform 1 0 556 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1626
timestamp 1677677812
transform 1 0 580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1723
timestamp 1677677812
transform 1 0 572 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1431
timestamp 1677677812
transform 1 0 588 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1724
timestamp 1677677812
transform 1 0 612 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1446
timestamp 1677677812
transform 1 0 620 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1494
timestamp 1677677812
transform 1 0 612 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1627
timestamp 1677677812
transform 1 0 636 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1628
timestamp 1677677812
transform 1 0 644 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1629
timestamp 1677677812
transform 1 0 668 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1630
timestamp 1677677812
transform 1 0 676 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1432
timestamp 1677677812
transform 1 0 636 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1725
timestamp 1677677812
transform 1 0 644 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1726
timestamp 1677677812
transform 1 0 660 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1433
timestamp 1677677812
transform 1 0 668 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1447
timestamp 1677677812
transform 1 0 660 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1478
timestamp 1677677812
transform 1 0 644 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1727
timestamp 1677677812
transform 1 0 684 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1728
timestamp 1677677812
transform 1 0 740 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1448
timestamp 1677677812
transform 1 0 740 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1415
timestamp 1677677812
transform 1 0 812 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1631
timestamp 1677677812
transform 1 0 836 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1729
timestamp 1677677812
transform 1 0 756 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1434
timestamp 1677677812
transform 1 0 764 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1730
timestamp 1677677812
transform 1 0 788 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1449
timestamp 1677677812
transform 1 0 788 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1416
timestamp 1677677812
transform 1 0 852 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1731
timestamp 1677677812
transform 1 0 852 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1732
timestamp 1677677812
transform 1 0 892 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1479
timestamp 1677677812
transform 1 0 892 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1632
timestamp 1677677812
transform 1 0 908 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1450
timestamp 1677677812
transform 1 0 908 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1633
timestamp 1677677812
transform 1 0 924 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1634
timestamp 1677677812
transform 1 0 956 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1733
timestamp 1677677812
transform 1 0 948 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1734
timestamp 1677677812
transform 1 0 964 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1451
timestamp 1677677812
transform 1 0 948 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1366
timestamp 1677677812
transform 1 0 980 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1387
timestamp 1677677812
transform 1 0 996 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1367
timestamp 1677677812
transform 1 0 1012 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1368
timestamp 1677677812
transform 1 0 1028 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1369
timestamp 1677677812
transform 1 0 1044 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1635
timestamp 1677677812
transform 1 0 1012 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1735
timestamp 1677677812
transform 1 0 1036 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1736
timestamp 1677677812
transform 1 0 1092 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1435
timestamp 1677677812
transform 1 0 1108 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1737
timestamp 1677677812
transform 1 0 1132 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1636
timestamp 1677677812
transform 1 0 1220 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1738
timestamp 1677677812
transform 1 0 1196 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1436
timestamp 1677677812
transform 1 0 1220 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1480
timestamp 1677677812
transform 1 0 1156 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1388
timestamp 1677677812
transform 1 0 1236 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1637
timestamp 1677677812
transform 1 0 1236 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1481
timestamp 1677677812
transform 1 0 1236 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1822
timestamp 1677677812
transform 1 0 1252 0 1 3915
box -2 -2 2 2
use M3_M2  M3_M2_1341
timestamp 1677677812
transform 1 0 1268 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1739
timestamp 1677677812
transform 1 0 1300 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1638
timestamp 1677677812
transform 1 0 1324 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1342
timestamp 1677677812
transform 1 0 1348 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1417
timestamp 1677677812
transform 1 0 1388 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1639
timestamp 1677677812
transform 1 0 1412 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1740
timestamp 1677677812
transform 1 0 1332 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1452
timestamp 1677677812
transform 1 0 1324 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1437
timestamp 1677677812
transform 1 0 1372 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1741
timestamp 1677677812
transform 1 0 1388 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1640
timestamp 1677677812
transform 1 0 1428 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1418
timestamp 1677677812
transform 1 0 1444 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1742
timestamp 1677677812
transform 1 0 1460 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1641
timestamp 1677677812
transform 1 0 1548 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1743
timestamp 1677677812
transform 1 0 1588 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1744
timestamp 1677677812
transform 1 0 1628 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1745
timestamp 1677677812
transform 1 0 1636 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1453
timestamp 1677677812
transform 1 0 1636 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1642
timestamp 1677677812
transform 1 0 1652 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1643
timestamp 1677677812
transform 1 0 1676 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1746
timestamp 1677677812
transform 1 0 1668 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1438
timestamp 1677677812
transform 1 0 1676 0 1 3925
box -3 -3 3 3
use M2_M1  M2_M1_1747
timestamp 1677677812
transform 1 0 1700 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1454
timestamp 1677677812
transform 1 0 1700 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1419
timestamp 1677677812
transform 1 0 1716 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1748
timestamp 1677677812
transform 1 0 1716 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1455
timestamp 1677677812
transform 1 0 1732 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1482
timestamp 1677677812
transform 1 0 1788 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1370
timestamp 1677677812
transform 1 0 1804 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1644
timestamp 1677677812
transform 1 0 1812 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1749
timestamp 1677677812
transform 1 0 1804 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1750
timestamp 1677677812
transform 1 0 1820 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1456
timestamp 1677677812
transform 1 0 1820 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1751
timestamp 1677677812
transform 1 0 1852 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1389
timestamp 1677677812
transform 1 0 1900 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1645
timestamp 1677677812
transform 1 0 1900 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1752
timestamp 1677677812
transform 1 0 1892 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1457
timestamp 1677677812
transform 1 0 1884 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1390
timestamp 1677677812
transform 1 0 1916 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1646
timestamp 1677677812
transform 1 0 1924 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1420
timestamp 1677677812
transform 1 0 1932 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1753
timestamp 1677677812
transform 1 0 1916 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1754
timestamp 1677677812
transform 1 0 1932 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1495
timestamp 1677677812
transform 1 0 1916 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1647
timestamp 1677677812
transform 1 0 1948 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1824
timestamp 1677677812
transform 1 0 1948 0 1 3885
box -2 -2 2 2
use M3_M2  M3_M2_1391
timestamp 1677677812
transform 1 0 1972 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1755
timestamp 1677677812
transform 1 0 1996 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1486
timestamp 1677677812
transform 1 0 1996 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1496
timestamp 1677677812
transform 1 0 1988 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1825
timestamp 1677677812
transform 1 0 1996 0 1 3885
box -2 -2 2 2
use M3_M2  M3_M2_1343
timestamp 1677677812
transform 1 0 2020 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1344
timestamp 1677677812
transform 1 0 2044 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1371
timestamp 1677677812
transform 1 0 2036 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1392
timestamp 1677677812
transform 1 0 2028 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1648
timestamp 1677677812
transform 1 0 2028 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1756
timestamp 1677677812
transform 1 0 2020 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1757
timestamp 1677677812
transform 1 0 2036 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1393
timestamp 1677677812
transform 1 0 2060 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1649
timestamp 1677677812
transform 1 0 2060 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1650
timestamp 1677677812
transform 1 0 2092 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1458
timestamp 1677677812
transform 1 0 2092 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1394
timestamp 1677677812
transform 1 0 2116 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1758
timestamp 1677677812
transform 1 0 2108 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1497
timestamp 1677677812
transform 1 0 2108 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1651
timestamp 1677677812
transform 1 0 2116 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1759
timestamp 1677677812
transform 1 0 2124 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1345
timestamp 1677677812
transform 1 0 2148 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1372
timestamp 1677677812
transform 1 0 2164 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1652
timestamp 1677677812
transform 1 0 2148 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1653
timestamp 1677677812
transform 1 0 2164 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1760
timestamp 1677677812
transform 1 0 2156 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1459
timestamp 1677677812
transform 1 0 2156 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1761
timestamp 1677677812
transform 1 0 2180 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1487
timestamp 1677677812
transform 1 0 2180 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1498
timestamp 1677677812
transform 1 0 2188 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1762
timestamp 1677677812
transform 1 0 2212 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1373
timestamp 1677677812
transform 1 0 2236 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1395
timestamp 1677677812
transform 1 0 2228 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1654
timestamp 1677677812
transform 1 0 2228 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1655
timestamp 1677677812
transform 1 0 2236 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1346
timestamp 1677677812
transform 1 0 2252 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1347
timestamp 1677677812
transform 1 0 2276 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1656
timestamp 1677677812
transform 1 0 2276 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1763
timestamp 1677677812
transform 1 0 2268 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1764
timestamp 1677677812
transform 1 0 2292 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1460
timestamp 1677677812
transform 1 0 2276 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1461
timestamp 1677677812
transform 1 0 2292 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1657
timestamp 1677677812
transform 1 0 2308 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1374
timestamp 1677677812
transform 1 0 2324 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1658
timestamp 1677677812
transform 1 0 2324 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1659
timestamp 1677677812
transform 1 0 2340 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1660
timestamp 1677677812
transform 1 0 2348 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1765
timestamp 1677677812
transform 1 0 2316 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1766
timestamp 1677677812
transform 1 0 2332 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1462
timestamp 1677677812
transform 1 0 2308 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1463
timestamp 1677677812
transform 1 0 2340 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1767
timestamp 1677677812
transform 1 0 2356 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1375
timestamp 1677677812
transform 1 0 2380 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1464
timestamp 1677677812
transform 1 0 2380 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1661
timestamp 1677677812
transform 1 0 2412 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1768
timestamp 1677677812
transform 1 0 2428 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1769
timestamp 1677677812
transform 1 0 2484 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1662
timestamp 1677677812
transform 1 0 2500 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1465
timestamp 1677677812
transform 1 0 2500 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1663
timestamp 1677677812
transform 1 0 2532 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1664
timestamp 1677677812
transform 1 0 2556 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1770
timestamp 1677677812
transform 1 0 2540 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1771
timestamp 1677677812
transform 1 0 2548 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1772
timestamp 1677677812
transform 1 0 2564 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1773
timestamp 1677677812
transform 1 0 2580 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1488
timestamp 1677677812
transform 1 0 2540 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1466
timestamp 1677677812
transform 1 0 2564 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1665
timestamp 1677677812
transform 1 0 2596 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1467
timestamp 1677677812
transform 1 0 2596 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1376
timestamp 1677677812
transform 1 0 2612 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1666
timestamp 1677677812
transform 1 0 2612 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1774
timestamp 1677677812
transform 1 0 2636 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1775
timestamp 1677677812
transform 1 0 2692 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1468
timestamp 1677677812
transform 1 0 2692 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1489
timestamp 1677677812
transform 1 0 2636 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1469
timestamp 1677677812
transform 1 0 2716 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1348
timestamp 1677677812
transform 1 0 2780 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1667
timestamp 1677677812
transform 1 0 2732 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1776
timestamp 1677677812
transform 1 0 2764 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1777
timestamp 1677677812
transform 1 0 2812 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1490
timestamp 1677677812
transform 1 0 2796 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1778
timestamp 1677677812
transform 1 0 2852 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1615
timestamp 1677677812
transform 1 0 2884 0 1 3945
box -2 -2 2 2
use M2_M1  M2_M1_1668
timestamp 1677677812
transform 1 0 2876 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1421
timestamp 1677677812
transform 1 0 2884 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1823
timestamp 1677677812
transform 1 0 2900 0 1 3915
box -2 -2 2 2
use M2_M1  M2_M1_1779
timestamp 1677677812
transform 1 0 2924 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1483
timestamp 1677677812
transform 1 0 2932 0 1 3905
box -3 -3 3 3
use M3_M2  M3_M2_1491
timestamp 1677677812
transform 1 0 2924 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1669
timestamp 1677677812
transform 1 0 2948 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1349
timestamp 1677677812
transform 1 0 2964 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1350
timestamp 1677677812
transform 1 0 3044 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1396
timestamp 1677677812
transform 1 0 2964 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1397
timestamp 1677677812
transform 1 0 3012 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1670
timestamp 1677677812
transform 1 0 2964 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1780
timestamp 1677677812
transform 1 0 3012 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1484
timestamp 1677677812
transform 1 0 2996 0 1 3905
box -3 -3 3 3
use M2_M1  M2_M1_1781
timestamp 1677677812
transform 1 0 3068 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1470
timestamp 1677677812
transform 1 0 3068 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1671
timestamp 1677677812
transform 1 0 3108 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1398
timestamp 1677677812
transform 1 0 3140 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1672
timestamp 1677677812
transform 1 0 3140 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1782
timestamp 1677677812
transform 1 0 3132 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1471
timestamp 1677677812
transform 1 0 3132 0 1 3915
box -3 -3 3 3
use M2_M1  M2_M1_1783
timestamp 1677677812
transform 1 0 3172 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1399
timestamp 1677677812
transform 1 0 3188 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1673
timestamp 1677677812
transform 1 0 3188 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1674
timestamp 1677677812
transform 1 0 3220 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1784
timestamp 1677677812
transform 1 0 3244 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1785
timestamp 1677677812
transform 1 0 3300 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1351
timestamp 1677677812
transform 1 0 3380 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1352
timestamp 1677677812
transform 1 0 3412 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1400
timestamp 1677677812
transform 1 0 3388 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1675
timestamp 1677677812
transform 1 0 3420 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1786
timestamp 1677677812
transform 1 0 3340 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1787
timestamp 1677677812
transform 1 0 3388 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1353
timestamp 1677677812
transform 1 0 3452 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1354
timestamp 1677677812
transform 1 0 3492 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1401
timestamp 1677677812
transform 1 0 3492 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1676
timestamp 1677677812
transform 1 0 3476 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1677
timestamp 1677677812
transform 1 0 3492 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1422
timestamp 1677677812
transform 1 0 3500 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1678
timestamp 1677677812
transform 1 0 3508 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1788
timestamp 1677677812
transform 1 0 3484 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1789
timestamp 1677677812
transform 1 0 3500 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1790
timestamp 1677677812
transform 1 0 3540 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1355
timestamp 1677677812
transform 1 0 3580 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1356
timestamp 1677677812
transform 1 0 3604 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1357
timestamp 1677677812
transform 1 0 3620 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1402
timestamp 1677677812
transform 1 0 3596 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1679
timestamp 1677677812
transform 1 0 3580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1680
timestamp 1677677812
transform 1 0 3596 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1423
timestamp 1677677812
transform 1 0 3604 0 1 3935
box -3 -3 3 3
use M3_M2  M3_M2_1377
timestamp 1677677812
transform 1 0 3716 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1403
timestamp 1677677812
transform 1 0 3652 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1681
timestamp 1677677812
transform 1 0 3612 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1682
timestamp 1677677812
transform 1 0 3700 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1683
timestamp 1677677812
transform 1 0 3716 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1791
timestamp 1677677812
transform 1 0 3588 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1792
timestamp 1677677812
transform 1 0 3604 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1793
timestamp 1677677812
transform 1 0 3612 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1794
timestamp 1677677812
transform 1 0 3652 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1499
timestamp 1677677812
transform 1 0 3604 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1439
timestamp 1677677812
transform 1 0 3700 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1500
timestamp 1677677812
transform 1 0 3644 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1501
timestamp 1677677812
transform 1 0 3660 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1404
timestamp 1677677812
transform 1 0 3748 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1684
timestamp 1677677812
transform 1 0 3748 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1795
timestamp 1677677812
transform 1 0 3740 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1358
timestamp 1677677812
transform 1 0 3788 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1796
timestamp 1677677812
transform 1 0 3828 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1359
timestamp 1677677812
transform 1 0 3860 0 1 3965
box -3 -3 3 3
use M2_M1  M2_M1_1685
timestamp 1677677812
transform 1 0 3844 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1686
timestamp 1677677812
transform 1 0 3860 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1797
timestamp 1677677812
transform 1 0 3852 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1798
timestamp 1677677812
transform 1 0 3868 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1502
timestamp 1677677812
transform 1 0 3844 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1687
timestamp 1677677812
transform 1 0 3884 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1688
timestamp 1677677812
transform 1 0 3892 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1689
timestamp 1677677812
transform 1 0 3916 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1799
timestamp 1677677812
transform 1 0 3956 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1800
timestamp 1677677812
transform 1 0 3996 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1503
timestamp 1677677812
transform 1 0 3924 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1378
timestamp 1677677812
transform 1 0 4052 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1405
timestamp 1677677812
transform 1 0 4020 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1690
timestamp 1677677812
transform 1 0 4020 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1801
timestamp 1677677812
transform 1 0 4060 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1802
timestamp 1677677812
transform 1 0 4100 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1691
timestamp 1677677812
transform 1 0 4132 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1803
timestamp 1677677812
transform 1 0 4180 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1472
timestamp 1677677812
transform 1 0 4180 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1504
timestamp 1677677812
transform 1 0 4180 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1379
timestamp 1677677812
transform 1 0 4236 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1406
timestamp 1677677812
transform 1 0 4228 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1407
timestamp 1677677812
transform 1 0 4276 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1692
timestamp 1677677812
transform 1 0 4236 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1693
timestamp 1677677812
transform 1 0 4252 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1694
timestamp 1677677812
transform 1 0 4268 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1695
timestamp 1677677812
transform 1 0 4276 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1804
timestamp 1677677812
transform 1 0 4228 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1805
timestamp 1677677812
transform 1 0 4236 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1806
timestamp 1677677812
transform 1 0 4244 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1807
timestamp 1677677812
transform 1 0 4260 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1505
timestamp 1677677812
transform 1 0 4220 0 1 3885
box -3 -3 3 3
use M3_M2  M3_M2_1473
timestamp 1677677812
transform 1 0 4252 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1492
timestamp 1677677812
transform 1 0 4260 0 1 3895
box -3 -3 3 3
use M2_M1  M2_M1_1808
timestamp 1677677812
transform 1 0 4276 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1493
timestamp 1677677812
transform 1 0 4276 0 1 3895
box -3 -3 3 3
use M3_M2  M3_M2_1506
timestamp 1677677812
transform 1 0 4268 0 1 3885
box -3 -3 3 3
use M2_M1  M2_M1_1696
timestamp 1677677812
transform 1 0 4316 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1697
timestamp 1677677812
transform 1 0 4356 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1424
timestamp 1677677812
transform 1 0 4364 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1698
timestamp 1677677812
transform 1 0 4372 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1809
timestamp 1677677812
transform 1 0 4348 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1810
timestamp 1677677812
transform 1 0 4364 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1474
timestamp 1677677812
transform 1 0 4356 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1360
timestamp 1677677812
transform 1 0 4396 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1361
timestamp 1677677812
transform 1 0 4436 0 1 3965
box -3 -3 3 3
use M3_M2  M3_M2_1380
timestamp 1677677812
transform 1 0 4476 0 1 3955
box -3 -3 3 3
use M2_M1  M2_M1_1699
timestamp 1677677812
transform 1 0 4396 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1811
timestamp 1677677812
transform 1 0 4420 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1440
timestamp 1677677812
transform 1 0 4468 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1475
timestamp 1677677812
transform 1 0 4420 0 1 3915
box -3 -3 3 3
use M3_M2  M3_M2_1425
timestamp 1677677812
transform 1 0 4492 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1700
timestamp 1677677812
transform 1 0 4500 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1812
timestamp 1677677812
transform 1 0 4492 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1813
timestamp 1677677812
transform 1 0 4500 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1441
timestamp 1677677812
transform 1 0 4516 0 1 3925
box -3 -3 3 3
use M3_M2  M3_M2_1381
timestamp 1677677812
transform 1 0 4556 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1408
timestamp 1677677812
transform 1 0 4540 0 1 3945
box -3 -3 3 3
use M3_M2  M3_M2_1409
timestamp 1677677812
transform 1 0 4564 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1701
timestamp 1677677812
transform 1 0 4548 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1814
timestamp 1677677812
transform 1 0 4540 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1815
timestamp 1677677812
transform 1 0 4556 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1816
timestamp 1677677812
transform 1 0 4572 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1702
timestamp 1677677812
transform 1 0 4580 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1703
timestamp 1677677812
transform 1 0 4604 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1426
timestamp 1677677812
transform 1 0 4620 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1817
timestamp 1677677812
transform 1 0 4612 0 1 3925
box -2 -2 2 2
use M3_M2  M3_M2_1410
timestamp 1677677812
transform 1 0 4652 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1704
timestamp 1677677812
transform 1 0 4636 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1427
timestamp 1677677812
transform 1 0 4644 0 1 3935
box -3 -3 3 3
use M2_M1  M2_M1_1705
timestamp 1677677812
transform 1 0 4652 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1706
timestamp 1677677812
transform 1 0 4668 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1818
timestamp 1677677812
transform 1 0 4636 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1819
timestamp 1677677812
transform 1 0 4660 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1707
timestamp 1677677812
transform 1 0 4684 0 1 3935
box -2 -2 2 2
use M3_M2  M3_M2_1382
timestamp 1677677812
transform 1 0 4764 0 1 3955
box -3 -3 3 3
use M3_M2  M3_M2_1411
timestamp 1677677812
transform 1 0 4724 0 1 3945
box -3 -3 3 3
use M2_M1  M2_M1_1708
timestamp 1677677812
transform 1 0 4700 0 1 3935
box -2 -2 2 2
use M2_M1  M2_M1_1820
timestamp 1677677812
transform 1 0 4724 0 1 3925
box -2 -2 2 2
use M2_M1  M2_M1_1821
timestamp 1677677812
transform 1 0 4780 0 1 3925
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_16
timestamp 1677677812
transform 1 0 24 0 1 3870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_100
timestamp 1677677812
transform 1 0 72 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_120
timestamp 1677677812
transform -1 0 184 0 -1 3970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_101
timestamp 1677677812
transform 1 0 184 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1279
timestamp 1677677812
transform 1 0 280 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1280
timestamp 1677677812
transform 1 0 288 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_65
timestamp 1677677812
transform 1 0 296 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1281
timestamp 1677677812
transform 1 0 336 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1282
timestamp 1677677812
transform 1 0 344 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_102
timestamp 1677677812
transform 1 0 352 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1283
timestamp 1677677812
transform 1 0 448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1284
timestamp 1677677812
transform 1 0 456 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_121
timestamp 1677677812
transform -1 0 480 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1285
timestamp 1677677812
transform 1 0 480 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_66
timestamp 1677677812
transform 1 0 488 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1286
timestamp 1677677812
transform 1 0 528 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1288
timestamp 1677677812
transform 1 0 536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1292
timestamp 1677677812
transform 1 0 544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1293
timestamp 1677677812
transform 1 0 552 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_66
timestamp 1677677812
transform -1 0 600 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1294
timestamp 1677677812
transform 1 0 600 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1296
timestamp 1677677812
transform 1 0 608 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1301
timestamp 1677677812
transform 1 0 616 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1302
timestamp 1677677812
transform 1 0 624 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1303
timestamp 1677677812
transform 1 0 632 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_69
timestamp 1677677812
transform 1 0 640 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1304
timestamp 1677677812
transform 1 0 680 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1307
timestamp 1677677812
transform 1 0 688 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1308
timestamp 1677677812
transform 1 0 696 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_122
timestamp 1677677812
transform 1 0 704 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1309
timestamp 1677677812
transform 1 0 720 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1310
timestamp 1677677812
transform 1 0 728 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1311
timestamp 1677677812
transform 1 0 736 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1315
timestamp 1677677812
transform 1 0 744 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_104
timestamp 1677677812
transform -1 0 848 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1316
timestamp 1677677812
transform 1 0 848 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1317
timestamp 1677677812
transform 1 0 856 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1318
timestamp 1677677812
transform 1 0 864 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_124
timestamp 1677677812
transform -1 0 888 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1319
timestamp 1677677812
transform 1 0 888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1320
timestamp 1677677812
transform 1 0 896 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1322
timestamp 1677677812
transform 1 0 904 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1324
timestamp 1677677812
transform 1 0 912 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1326
timestamp 1677677812
transform 1 0 920 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_70
timestamp 1677677812
transform 1 0 928 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1333
timestamp 1677677812
transform 1 0 968 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1335
timestamp 1677677812
transform 1 0 976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1336
timestamp 1677677812
transform 1 0 984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1337
timestamp 1677677812
transform 1 0 992 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_105
timestamp 1677677812
transform 1 0 1000 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1346
timestamp 1677677812
transform 1 0 1096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1348
timestamp 1677677812
transform 1 0 1104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1350
timestamp 1677677812
transform 1 0 1112 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1352
timestamp 1677677812
transform 1 0 1120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1359
timestamp 1677677812
transform 1 0 1128 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_106
timestamp 1677677812
transform -1 0 1232 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1360
timestamp 1677677812
transform 1 0 1232 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1361
timestamp 1677677812
transform 1 0 1240 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1363
timestamp 1677677812
transform 1 0 1248 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_37
timestamp 1677677812
transform -1 0 1288 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1376
timestamp 1677677812
transform 1 0 1288 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1377
timestamp 1677677812
transform 1 0 1296 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1378
timestamp 1677677812
transform 1 0 1304 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1379
timestamp 1677677812
transform 1 0 1312 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1380
timestamp 1677677812
transform 1 0 1320 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_107
timestamp 1677677812
transform -1 0 1424 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1381
timestamp 1677677812
transform 1 0 1424 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1382
timestamp 1677677812
transform 1 0 1432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1383
timestamp 1677677812
transform 1 0 1440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1384
timestamp 1677677812
transform 1 0 1448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1385
timestamp 1677677812
transform 1 0 1456 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1386
timestamp 1677677812
transform 1 0 1464 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_127
timestamp 1677677812
transform 1 0 1472 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1390
timestamp 1677677812
transform 1 0 1488 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1392
timestamp 1677677812
transform 1 0 1496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1394
timestamp 1677677812
transform 1 0 1504 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1396
timestamp 1677677812
transform 1 0 1512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1398
timestamp 1677677812
transform 1 0 1520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1400
timestamp 1677677812
transform 1 0 1528 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_109
timestamp 1677677812
transform 1 0 1536 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1402
timestamp 1677677812
transform 1 0 1632 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1404
timestamp 1677677812
transform 1 0 1640 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_129
timestamp 1677677812
transform 1 0 1648 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1407
timestamp 1677677812
transform 1 0 1664 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1408
timestamp 1677677812
transform 1 0 1672 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1409
timestamp 1677677812
transform 1 0 1680 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_130
timestamp 1677677812
transform 1 0 1688 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1410
timestamp 1677677812
transform 1 0 1704 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1411
timestamp 1677677812
transform 1 0 1712 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1413
timestamp 1677677812
transform 1 0 1720 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1415
timestamp 1677677812
transform 1 0 1728 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1417
timestamp 1677677812
transform 1 0 1736 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1419
timestamp 1677677812
transform 1 0 1744 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1421
timestamp 1677677812
transform 1 0 1752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1423
timestamp 1677677812
transform 1 0 1760 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1425
timestamp 1677677812
transform 1 0 1768 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1427
timestamp 1677677812
transform 1 0 1776 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1429
timestamp 1677677812
transform 1 0 1784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1436
timestamp 1677677812
transform 1 0 1792 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_73
timestamp 1677677812
transform 1 0 1800 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1437
timestamp 1677677812
transform 1 0 1840 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1438
timestamp 1677677812
transform 1 0 1848 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1439
timestamp 1677677812
transform 1 0 1856 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1440
timestamp 1677677812
transform 1 0 1864 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1441
timestamp 1677677812
transform 1 0 1872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1442
timestamp 1677677812
transform 1 0 1880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1443
timestamp 1677677812
transform 1 0 1888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1444
timestamp 1677677812
transform 1 0 1896 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_70
timestamp 1677677812
transform 1 0 1904 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1445
timestamp 1677677812
transform 1 0 1944 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1446
timestamp 1677677812
transform 1 0 1952 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1447
timestamp 1677677812
transform 1 0 1960 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1448
timestamp 1677677812
transform 1 0 1968 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1449
timestamp 1677677812
transform 1 0 1976 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1450
timestamp 1677677812
transform 1 0 1984 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1451
timestamp 1677677812
transform 1 0 1992 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_74
timestamp 1677677812
transform -1 0 2040 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1452
timestamp 1677677812
transform 1 0 2040 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1454
timestamp 1677677812
transform 1 0 2048 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1455
timestamp 1677677812
transform 1 0 2056 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1456
timestamp 1677677812
transform 1 0 2064 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1459
timestamp 1677677812
transform 1 0 2072 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1460
timestamp 1677677812
transform 1 0 2080 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_133
timestamp 1677677812
transform 1 0 2088 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1461
timestamp 1677677812
transform 1 0 2104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1462
timestamp 1677677812
transform 1 0 2112 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1463
timestamp 1677677812
transform 1 0 2120 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1464
timestamp 1677677812
transform 1 0 2128 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_75
timestamp 1677677812
transform 1 0 2136 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1465
timestamp 1677677812
transform 1 0 2176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1468
timestamp 1677677812
transform 1 0 2184 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1507
timestamp 1677677812
transform 1 0 2204 0 1 3875
box -3 -3 3 3
use FILL  FILL_1469
timestamp 1677677812
transform 1 0 2192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1470
timestamp 1677677812
transform 1 0 2200 0 -1 3970
box -8 -3 16 105
use BUFX2  BUFX2_5
timestamp 1677677812
transform 1 0 2208 0 -1 3970
box -5 -3 28 105
use FILL  FILL_1471
timestamp 1677677812
transform 1 0 2232 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1472
timestamp 1677677812
transform 1 0 2240 0 -1 3970
box -8 -3 16 105
use M3_M2  M3_M2_1508
timestamp 1677677812
transform 1 0 2260 0 1 3875
box -3 -3 3 3
use FILL  FILL_1475
timestamp 1677677812
transform 1 0 2248 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_71
timestamp 1677677812
transform -1 0 2296 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1476
timestamp 1677677812
transform 1 0 2296 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1478
timestamp 1677677812
transform 1 0 2304 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_77
timestamp 1677677812
transform 1 0 2312 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1482
timestamp 1677677812
transform 1 0 2352 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1484
timestamp 1677677812
transform 1 0 2360 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1486
timestamp 1677677812
transform 1 0 2368 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1488
timestamp 1677677812
transform 1 0 2376 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1489
timestamp 1677677812
transform 1 0 2384 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_134
timestamp 1677677812
transform 1 0 2392 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1490
timestamp 1677677812
transform 1 0 2408 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1491
timestamp 1677677812
transform 1 0 2416 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1493
timestamp 1677677812
transform 1 0 2424 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1495
timestamp 1677677812
transform 1 0 2432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1509
timestamp 1677677812
transform 1 0 2440 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_135
timestamp 1677677812
transform 1 0 2448 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1510
timestamp 1677677812
transform 1 0 2464 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1511
timestamp 1677677812
transform 1 0 2472 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1512
timestamp 1677677812
transform 1 0 2480 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1513
timestamp 1677677812
transform 1 0 2488 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_136
timestamp 1677677812
transform 1 0 2496 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1514
timestamp 1677677812
transform 1 0 2512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1515
timestamp 1677677812
transform 1 0 2520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1516
timestamp 1677677812
transform 1 0 2528 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1517
timestamp 1677677812
transform 1 0 2536 0 -1 3970
box -8 -3 16 105
use AOI22X1  AOI22X1_81
timestamp 1677677812
transform 1 0 2544 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1518
timestamp 1677677812
transform 1 0 2584 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1519
timestamp 1677677812
transform 1 0 2592 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_114
timestamp 1677677812
transform 1 0 2600 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1520
timestamp 1677677812
transform 1 0 2696 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1521
timestamp 1677677812
transform 1 0 2704 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1522
timestamp 1677677812
transform 1 0 2712 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_115
timestamp 1677677812
transform 1 0 2720 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1534
timestamp 1677677812
transform 1 0 2816 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1536
timestamp 1677677812
transform 1 0 2824 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1538
timestamp 1677677812
transform 1 0 2832 0 -1 3970
box -8 -3 16 105
use OAI21X1  OAI21X1_39
timestamp 1677677812
transform 1 0 2840 0 -1 3970
box -8 -3 34 105
use FILL  FILL_1542
timestamp 1677677812
transform 1 0 2872 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1543
timestamp 1677677812
transform 1 0 2880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1544
timestamp 1677677812
transform 1 0 2888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1546
timestamp 1677677812
transform 1 0 2896 0 -1 3970
box -8 -3 16 105
use NOR2X1  NOR2X1_18
timestamp 1677677812
transform 1 0 2904 0 -1 3970
box -8 -3 32 105
use FILL  FILL_1551
timestamp 1677677812
transform 1 0 2928 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1553
timestamp 1677677812
transform 1 0 2936 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1555
timestamp 1677677812
transform 1 0 2944 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_117
timestamp 1677677812
transform 1 0 2952 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1567
timestamp 1677677812
transform 1 0 3048 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_138
timestamp 1677677812
transform 1 0 3056 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1568
timestamp 1677677812
transform 1 0 3072 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1569
timestamp 1677677812
transform 1 0 3080 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1570
timestamp 1677677812
transform 1 0 3088 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1571
timestamp 1677677812
transform 1 0 3096 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1572
timestamp 1677677812
transform 1 0 3104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1573
timestamp 1677677812
transform 1 0 3112 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_73
timestamp 1677677812
transform -1 0 3160 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1574
timestamp 1677677812
transform 1 0 3160 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1575
timestamp 1677677812
transform 1 0 3168 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1576
timestamp 1677677812
transform 1 0 3176 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1577
timestamp 1677677812
transform 1 0 3184 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1578
timestamp 1677677812
transform 1 0 3192 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1579
timestamp 1677677812
transform 1 0 3200 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_119
timestamp 1677677812
transform 1 0 3208 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1589
timestamp 1677677812
transform 1 0 3304 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1590
timestamp 1677677812
transform 1 0 3312 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1591
timestamp 1677677812
transform 1 0 3320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1592
timestamp 1677677812
transform 1 0 3328 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_120
timestamp 1677677812
transform -1 0 3432 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1593
timestamp 1677677812
transform 1 0 3432 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1594
timestamp 1677677812
transform 1 0 3440 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1610
timestamp 1677677812
transform 1 0 3448 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1611
timestamp 1677677812
transform 1 0 3456 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1612
timestamp 1677677812
transform 1 0 3464 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_75
timestamp 1677677812
transform -1 0 3512 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1613
timestamp 1677677812
transform 1 0 3512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1614
timestamp 1677677812
transform 1 0 3520 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1615
timestamp 1677677812
transform 1 0 3528 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1616
timestamp 1677677812
transform 1 0 3536 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1617
timestamp 1677677812
transform 1 0 3544 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1618
timestamp 1677677812
transform 1 0 3552 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1619
timestamp 1677677812
transform 1 0 3560 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1620
timestamp 1677677812
transform 1 0 3568 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_76
timestamp 1677677812
transform -1 0 3616 0 -1 3970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_122
timestamp 1677677812
transform -1 0 3712 0 -1 3970
box -8 -3 104 105
use BUFX2  BUFX2_9
timestamp 1677677812
transform -1 0 3736 0 -1 3970
box -5 -3 28 105
use FILL  FILL_1621
timestamp 1677677812
transform 1 0 3736 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1623
timestamp 1677677812
transform 1 0 3744 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1627
timestamp 1677677812
transform 1 0 3752 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1628
timestamp 1677677812
transform 1 0 3760 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1629
timestamp 1677677812
transform 1 0 3768 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1630
timestamp 1677677812
transform 1 0 3776 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1631
timestamp 1677677812
transform 1 0 3784 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1632
timestamp 1677677812
transform 1 0 3792 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1633
timestamp 1677677812
transform 1 0 3800 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1634
timestamp 1677677812
transform 1 0 3808 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1635
timestamp 1677677812
transform 1 0 3816 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1636
timestamp 1677677812
transform 1 0 3824 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1637
timestamp 1677677812
transform 1 0 3832 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_77
timestamp 1677677812
transform 1 0 3840 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1638
timestamp 1677677812
transform 1 0 3880 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1640
timestamp 1677677812
transform 1 0 3888 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1650
timestamp 1677677812
transform 1 0 3896 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_126
timestamp 1677677812
transform 1 0 3904 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1651
timestamp 1677677812
transform 1 0 4000 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_127
timestamp 1677677812
transform 1 0 4008 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1652
timestamp 1677677812
transform 1 0 4104 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1653
timestamp 1677677812
transform 1 0 4112 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_128
timestamp 1677677812
transform 1 0 4120 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1654
timestamp 1677677812
transform 1 0 4216 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1656
timestamp 1677677812
transform 1 0 4224 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_79
timestamp 1677677812
transform 1 0 4232 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1658
timestamp 1677677812
transform 1 0 4272 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_144
timestamp 1677677812
transform 1 0 4280 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1671
timestamp 1677677812
transform 1 0 4296 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1672
timestamp 1677677812
transform 1 0 4304 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1673
timestamp 1677677812
transform 1 0 4312 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1674
timestamp 1677677812
transform 1 0 4320 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1675
timestamp 1677677812
transform 1 0 4328 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_81
timestamp 1677677812
transform 1 0 4336 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1676
timestamp 1677677812
transform 1 0 4376 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_130
timestamp 1677677812
transform 1 0 4384 0 -1 3970
box -8 -3 104 105
use INVX2  INVX2_145
timestamp 1677677812
transform 1 0 4480 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1677
timestamp 1677677812
transform 1 0 4496 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1678
timestamp 1677677812
transform 1 0 4504 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1679
timestamp 1677677812
transform 1 0 4512 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1680
timestamp 1677677812
transform 1 0 4520 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_82
timestamp 1677677812
transform 1 0 4528 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1681
timestamp 1677677812
transform 1 0 4568 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1682
timestamp 1677677812
transform 1 0 4576 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1683
timestamp 1677677812
transform 1 0 4584 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1684
timestamp 1677677812
transform 1 0 4592 0 -1 3970
box -8 -3 16 105
use INVX2  INVX2_147
timestamp 1677677812
transform 1 0 4600 0 -1 3970
box -9 -3 26 105
use FILL  FILL_1688
timestamp 1677677812
transform 1 0 4616 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1689
timestamp 1677677812
transform 1 0 4624 0 -1 3970
box -8 -3 16 105
use OAI22X1  OAI22X1_83
timestamp 1677677812
transform 1 0 4632 0 -1 3970
box -8 -3 46 105
use FILL  FILL_1690
timestamp 1677677812
transform 1 0 4672 0 -1 3970
box -8 -3 16 105
use FILL  FILL_1692
timestamp 1677677812
transform 1 0 4680 0 -1 3970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_131
timestamp 1677677812
transform 1 0 4688 0 -1 3970
box -8 -3 104 105
use FILL  FILL_1704
timestamp 1677677812
transform 1 0 4784 0 -1 3970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_17
timestamp 1677677812
transform 1 0 4843 0 1 3870
box -10 -3 10 3
use M2_M1  M2_M1_1835
timestamp 1677677812
transform 1 0 124 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1938
timestamp 1677677812
transform 1 0 92 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1836
timestamp 1677677812
transform 1 0 188 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1837
timestamp 1677677812
transform 1 0 196 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1939
timestamp 1677677812
transform 1 0 180 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1588
timestamp 1677677812
transform 1 0 204 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1838
timestamp 1677677812
transform 1 0 212 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1940
timestamp 1677677812
transform 1 0 196 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1941
timestamp 1677677812
transform 1 0 220 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1942
timestamp 1677677812
transform 1 0 228 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1627
timestamp 1677677812
transform 1 0 188 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1628
timestamp 1677677812
transform 1 0 220 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1559
timestamp 1677677812
transform 1 0 252 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1839
timestamp 1677677812
transform 1 0 244 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1546
timestamp 1677677812
transform 1 0 268 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1589
timestamp 1677677812
transform 1 0 276 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1547
timestamp 1677677812
transform 1 0 324 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1560
timestamp 1677677812
transform 1 0 308 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1840
timestamp 1677677812
transform 1 0 292 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1590
timestamp 1677677812
transform 1 0 300 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1841
timestamp 1677677812
transform 1 0 308 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1591
timestamp 1677677812
transform 1 0 316 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1561
timestamp 1677677812
transform 1 0 388 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1562
timestamp 1677677812
transform 1 0 428 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1842
timestamp 1677677812
transform 1 0 388 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1843
timestamp 1677677812
transform 1 0 420 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1844
timestamp 1677677812
transform 1 0 428 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1943
timestamp 1677677812
transform 1 0 292 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1944
timestamp 1677677812
transform 1 0 300 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1945
timestamp 1677677812
transform 1 0 316 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1946
timestamp 1677677812
transform 1 0 324 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1947
timestamp 1677677812
transform 1 0 340 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1629
timestamp 1677677812
transform 1 0 324 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1630
timestamp 1677677812
transform 1 0 420 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1563
timestamp 1677677812
transform 1 0 444 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1548
timestamp 1677677812
transform 1 0 484 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1564
timestamp 1677677812
transform 1 0 492 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1845
timestamp 1677677812
transform 1 0 484 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1846
timestamp 1677677812
transform 1 0 500 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1847
timestamp 1677677812
transform 1 0 516 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1948
timestamp 1677677812
transform 1 0 484 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1949
timestamp 1677677812
transform 1 0 492 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1950
timestamp 1677677812
transform 1 0 508 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1631
timestamp 1677677812
transform 1 0 508 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1519
timestamp 1677677812
transform 1 0 572 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1565
timestamp 1677677812
transform 1 0 580 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1848
timestamp 1677677812
transform 1 0 580 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1951
timestamp 1677677812
transform 1 0 588 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1849
timestamp 1677677812
transform 1 0 612 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1549
timestamp 1677677812
transform 1 0 636 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1850
timestamp 1677677812
transform 1 0 636 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1613
timestamp 1677677812
transform 1 0 636 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1952
timestamp 1677677812
transform 1 0 644 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1632
timestamp 1677677812
transform 1 0 644 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1851
timestamp 1677677812
transform 1 0 668 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1953
timestamp 1677677812
transform 1 0 660 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1954
timestamp 1677677812
transform 1 0 676 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1633
timestamp 1677677812
transform 1 0 676 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1852
timestamp 1677677812
transform 1 0 692 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1550
timestamp 1677677812
transform 1 0 812 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1853
timestamp 1677677812
transform 1 0 772 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1955
timestamp 1677677812
transform 1 0 812 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1668
timestamp 1677677812
transform 1 0 812 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1551
timestamp 1677677812
transform 1 0 836 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1854
timestamp 1677677812
transform 1 0 828 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1634
timestamp 1677677812
transform 1 0 828 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1635
timestamp 1677677812
transform 1 0 844 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1532
timestamp 1677677812
transform 1 0 884 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1552
timestamp 1677677812
transform 1 0 884 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1855
timestamp 1677677812
transform 1 0 892 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1956
timestamp 1677677812
transform 1 0 884 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1957
timestamp 1677677812
transform 1 0 908 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1553
timestamp 1677677812
transform 1 0 924 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1592
timestamp 1677677812
transform 1 0 924 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2035
timestamp 1677677812
transform 1 0 924 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1533
timestamp 1677677812
transform 1 0 940 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1554
timestamp 1677677812
transform 1 0 948 0 1 3835
box -3 -3 3 3
use M3_M2  M3_M2_1555
timestamp 1677677812
transform 1 0 964 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1856
timestamp 1677677812
transform 1 0 948 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1593
timestamp 1677677812
transform 1 0 956 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1566
timestamp 1677677812
transform 1 0 972 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_2036
timestamp 1677677812
transform 1 0 972 0 1 3795
box -2 -2 2 2
use M2_M1  M2_M1_1857
timestamp 1677677812
transform 1 0 996 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1958
timestamp 1677677812
transform 1 0 996 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1509
timestamp 1677677812
transform 1 0 1012 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1594
timestamp 1677677812
transform 1 0 1036 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1959
timestamp 1677677812
transform 1 0 1028 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1960
timestamp 1677677812
transform 1 0 1036 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1567
timestamp 1677677812
transform 1 0 1084 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1858
timestamp 1677677812
transform 1 0 1084 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1859
timestamp 1677677812
transform 1 0 1092 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1614
timestamp 1677677812
transform 1 0 1092 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1568
timestamp 1677677812
transform 1 0 1116 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1961
timestamp 1677677812
transform 1 0 1116 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1827
timestamp 1677677812
transform 1 0 1156 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1615
timestamp 1677677812
transform 1 0 1148 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1556
timestamp 1677677812
transform 1 0 1172 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1962
timestamp 1677677812
transform 1 0 1172 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1636
timestamp 1677677812
transform 1 0 1172 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1860
timestamp 1677677812
transform 1 0 1196 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1637
timestamp 1677677812
transform 1 0 1196 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1669
timestamp 1677677812
transform 1 0 1212 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1963
timestamp 1677677812
transform 1 0 1236 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1828
timestamp 1677677812
transform 1 0 1252 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1861
timestamp 1677677812
transform 1 0 1268 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1510
timestamp 1677677812
transform 1 0 1292 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1595
timestamp 1677677812
transform 1 0 1308 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1964
timestamp 1677677812
transform 1 0 1308 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1511
timestamp 1677677812
transform 1 0 1380 0 1 3865
box -3 -3 3 3
use M2_M1  M2_M1_1862
timestamp 1677677812
transform 1 0 1364 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1965
timestamp 1677677812
transform 1 0 1324 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1638
timestamp 1677677812
transform 1 0 1364 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1512
timestamp 1677677812
transform 1 0 1420 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1596
timestamp 1677677812
transform 1 0 1436 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1863
timestamp 1677677812
transform 1 0 1444 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1616
timestamp 1677677812
transform 1 0 1444 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1966
timestamp 1677677812
transform 1 0 1484 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1597
timestamp 1677677812
transform 1 0 1500 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1864
timestamp 1677677812
transform 1 0 1508 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1865
timestamp 1677677812
transform 1 0 1524 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1967
timestamp 1677677812
transform 1 0 1516 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1639
timestamp 1677677812
transform 1 0 1516 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1866
timestamp 1677677812
transform 1 0 1540 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1617
timestamp 1677677812
transform 1 0 1548 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1968
timestamp 1677677812
transform 1 0 1580 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1640
timestamp 1677677812
transform 1 0 1588 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1867
timestamp 1677677812
transform 1 0 1620 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1969
timestamp 1677677812
transform 1 0 1628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1970
timestamp 1677677812
transform 1 0 1636 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1641
timestamp 1677677812
transform 1 0 1628 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1618
timestamp 1677677812
transform 1 0 1700 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1971
timestamp 1677677812
transform 1 0 1708 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1569
timestamp 1677677812
transform 1 0 1724 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1868
timestamp 1677677812
transform 1 0 1724 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1570
timestamp 1677677812
transform 1 0 1748 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1869
timestamp 1677677812
transform 1 0 1748 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1870
timestamp 1677677812
transform 1 0 1756 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1642
timestamp 1677677812
transform 1 0 1780 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_1871
timestamp 1677677812
transform 1 0 1796 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1670
timestamp 1677677812
transform 1 0 1796 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1513
timestamp 1677677812
transform 1 0 1812 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1514
timestamp 1677677812
transform 1 0 1836 0 1 3865
box -3 -3 3 3
use M2_M1  M2_M1_1872
timestamp 1677677812
transform 1 0 1844 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1873
timestamp 1677677812
transform 1 0 1860 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1972
timestamp 1677677812
transform 1 0 1828 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1973
timestamp 1677677812
transform 1 0 1836 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1974
timestamp 1677677812
transform 1 0 1852 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1643
timestamp 1677677812
transform 1 0 1852 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1515
timestamp 1677677812
transform 1 0 1924 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1516
timestamp 1677677812
transform 1 0 1940 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1520
timestamp 1677677812
transform 1 0 1932 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1874
timestamp 1677677812
transform 1 0 1884 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1875
timestamp 1677677812
transform 1 0 1892 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1876
timestamp 1677677812
transform 1 0 1940 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1619
timestamp 1677677812
transform 1 0 1932 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1975
timestamp 1677677812
transform 1 0 1972 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1877
timestamp 1677677812
transform 1 0 1988 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1598
timestamp 1677677812
transform 1 0 2004 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1521
timestamp 1677677812
transform 1 0 2036 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1878
timestamp 1677677812
transform 1 0 2028 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1976
timestamp 1677677812
transform 1 0 2004 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1977
timestamp 1677677812
transform 1 0 2020 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1644
timestamp 1677677812
transform 1 0 1996 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1671
timestamp 1677677812
transform 1 0 1988 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1620
timestamp 1677677812
transform 1 0 2028 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1978
timestamp 1677677812
transform 1 0 2036 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1645
timestamp 1677677812
transform 1 0 2036 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1621
timestamp 1677677812
transform 1 0 2052 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1622
timestamp 1677677812
transform 1 0 2068 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1879
timestamp 1677677812
transform 1 0 2132 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1979
timestamp 1677677812
transform 1 0 2084 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1672
timestamp 1677677812
transform 1 0 2124 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1880
timestamp 1677677812
transform 1 0 2180 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1881
timestamp 1677677812
transform 1 0 2188 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1673
timestamp 1677677812
transform 1 0 2172 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1674
timestamp 1677677812
transform 1 0 2196 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1980
timestamp 1677677812
transform 1 0 2252 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1675
timestamp 1677677812
transform 1 0 2268 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1534
timestamp 1677677812
transform 1 0 2284 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1571
timestamp 1677677812
transform 1 0 2292 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1535
timestamp 1677677812
transform 1 0 2324 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1882
timestamp 1677677812
transform 1 0 2292 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1883
timestamp 1677677812
transform 1 0 2308 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1599
timestamp 1677677812
transform 1 0 2316 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1884
timestamp 1677677812
transform 1 0 2324 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1600
timestamp 1677677812
transform 1 0 2332 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1981
timestamp 1677677812
transform 1 0 2292 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1982
timestamp 1677677812
transform 1 0 2316 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1983
timestamp 1677677812
transform 1 0 2324 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1676
timestamp 1677677812
transform 1 0 2316 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1885
timestamp 1677677812
transform 1 0 2356 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1886
timestamp 1677677812
transform 1 0 2380 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1887
timestamp 1677677812
transform 1 0 2428 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1601
timestamp 1677677812
transform 1 0 2460 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1888
timestamp 1677677812
transform 1 0 2476 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1984
timestamp 1677677812
transform 1 0 2460 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1572
timestamp 1677677812
transform 1 0 2500 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1889
timestamp 1677677812
transform 1 0 2500 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1602
timestamp 1677677812
transform 1 0 2508 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1522
timestamp 1677677812
transform 1 0 2548 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1536
timestamp 1677677812
transform 1 0 2524 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1890
timestamp 1677677812
transform 1 0 2540 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1603
timestamp 1677677812
transform 1 0 2548 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1985
timestamp 1677677812
transform 1 0 2524 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1986
timestamp 1677677812
transform 1 0 2532 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1987
timestamp 1677677812
transform 1 0 2548 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1988
timestamp 1677677812
transform 1 0 2556 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1891
timestamp 1677677812
transform 1 0 2572 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1573
timestamp 1677677812
transform 1 0 2612 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1892
timestamp 1677677812
transform 1 0 2612 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1574
timestamp 1677677812
transform 1 0 2652 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1893
timestamp 1677677812
transform 1 0 2652 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1604
timestamp 1677677812
transform 1 0 2700 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1894
timestamp 1677677812
transform 1 0 2708 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1989
timestamp 1677677812
transform 1 0 2628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1990
timestamp 1677677812
transform 1 0 2716 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1646
timestamp 1677677812
transform 1 0 2628 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1647
timestamp 1677677812
transform 1 0 2660 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1648
timestamp 1677677812
transform 1 0 2708 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1537
timestamp 1677677812
transform 1 0 2732 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1895
timestamp 1677677812
transform 1 0 2756 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1677
timestamp 1677677812
transform 1 0 2756 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1829
timestamp 1677677812
transform 1 0 2788 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1605
timestamp 1677677812
transform 1 0 2788 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2037
timestamp 1677677812
transform 1 0 2780 0 1 3795
box -2 -2 2 2
use M3_M2  M3_M2_1557
timestamp 1677677812
transform 1 0 2804 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1991
timestamp 1677677812
transform 1 0 2796 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1992
timestamp 1677677812
transform 1 0 2804 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1993
timestamp 1677677812
transform 1 0 2812 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1678
timestamp 1677677812
transform 1 0 2788 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1649
timestamp 1677677812
transform 1 0 2812 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1523
timestamp 1677677812
transform 1 0 2828 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1896
timestamp 1677677812
transform 1 0 2828 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1575
timestamp 1677677812
transform 1 0 2844 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1897
timestamp 1677677812
transform 1 0 2844 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1994
timestamp 1677677812
transform 1 0 2860 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1524
timestamp 1677677812
transform 1 0 2876 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1830
timestamp 1677677812
transform 1 0 2884 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1650
timestamp 1677677812
transform 1 0 2884 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1576
timestamp 1677677812
transform 1 0 2916 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1898
timestamp 1677677812
transform 1 0 2908 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1606
timestamp 1677677812
transform 1 0 2924 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1995
timestamp 1677677812
transform 1 0 2916 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1996
timestamp 1677677812
transform 1 0 2924 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1679
timestamp 1677677812
transform 1 0 2908 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1831
timestamp 1677677812
transform 1 0 2940 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1680
timestamp 1677677812
transform 1 0 2932 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1832
timestamp 1677677812
transform 1 0 2956 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1899
timestamp 1677677812
transform 1 0 2972 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1651
timestamp 1677677812
transform 1 0 2956 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1681
timestamp 1677677812
transform 1 0 2972 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1538
timestamp 1677677812
transform 1 0 2996 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1525
timestamp 1677677812
transform 1 0 3012 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1607
timestamp 1677677812
transform 1 0 3004 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1577
timestamp 1677677812
transform 1 0 3020 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1578
timestamp 1677677812
transform 1 0 3044 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1900
timestamp 1677677812
transform 1 0 3020 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1901
timestamp 1677677812
transform 1 0 3044 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1997
timestamp 1677677812
transform 1 0 3004 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1998
timestamp 1677677812
transform 1 0 3012 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1999
timestamp 1677677812
transform 1 0 3028 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1623
timestamp 1677677812
transform 1 0 3036 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_2000
timestamp 1677677812
transform 1 0 3044 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2001
timestamp 1677677812
transform 1 0 3052 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1652
timestamp 1677677812
transform 1 0 3028 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1608
timestamp 1677677812
transform 1 0 3068 0 1 3815
box -3 -3 3 3
use M3_M2  M3_M2_1526
timestamp 1677677812
transform 1 0 3108 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1579
timestamp 1677677812
transform 1 0 3132 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1902
timestamp 1677677812
transform 1 0 3108 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2002
timestamp 1677677812
transform 1 0 3156 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1653
timestamp 1677677812
transform 1 0 3108 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1580
timestamp 1677677812
transform 1 0 3172 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1903
timestamp 1677677812
transform 1 0 3172 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1527
timestamp 1677677812
transform 1 0 3236 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1539
timestamp 1677677812
transform 1 0 3228 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1904
timestamp 1677677812
transform 1 0 3228 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2003
timestamp 1677677812
transform 1 0 3204 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2004
timestamp 1677677812
transform 1 0 3220 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2005
timestamp 1677677812
transform 1 0 3236 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1654
timestamp 1677677812
transform 1 0 3204 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1655
timestamp 1677677812
transform 1 0 3268 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1540
timestamp 1677677812
transform 1 0 3284 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1905
timestamp 1677677812
transform 1 0 3284 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2006
timestamp 1677677812
transform 1 0 3300 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2007
timestamp 1677677812
transform 1 0 3340 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1682
timestamp 1677677812
transform 1 0 3364 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1656
timestamp 1677677812
transform 1 0 3380 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1657
timestamp 1677677812
transform 1 0 3404 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1541
timestamp 1677677812
transform 1 0 3476 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1581
timestamp 1677677812
transform 1 0 3460 0 1 3825
box -3 -3 3 3
use M3_M2  M3_M2_1582
timestamp 1677677812
transform 1 0 3484 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1906
timestamp 1677677812
transform 1 0 3452 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1907
timestamp 1677677812
transform 1 0 3468 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2008
timestamp 1677677812
transform 1 0 3460 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1683
timestamp 1677677812
transform 1 0 3468 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1908
timestamp 1677677812
transform 1 0 3516 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1542
timestamp 1677677812
transform 1 0 3540 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1909
timestamp 1677677812
transform 1 0 3588 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1910
timestamp 1677677812
transform 1 0 3628 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1911
timestamp 1677677812
transform 1 0 3644 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2009
timestamp 1677677812
transform 1 0 3612 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2010
timestamp 1677677812
transform 1 0 3620 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2011
timestamp 1677677812
transform 1 0 3636 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2012
timestamp 1677677812
transform 1 0 3652 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1517
timestamp 1677677812
transform 1 0 3764 0 1 3865
box -3 -3 3 3
use M3_M2  M3_M2_1518
timestamp 1677677812
transform 1 0 3844 0 1 3865
box -3 -3 3 3
use M2_M1  M2_M1_1912
timestamp 1677677812
transform 1 0 3764 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1913
timestamp 1677677812
transform 1 0 3820 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2013
timestamp 1677677812
transform 1 0 3844 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1658
timestamp 1677677812
transform 1 0 3844 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1543
timestamp 1677677812
transform 1 0 3860 0 1 3845
box -3 -3 3 3
use M3_M2  M3_M2_1684
timestamp 1677677812
transform 1 0 3820 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1685
timestamp 1677677812
transform 1 0 3852 0 1 3785
box -3 -3 3 3
use M2_M1  M2_M1_1914
timestamp 1677677812
transform 1 0 3868 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1915
timestamp 1677677812
transform 1 0 3876 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1916
timestamp 1677677812
transform 1 0 3908 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2014
timestamp 1677677812
transform 1 0 3916 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2015
timestamp 1677677812
transform 1 0 3924 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1659
timestamp 1677677812
transform 1 0 3900 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1660
timestamp 1677677812
transform 1 0 3916 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1686
timestamp 1677677812
transform 1 0 3892 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1583
timestamp 1677677812
transform 1 0 3948 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1917
timestamp 1677677812
transform 1 0 3940 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1918
timestamp 1677677812
transform 1 0 3948 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1919
timestamp 1677677812
transform 1 0 3964 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2016
timestamp 1677677812
transform 1 0 3956 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1661
timestamp 1677677812
transform 1 0 3964 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1584
timestamp 1677677812
transform 1 0 3980 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1920
timestamp 1677677812
transform 1 0 3980 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2017
timestamp 1677677812
transform 1 0 3988 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2018
timestamp 1677677812
transform 1 0 3996 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1662
timestamp 1677677812
transform 1 0 3988 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1585
timestamp 1677677812
transform 1 0 4012 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1921
timestamp 1677677812
transform 1 0 4012 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1528
timestamp 1677677812
transform 1 0 4036 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_2019
timestamp 1677677812
transform 1 0 4036 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1529
timestamp 1677677812
transform 1 0 4052 0 1 3855
box -3 -3 3 3
use M2_M1  M2_M1_1922
timestamp 1677677812
transform 1 0 4068 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1609
timestamp 1677677812
transform 1 0 4076 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1923
timestamp 1677677812
transform 1 0 4084 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2020
timestamp 1677677812
transform 1 0 4060 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2021
timestamp 1677677812
transform 1 0 4076 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1663
timestamp 1677677812
transform 1 0 4076 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_2022
timestamp 1677677812
transform 1 0 4100 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1544
timestamp 1677677812
transform 1 0 4116 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1924
timestamp 1677677812
transform 1 0 4116 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1624
timestamp 1677677812
transform 1 0 4140 0 1 3805
box -3 -3 3 3
use M2_M1  M2_M1_1925
timestamp 1677677812
transform 1 0 4172 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2023
timestamp 1677677812
transform 1 0 4148 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2024
timestamp 1677677812
transform 1 0 4164 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2025
timestamp 1677677812
transform 1 0 4180 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1687
timestamp 1677677812
transform 1 0 4180 0 1 3785
box -3 -3 3 3
use M3_M2  M3_M2_1530
timestamp 1677677812
transform 1 0 4220 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1545
timestamp 1677677812
transform 1 0 4236 0 1 3845
box -3 -3 3 3
use M2_M1  M2_M1_1926
timestamp 1677677812
transform 1 0 4252 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1586
timestamp 1677677812
transform 1 0 4276 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1927
timestamp 1677677812
transform 1 0 4276 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1610
timestamp 1677677812
transform 1 0 4284 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2026
timestamp 1677677812
transform 1 0 4260 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2027
timestamp 1677677812
transform 1 0 4284 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1928
timestamp 1677677812
transform 1 0 4308 0 1 3815
box -2 -2 2 2
use M3_M2  M3_M2_1531
timestamp 1677677812
transform 1 0 4332 0 1 3855
box -3 -3 3 3
use M3_M2  M3_M2_1558
timestamp 1677677812
transform 1 0 4332 0 1 3835
box -3 -3 3 3
use M2_M1  M2_M1_1826
timestamp 1677677812
transform 1 0 4340 0 1 3835
box -2 -2 2 2
use M2_M1  M2_M1_1833
timestamp 1677677812
transform 1 0 4332 0 1 3825
box -2 -2 2 2
use M3_M2  M3_M2_1587
timestamp 1677677812
transform 1 0 4340 0 1 3825
box -3 -3 3 3
use M2_M1  M2_M1_1834
timestamp 1677677812
transform 1 0 4348 0 1 3825
box -2 -2 2 2
use M2_M1  M2_M1_1929
timestamp 1677677812
transform 1 0 4348 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1930
timestamp 1677677812
transform 1 0 4420 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1931
timestamp 1677677812
transform 1 0 4468 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2028
timestamp 1677677812
transform 1 0 4388 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1611
timestamp 1677677812
transform 1 0 4476 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_1932
timestamp 1677677812
transform 1 0 4548 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1933
timestamp 1677677812
transform 1 0 4604 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2029
timestamp 1677677812
transform 1 0 4516 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1625
timestamp 1677677812
transform 1 0 4556 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1626
timestamp 1677677812
transform 1 0 4596 0 1 3805
box -3 -3 3 3
use M3_M2  M3_M2_1664
timestamp 1677677812
transform 1 0 4516 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1665
timestamp 1677677812
transform 1 0 4596 0 1 3795
box -3 -3 3 3
use M3_M2  M3_M2_1612
timestamp 1677677812
transform 1 0 4612 0 1 3815
box -3 -3 3 3
use M2_M1  M2_M1_2030
timestamp 1677677812
transform 1 0 4612 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1934
timestamp 1677677812
transform 1 0 4636 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1935
timestamp 1677677812
transform 1 0 4652 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2031
timestamp 1677677812
transform 1 0 4628 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_2032
timestamp 1677677812
transform 1 0 4644 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1666
timestamp 1677677812
transform 1 0 4644 0 1 3795
box -3 -3 3 3
use M2_M1  M2_M1_2033
timestamp 1677677812
transform 1 0 4668 0 1 3805
box -2 -2 2 2
use M2_M1  M2_M1_1936
timestamp 1677677812
transform 1 0 4724 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_1937
timestamp 1677677812
transform 1 0 4780 0 1 3815
box -2 -2 2 2
use M2_M1  M2_M1_2034
timestamp 1677677812
transform 1 0 4700 0 1 3805
box -2 -2 2 2
use M3_M2  M3_M2_1667
timestamp 1677677812
transform 1 0 4724 0 1 3795
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_18
timestamp 1677677812
transform 1 0 48 0 1 3770
box -10 -3 10 3
use FILL  FILL_1705
timestamp 1677677812
transform 1 0 72 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_132
timestamp 1677677812
transform 1 0 80 0 1 3770
box -8 -3 104 105
use FILL  FILL_1707
timestamp 1677677812
transform 1 0 176 0 1 3770
box -8 -3 16 105
use FILL  FILL_1708
timestamp 1677677812
transform 1 0 184 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_84
timestamp 1677677812
transform 1 0 192 0 1 3770
box -8 -3 46 105
use FILL  FILL_1709
timestamp 1677677812
transform 1 0 232 0 1 3770
box -8 -3 16 105
use FILL  FILL_1721
timestamp 1677677812
transform 1 0 240 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1688
timestamp 1677677812
transform 1 0 260 0 1 3775
box -3 -3 3 3
use INVX2  INVX2_151
timestamp 1677677812
transform -1 0 264 0 1 3770
box -9 -3 26 105
use FILL  FILL_1722
timestamp 1677677812
transform 1 0 264 0 1 3770
box -8 -3 16 105
use FILL  FILL_1723
timestamp 1677677812
transform 1 0 272 0 1 3770
box -8 -3 16 105
use FILL  FILL_1724
timestamp 1677677812
transform 1 0 280 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_86
timestamp 1677677812
transform -1 0 328 0 1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_133
timestamp 1677677812
transform 1 0 328 0 1 3770
box -8 -3 104 105
use INVX2  INVX2_152
timestamp 1677677812
transform -1 0 440 0 1 3770
box -9 -3 26 105
use FILL  FILL_1725
timestamp 1677677812
transform 1 0 440 0 1 3770
box -8 -3 16 105
use FILL  FILL_1726
timestamp 1677677812
transform 1 0 448 0 1 3770
box -8 -3 16 105
use FILL  FILL_1727
timestamp 1677677812
transform 1 0 456 0 1 3770
box -8 -3 16 105
use FILL  FILL_1728
timestamp 1677677812
transform 1 0 464 0 1 3770
box -8 -3 16 105
use FILL  FILL_1729
timestamp 1677677812
transform 1 0 472 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_87
timestamp 1677677812
transform 1 0 480 0 1 3770
box -8 -3 46 105
use FILL  FILL_1730
timestamp 1677677812
transform 1 0 520 0 1 3770
box -8 -3 16 105
use FILL  FILL_1731
timestamp 1677677812
transform 1 0 528 0 1 3770
box -8 -3 16 105
use FILL  FILL_1732
timestamp 1677677812
transform 1 0 536 0 1 3770
box -8 -3 16 105
use FILL  FILL_1733
timestamp 1677677812
transform 1 0 544 0 1 3770
box -8 -3 16 105
use FILL  FILL_1734
timestamp 1677677812
transform 1 0 552 0 1 3770
box -8 -3 16 105
use FILL  FILL_1735
timestamp 1677677812
transform 1 0 560 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_84
timestamp 1677677812
transform -1 0 608 0 1 3770
box -8 -3 46 105
use FILL  FILL_1736
timestamp 1677677812
transform 1 0 608 0 1 3770
box -8 -3 16 105
use FILL  FILL_1748
timestamp 1677677812
transform 1 0 616 0 1 3770
box -8 -3 16 105
use FILL  FILL_1750
timestamp 1677677812
transform 1 0 624 0 1 3770
box -8 -3 16 105
use FILL  FILL_1752
timestamp 1677677812
transform 1 0 632 0 1 3770
box -8 -3 16 105
use FILL  FILL_1753
timestamp 1677677812
transform 1 0 640 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_89
timestamp 1677677812
transform 1 0 648 0 1 3770
box -8 -3 46 105
use FILL  FILL_1754
timestamp 1677677812
transform 1 0 688 0 1 3770
box -8 -3 16 105
use FILL  FILL_1758
timestamp 1677677812
transform 1 0 696 0 1 3770
box -8 -3 16 105
use FILL  FILL_1760
timestamp 1677677812
transform 1 0 704 0 1 3770
box -8 -3 16 105
use FILL  FILL_1762
timestamp 1677677812
transform 1 0 712 0 1 3770
box -8 -3 16 105
use FILL  FILL_1764
timestamp 1677677812
transform 1 0 720 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_136
timestamp 1677677812
transform -1 0 824 0 1 3770
box -8 -3 104 105
use FILL  FILL_1765
timestamp 1677677812
transform 1 0 824 0 1 3770
box -8 -3 16 105
use FILL  FILL_1766
timestamp 1677677812
transform 1 0 832 0 1 3770
box -8 -3 16 105
use FILL  FILL_1767
timestamp 1677677812
transform 1 0 840 0 1 3770
box -8 -3 16 105
use FILL  FILL_1768
timestamp 1677677812
transform 1 0 848 0 1 3770
box -8 -3 16 105
use FILL  FILL_1769
timestamp 1677677812
transform 1 0 856 0 1 3770
box -8 -3 16 105
use FILL  FILL_1770
timestamp 1677677812
transform 1 0 864 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_91
timestamp 1677677812
transform 1 0 872 0 1 3770
box -8 -3 46 105
use M3_M2  M3_M2_1689
timestamp 1677677812
transform 1 0 924 0 1 3775
box -3 -3 3 3
use FILL  FILL_1771
timestamp 1677677812
transform 1 0 912 0 1 3770
box -8 -3 16 105
use FILL  FILL_1779
timestamp 1677677812
transform 1 0 920 0 1 3770
box -8 -3 16 105
use FILL  FILL_1781
timestamp 1677677812
transform 1 0 928 0 1 3770
box -8 -3 16 105
use FILL  FILL_1783
timestamp 1677677812
transform 1 0 936 0 1 3770
box -8 -3 16 105
use FILL  FILL_1785
timestamp 1677677812
transform 1 0 944 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_19
timestamp 1677677812
transform 1 0 952 0 1 3770
box -8 -3 32 105
use FILL  FILL_1786
timestamp 1677677812
transform 1 0 976 0 1 3770
box -8 -3 16 105
use FILL  FILL_1787
timestamp 1677677812
transform 1 0 984 0 1 3770
box -8 -3 16 105
use FILL  FILL_1788
timestamp 1677677812
transform 1 0 992 0 1 3770
box -8 -3 16 105
use FILL  FILL_1789
timestamp 1677677812
transform 1 0 1000 0 1 3770
box -8 -3 16 105
use FILL  FILL_1790
timestamp 1677677812
transform 1 0 1008 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_21
timestamp 1677677812
transform 1 0 1016 0 1 3770
box -8 -3 32 105
use FILL  FILL_1793
timestamp 1677677812
transform 1 0 1040 0 1 3770
box -8 -3 16 105
use FILL  FILL_1798
timestamp 1677677812
transform 1 0 1048 0 1 3770
box -8 -3 16 105
use FILL  FILL_1800
timestamp 1677677812
transform 1 0 1056 0 1 3770
box -8 -3 16 105
use FILL  FILL_1801
timestamp 1677677812
transform 1 0 1064 0 1 3770
box -8 -3 16 105
use FILL  FILL_1802
timestamp 1677677812
transform 1 0 1072 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_42
timestamp 1677677812
transform 1 0 1080 0 1 3770
box -8 -3 34 105
use FILL  FILL_1803
timestamp 1677677812
transform 1 0 1112 0 1 3770
box -8 -3 16 105
use FILL  FILL_1804
timestamp 1677677812
transform 1 0 1120 0 1 3770
box -8 -3 16 105
use FILL  FILL_1805
timestamp 1677677812
transform 1 0 1128 0 1 3770
box -8 -3 16 105
use FILL  FILL_1806
timestamp 1677677812
transform 1 0 1136 0 1 3770
box -8 -3 16 105
use FILL  FILL_1811
timestamp 1677677812
transform 1 0 1144 0 1 3770
box -8 -3 16 105
use FILL  FILL_1813
timestamp 1677677812
transform 1 0 1152 0 1 3770
box -8 -3 16 105
use FILL  FILL_1815
timestamp 1677677812
transform 1 0 1160 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_157
timestamp 1677677812
transform 1 0 1168 0 1 3770
box -9 -3 26 105
use FILL  FILL_1817
timestamp 1677677812
transform 1 0 1184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1818
timestamp 1677677812
transform 1 0 1192 0 1 3770
box -8 -3 16 105
use FILL  FILL_1819
timestamp 1677677812
transform 1 0 1200 0 1 3770
box -8 -3 16 105
use FILL  FILL_1820
timestamp 1677677812
transform 1 0 1208 0 1 3770
box -8 -3 16 105
use FILL  FILL_1821
timestamp 1677677812
transform 1 0 1216 0 1 3770
box -8 -3 16 105
use FILL  FILL_1824
timestamp 1677677812
transform 1 0 1224 0 1 3770
box -8 -3 16 105
use FILL  FILL_1826
timestamp 1677677812
transform 1 0 1232 0 1 3770
box -8 -3 16 105
use FILL  FILL_1828
timestamp 1677677812
transform 1 0 1240 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_44
timestamp 1677677812
transform -1 0 1280 0 1 3770
box -8 -3 34 105
use FILL  FILL_1829
timestamp 1677677812
transform 1 0 1280 0 1 3770
box -8 -3 16 105
use FILL  FILL_1834
timestamp 1677677812
transform 1 0 1288 0 1 3770
box -8 -3 16 105
use FILL  FILL_1835
timestamp 1677677812
transform 1 0 1296 0 1 3770
box -8 -3 16 105
use FILL  FILL_1836
timestamp 1677677812
transform 1 0 1304 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1690
timestamp 1677677812
transform 1 0 1324 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1691
timestamp 1677677812
transform 1 0 1412 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_138
timestamp 1677677812
transform 1 0 1312 0 1 3770
box -8 -3 104 105
use FILL  FILL_1837
timestamp 1677677812
transform 1 0 1408 0 1 3770
box -8 -3 16 105
use FILL  FILL_1844
timestamp 1677677812
transform 1 0 1416 0 1 3770
box -8 -3 16 105
use FILL  FILL_1846
timestamp 1677677812
transform 1 0 1424 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_160
timestamp 1677677812
transform 1 0 1432 0 1 3770
box -9 -3 26 105
use FILL  FILL_1848
timestamp 1677677812
transform 1 0 1448 0 1 3770
box -8 -3 16 105
use FILL  FILL_1849
timestamp 1677677812
transform 1 0 1456 0 1 3770
box -8 -3 16 105
use FILL  FILL_1850
timestamp 1677677812
transform 1 0 1464 0 1 3770
box -8 -3 16 105
use FILL  FILL_1851
timestamp 1677677812
transform 1 0 1472 0 1 3770
box -8 -3 16 105
use FILL  FILL_1852
timestamp 1677677812
transform 1 0 1480 0 1 3770
box -8 -3 16 105
use FILL  FILL_1853
timestamp 1677677812
transform 1 0 1488 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_86
timestamp 1677677812
transform -1 0 1536 0 1 3770
box -8 -3 46 105
use FILL  FILL_1854
timestamp 1677677812
transform 1 0 1536 0 1 3770
box -8 -3 16 105
use FILL  FILL_1857
timestamp 1677677812
transform 1 0 1544 0 1 3770
box -8 -3 16 105
use FILL  FILL_1858
timestamp 1677677812
transform 1 0 1552 0 1 3770
box -8 -3 16 105
use FILL  FILL_1859
timestamp 1677677812
transform 1 0 1560 0 1 3770
box -8 -3 16 105
use FILL  FILL_1861
timestamp 1677677812
transform 1 0 1568 0 1 3770
box -8 -3 16 105
use FILL  FILL_1863
timestamp 1677677812
transform 1 0 1576 0 1 3770
box -8 -3 16 105
use FILL  FILL_1865
timestamp 1677677812
transform 1 0 1584 0 1 3770
box -8 -3 16 105
use FILL  FILL_1867
timestamp 1677677812
transform 1 0 1592 0 1 3770
box -8 -3 16 105
use FILL  FILL_1869
timestamp 1677677812
transform 1 0 1600 0 1 3770
box -8 -3 16 105
use FILL  FILL_1870
timestamp 1677677812
transform 1 0 1608 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1692
timestamp 1677677812
transform 1 0 1636 0 1 3775
box -3 -3 3 3
use INVX2  INVX2_162
timestamp 1677677812
transform -1 0 1632 0 1 3770
box -9 -3 26 105
use FILL  FILL_1871
timestamp 1677677812
transform 1 0 1632 0 1 3770
box -8 -3 16 105
use FILL  FILL_1872
timestamp 1677677812
transform 1 0 1640 0 1 3770
box -8 -3 16 105
use FILL  FILL_1873
timestamp 1677677812
transform 1 0 1648 0 1 3770
box -8 -3 16 105
use FILL  FILL_1876
timestamp 1677677812
transform 1 0 1656 0 1 3770
box -8 -3 16 105
use FILL  FILL_1878
timestamp 1677677812
transform 1 0 1664 0 1 3770
box -8 -3 16 105
use FILL  FILL_1880
timestamp 1677677812
transform 1 0 1672 0 1 3770
box -8 -3 16 105
use BUFX2  BUFX2_12
timestamp 1677677812
transform -1 0 1704 0 1 3770
box -5 -3 28 105
use FILL  FILL_1881
timestamp 1677677812
transform 1 0 1704 0 1 3770
box -8 -3 16 105
use FILL  FILL_1882
timestamp 1677677812
transform 1 0 1712 0 1 3770
box -8 -3 16 105
use FILL  FILL_1883
timestamp 1677677812
transform 1 0 1720 0 1 3770
box -8 -3 16 105
use BUFX2  BUFX2_13
timestamp 1677677812
transform -1 0 1752 0 1 3770
box -5 -3 28 105
use FILL  FILL_1884
timestamp 1677677812
transform 1 0 1752 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1693
timestamp 1677677812
transform 1 0 1772 0 1 3775
box -3 -3 3 3
use FILL  FILL_1885
timestamp 1677677812
transform 1 0 1760 0 1 3770
box -8 -3 16 105
use FILL  FILL_1886
timestamp 1677677812
transform 1 0 1768 0 1 3770
box -8 -3 16 105
use FILL  FILL_1887
timestamp 1677677812
transform 1 0 1776 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_163
timestamp 1677677812
transform -1 0 1800 0 1 3770
box -9 -3 26 105
use FILL  FILL_1888
timestamp 1677677812
transform 1 0 1800 0 1 3770
box -8 -3 16 105
use FILL  FILL_1892
timestamp 1677677812
transform 1 0 1808 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1694
timestamp 1677677812
transform 1 0 1828 0 1 3775
box -3 -3 3 3
use FILL  FILL_1894
timestamp 1677677812
transform 1 0 1816 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_93
timestamp 1677677812
transform 1 0 1824 0 1 3770
box -8 -3 46 105
use FILL  FILL_1895
timestamp 1677677812
transform 1 0 1864 0 1 3770
box -8 -3 16 105
use FILL  FILL_1896
timestamp 1677677812
transform 1 0 1872 0 1 3770
box -8 -3 16 105
use FILL  FILL_1897
timestamp 1677677812
transform 1 0 1880 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_141
timestamp 1677677812
transform -1 0 1984 0 1 3770
box -8 -3 104 105
use M3_M2  M3_M2_1695
timestamp 1677677812
transform 1 0 2004 0 1 3775
box -3 -3 3 3
use FILL  FILL_1898
timestamp 1677677812
transform 1 0 1984 0 1 3770
box -8 -3 16 105
use FILL  FILL_1899
timestamp 1677677812
transform 1 0 1992 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1696
timestamp 1677677812
transform 1 0 2028 0 1 3775
box -3 -3 3 3
use OAI22X1  OAI22X1_88
timestamp 1677677812
transform 1 0 2000 0 1 3770
box -8 -3 46 105
use FILL  FILL_1900
timestamp 1677677812
transform 1 0 2040 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1697
timestamp 1677677812
transform 1 0 2060 0 1 3775
box -3 -3 3 3
use FILL  FILL_1901
timestamp 1677677812
transform 1 0 2048 0 1 3770
box -8 -3 16 105
use FILL  FILL_1902
timestamp 1677677812
transform 1 0 2056 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1698
timestamp 1677677812
transform 1 0 2076 0 1 3775
box -3 -3 3 3
use FILL  FILL_1903
timestamp 1677677812
transform 1 0 2064 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_142
timestamp 1677677812
transform 1 0 2072 0 1 3770
box -8 -3 104 105
use FILL  FILL_1904
timestamp 1677677812
transform 1 0 2168 0 1 3770
box -8 -3 16 105
use FILL  FILL_1905
timestamp 1677677812
transform 1 0 2176 0 1 3770
box -8 -3 16 105
use FILL  FILL_1906
timestamp 1677677812
transform 1 0 2184 0 1 3770
box -8 -3 16 105
use FILL  FILL_1907
timestamp 1677677812
transform 1 0 2192 0 1 3770
box -8 -3 16 105
use FILL  FILL_1916
timestamp 1677677812
transform 1 0 2200 0 1 3770
box -8 -3 16 105
use FILL  FILL_1918
timestamp 1677677812
transform 1 0 2208 0 1 3770
box -8 -3 16 105
use FILL  FILL_1920
timestamp 1677677812
transform 1 0 2216 0 1 3770
box -8 -3 16 105
use FILL  FILL_1922
timestamp 1677677812
transform 1 0 2224 0 1 3770
box -8 -3 16 105
use FILL  FILL_1924
timestamp 1677677812
transform 1 0 2232 0 1 3770
box -8 -3 16 105
use FILL  FILL_1925
timestamp 1677677812
transform 1 0 2240 0 1 3770
box -8 -3 16 105
use FILL  FILL_1926
timestamp 1677677812
transform 1 0 2248 0 1 3770
box -8 -3 16 105
use FILL  FILL_1928
timestamp 1677677812
transform 1 0 2256 0 1 3770
box -8 -3 16 105
use FILL  FILL_1930
timestamp 1677677812
transform 1 0 2264 0 1 3770
box -8 -3 16 105
use FILL  FILL_1932
timestamp 1677677812
transform 1 0 2272 0 1 3770
box -8 -3 16 105
use FILL  FILL_1934
timestamp 1677677812
transform 1 0 2280 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_96
timestamp 1677677812
transform 1 0 2288 0 1 3770
box -8 -3 46 105
use FILL  FILL_1936
timestamp 1677677812
transform 1 0 2328 0 1 3770
box -8 -3 16 105
use FILL  FILL_1938
timestamp 1677677812
transform 1 0 2336 0 1 3770
box -8 -3 16 105
use FILL  FILL_1940
timestamp 1677677812
transform 1 0 2344 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_169
timestamp 1677677812
transform 1 0 2352 0 1 3770
box -9 -3 26 105
use FILL  FILL_1942
timestamp 1677677812
transform 1 0 2368 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_145
timestamp 1677677812
transform -1 0 2472 0 1 3770
box -8 -3 104 105
use BUFX2  BUFX2_14
timestamp 1677677812
transform 1 0 2472 0 1 3770
box -5 -3 28 105
use FILL  FILL_1943
timestamp 1677677812
transform 1 0 2496 0 1 3770
box -8 -3 16 105
use FILL  FILL_1951
timestamp 1677677812
transform 1 0 2504 0 1 3770
box -8 -3 16 105
use FILL  FILL_1953
timestamp 1677677812
transform 1 0 2512 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_97
timestamp 1677677812
transform 1 0 2520 0 1 3770
box -8 -3 46 105
use FILL  FILL_1955
timestamp 1677677812
transform 1 0 2560 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_170
timestamp 1677677812
transform 1 0 2568 0 1 3770
box -9 -3 26 105
use FILL  FILL_1956
timestamp 1677677812
transform 1 0 2584 0 1 3770
box -8 -3 16 105
use FILL  FILL_1957
timestamp 1677677812
transform 1 0 2592 0 1 3770
box -8 -3 16 105
use FILL  FILL_1963
timestamp 1677677812
transform 1 0 2600 0 1 3770
box -8 -3 16 105
use FILL  FILL_1965
timestamp 1677677812
transform 1 0 2608 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_147
timestamp 1677677812
transform 1 0 2616 0 1 3770
box -8 -3 104 105
use FILL  FILL_1966
timestamp 1677677812
transform 1 0 2712 0 1 3770
box -8 -3 16 105
use FILL  FILL_1967
timestamp 1677677812
transform 1 0 2720 0 1 3770
box -8 -3 16 105
use FILL  FILL_1968
timestamp 1677677812
transform 1 0 2728 0 1 3770
box -8 -3 16 105
use FILL  FILL_1969
timestamp 1677677812
transform 1 0 2736 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_47
timestamp 1677677812
transform 1 0 2744 0 1 3770
box -8 -3 34 105
use FILL  FILL_1970
timestamp 1677677812
transform 1 0 2776 0 1 3770
box -8 -3 16 105
use FILL  FILL_1979
timestamp 1677677812
transform 1 0 2784 0 1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_23
timestamp 1677677812
transform 1 0 2792 0 1 3770
box -8 -3 32 105
use FILL  FILL_1981
timestamp 1677677812
transform 1 0 2816 0 1 3770
box -8 -3 16 105
use FILL  FILL_1983
timestamp 1677677812
transform 1 0 2824 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_48
timestamp 1677677812
transform 1 0 2832 0 1 3770
box -8 -3 34 105
use FILL  FILL_1985
timestamp 1677677812
transform 1 0 2864 0 1 3770
box -8 -3 16 105
use FILL  FILL_1988
timestamp 1677677812
transform 1 0 2872 0 1 3770
box -8 -3 16 105
use FILL  FILL_1990
timestamp 1677677812
transform 1 0 2880 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_49
timestamp 1677677812
transform -1 0 2920 0 1 3770
box -8 -3 34 105
use FILL  FILL_1991
timestamp 1677677812
transform 1 0 2920 0 1 3770
box -8 -3 16 105
use FILL  FILL_1996
timestamp 1677677812
transform 1 0 2928 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1699
timestamp 1677677812
transform 1 0 2948 0 1 3775
box -3 -3 3 3
use FILL  FILL_1997
timestamp 1677677812
transform 1 0 2936 0 1 3770
box -8 -3 16 105
use FILL  FILL_1998
timestamp 1677677812
transform 1 0 2944 0 1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_50
timestamp 1677677812
transform -1 0 2984 0 1 3770
box -8 -3 34 105
use FILL  FILL_1999
timestamp 1677677812
transform 1 0 2984 0 1 3770
box -8 -3 16 105
use FILL  FILL_2000
timestamp 1677677812
transform 1 0 2992 0 1 3770
box -8 -3 16 105
use FILL  FILL_2001
timestamp 1677677812
transform 1 0 3000 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_90
timestamp 1677677812
transform -1 0 3048 0 1 3770
box -8 -3 46 105
use FILL  FILL_2002
timestamp 1677677812
transform 1 0 3048 0 1 3770
box -8 -3 16 105
use FILL  FILL_2003
timestamp 1677677812
transform 1 0 3056 0 1 3770
box -8 -3 16 105
use FILL  FILL_2004
timestamp 1677677812
transform 1 0 3064 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_149
timestamp 1677677812
transform -1 0 3168 0 1 3770
box -8 -3 104 105
use FILL  FILL_2005
timestamp 1677677812
transform 1 0 3168 0 1 3770
box -8 -3 16 105
use FILL  FILL_2006
timestamp 1677677812
transform 1 0 3176 0 1 3770
box -8 -3 16 105
use FILL  FILL_2007
timestamp 1677677812
transform 1 0 3184 0 1 3770
box -8 -3 16 105
use FILL  FILL_2008
timestamp 1677677812
transform 1 0 3192 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_91
timestamp 1677677812
transform 1 0 3200 0 1 3770
box -8 -3 46 105
use FILL  FILL_2009
timestamp 1677677812
transform 1 0 3240 0 1 3770
box -8 -3 16 105
use FILL  FILL_2010
timestamp 1677677812
transform 1 0 3248 0 1 3770
box -8 -3 16 105
use FILL  FILL_2011
timestamp 1677677812
transform 1 0 3256 0 1 3770
box -8 -3 16 105
use FILL  FILL_2032
timestamp 1677677812
transform 1 0 3264 0 1 3770
box -8 -3 16 105
use FILL  FILL_2034
timestamp 1677677812
transform 1 0 3272 0 1 3770
box -8 -3 16 105
use FILL  FILL_2036
timestamp 1677677812
transform 1 0 3280 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_176
timestamp 1677677812
transform -1 0 3304 0 1 3770
box -9 -3 26 105
use FILL  FILL_2037
timestamp 1677677812
transform 1 0 3304 0 1 3770
box -8 -3 16 105
use FILL  FILL_2042
timestamp 1677677812
transform 1 0 3312 0 1 3770
box -8 -3 16 105
use FILL  FILL_2044
timestamp 1677677812
transform 1 0 3320 0 1 3770
box -8 -3 16 105
use FILL  FILL_2046
timestamp 1677677812
transform 1 0 3328 0 1 3770
box -8 -3 16 105
use FILL  FILL_2048
timestamp 1677677812
transform 1 0 3336 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1700
timestamp 1677677812
transform 1 0 3372 0 1 3775
box -3 -3 3 3
use INVX2  INVX2_177
timestamp 1677677812
transform 1 0 3344 0 1 3770
box -9 -3 26 105
use FILL  FILL_2049
timestamp 1677677812
transform 1 0 3360 0 1 3770
box -8 -3 16 105
use FILL  FILL_2050
timestamp 1677677812
transform 1 0 3368 0 1 3770
box -8 -3 16 105
use FILL  FILL_2051
timestamp 1677677812
transform 1 0 3376 0 1 3770
box -8 -3 16 105
use FILL  FILL_2054
timestamp 1677677812
transform 1 0 3384 0 1 3770
box -8 -3 16 105
use FILL  FILL_2056
timestamp 1677677812
transform 1 0 3392 0 1 3770
box -8 -3 16 105
use FILL  FILL_2058
timestamp 1677677812
transform 1 0 3400 0 1 3770
box -8 -3 16 105
use FILL  FILL_2060
timestamp 1677677812
transform 1 0 3408 0 1 3770
box -8 -3 16 105
use FILL  FILL_2062
timestamp 1677677812
transform 1 0 3416 0 1 3770
box -8 -3 16 105
use FILL  FILL_2064
timestamp 1677677812
transform 1 0 3424 0 1 3770
box -8 -3 16 105
use FILL  FILL_2065
timestamp 1677677812
transform 1 0 3432 0 1 3770
box -8 -3 16 105
use FILL  FILL_2066
timestamp 1677677812
transform 1 0 3440 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_99
timestamp 1677677812
transform 1 0 3448 0 1 3770
box -8 -3 46 105
use FILL  FILL_2067
timestamp 1677677812
transform 1 0 3488 0 1 3770
box -8 -3 16 105
use FILL  FILL_2068
timestamp 1677677812
transform 1 0 3496 0 1 3770
box -8 -3 16 105
use FILL  FILL_2069
timestamp 1677677812
transform 1 0 3504 0 1 3770
box -8 -3 16 105
use FILL  FILL_2070
timestamp 1677677812
transform 1 0 3512 0 1 3770
box -8 -3 16 105
use FILL  FILL_2071
timestamp 1677677812
transform 1 0 3520 0 1 3770
box -8 -3 16 105
use FILL  FILL_2073
timestamp 1677677812
transform 1 0 3528 0 1 3770
box -8 -3 16 105
use FILL  FILL_2075
timestamp 1677677812
transform 1 0 3536 0 1 3770
box -8 -3 16 105
use FILL  FILL_2077
timestamp 1677677812
transform 1 0 3544 0 1 3770
box -8 -3 16 105
use FILL  FILL_2079
timestamp 1677677812
transform 1 0 3552 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_178
timestamp 1677677812
transform -1 0 3576 0 1 3770
box -9 -3 26 105
use FILL  FILL_2080
timestamp 1677677812
transform 1 0 3576 0 1 3770
box -8 -3 16 105
use FILL  FILL_2081
timestamp 1677677812
transform 1 0 3584 0 1 3770
box -8 -3 16 105
use FILL  FILL_2085
timestamp 1677677812
transform 1 0 3592 0 1 3770
box -8 -3 16 105
use FILL  FILL_2087
timestamp 1677677812
transform 1 0 3600 0 1 3770
box -8 -3 16 105
use FILL  FILL_2089
timestamp 1677677812
transform 1 0 3608 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_92
timestamp 1677677812
transform -1 0 3656 0 1 3770
box -8 -3 46 105
use FILL  FILL_2090
timestamp 1677677812
transform 1 0 3656 0 1 3770
box -8 -3 16 105
use FILL  FILL_2091
timestamp 1677677812
transform 1 0 3664 0 1 3770
box -8 -3 16 105
use FILL  FILL_2092
timestamp 1677677812
transform 1 0 3672 0 1 3770
box -8 -3 16 105
use FILL  FILL_2093
timestamp 1677677812
transform 1 0 3680 0 1 3770
box -8 -3 16 105
use FILL  FILL_2094
timestamp 1677677812
transform 1 0 3688 0 1 3770
box -8 -3 16 105
use FILL  FILL_2095
timestamp 1677677812
transform 1 0 3696 0 1 3770
box -8 -3 16 105
use FILL  FILL_2096
timestamp 1677677812
transform 1 0 3704 0 1 3770
box -8 -3 16 105
use FILL  FILL_2097
timestamp 1677677812
transform 1 0 3712 0 1 3770
box -8 -3 16 105
use FILL  FILL_2098
timestamp 1677677812
transform 1 0 3720 0 1 3770
box -8 -3 16 105
use FILL  FILL_2099
timestamp 1677677812
transform 1 0 3728 0 1 3770
box -8 -3 16 105
use FILL  FILL_2104
timestamp 1677677812
transform 1 0 3736 0 1 3770
box -8 -3 16 105
use FILL  FILL_2106
timestamp 1677677812
transform 1 0 3744 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1701
timestamp 1677677812
transform 1 0 3764 0 1 3775
box -3 -3 3 3
use FILL  FILL_2108
timestamp 1677677812
transform 1 0 3752 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1702
timestamp 1677677812
transform 1 0 3788 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_153
timestamp 1677677812
transform -1 0 3856 0 1 3770
box -8 -3 104 105
use FILL  FILL_2109
timestamp 1677677812
transform 1 0 3856 0 1 3770
box -8 -3 16 105
use FILL  FILL_2110
timestamp 1677677812
transform 1 0 3864 0 1 3770
box -8 -3 16 105
use FILL  FILL_2111
timestamp 1677677812
transform 1 0 3872 0 1 3770
box -8 -3 16 105
use FILL  FILL_2119
timestamp 1677677812
transform 1 0 3880 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_100
timestamp 1677677812
transform -1 0 3928 0 1 3770
box -8 -3 46 105
use FILL  FILL_2120
timestamp 1677677812
transform 1 0 3928 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_94
timestamp 1677677812
transform 1 0 3936 0 1 3770
box -8 -3 46 105
use FILL  FILL_2128
timestamp 1677677812
transform 1 0 3976 0 1 3770
box -8 -3 16 105
use FILL  FILL_2129
timestamp 1677677812
transform 1 0 3984 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_182
timestamp 1677677812
transform 1 0 3992 0 1 3770
box -9 -3 26 105
use FILL  FILL_2130
timestamp 1677677812
transform 1 0 4008 0 1 3770
box -8 -3 16 105
use FILL  FILL_2131
timestamp 1677677812
transform 1 0 4016 0 1 3770
box -8 -3 16 105
use FILL  FILL_2132
timestamp 1677677812
transform 1 0 4024 0 1 3770
box -8 -3 16 105
use FILL  FILL_2133
timestamp 1677677812
transform 1 0 4032 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_95
timestamp 1677677812
transform 1 0 4040 0 1 3770
box -8 -3 46 105
use FILL  FILL_2134
timestamp 1677677812
transform 1 0 4080 0 1 3770
box -8 -3 16 105
use FILL  FILL_2142
timestamp 1677677812
transform 1 0 4088 0 1 3770
box -8 -3 16 105
use INVX2  INVX2_183
timestamp 1677677812
transform 1 0 4096 0 1 3770
box -9 -3 26 105
use FILL  FILL_2144
timestamp 1677677812
transform 1 0 4112 0 1 3770
box -8 -3 16 105
use FILL  FILL_2148
timestamp 1677677812
transform 1 0 4120 0 1 3770
box -8 -3 16 105
use FILL  FILL_2150
timestamp 1677677812
transform 1 0 4128 0 1 3770
box -8 -3 16 105
use FILL  FILL_2152
timestamp 1677677812
transform 1 0 4136 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_96
timestamp 1677677812
transform 1 0 4144 0 1 3770
box -8 -3 46 105
use FILL  FILL_2154
timestamp 1677677812
transform 1 0 4184 0 1 3770
box -8 -3 16 105
use FILL  FILL_2161
timestamp 1677677812
transform 1 0 4192 0 1 3770
box -8 -3 16 105
use FILL  FILL_2163
timestamp 1677677812
transform 1 0 4200 0 1 3770
box -8 -3 16 105
use FILL  FILL_2165
timestamp 1677677812
transform 1 0 4208 0 1 3770
box -8 -3 16 105
use FILL  FILL_2167
timestamp 1677677812
transform 1 0 4216 0 1 3770
box -8 -3 16 105
use FILL  FILL_2168
timestamp 1677677812
transform 1 0 4224 0 1 3770
box -8 -3 16 105
use FILL  FILL_2169
timestamp 1677677812
transform 1 0 4232 0 1 3770
box -8 -3 16 105
use FILL  FILL_2170
timestamp 1677677812
transform 1 0 4240 0 1 3770
box -8 -3 16 105
use FILL  FILL_2173
timestamp 1677677812
transform 1 0 4248 0 1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_101
timestamp 1677677812
transform -1 0 4296 0 1 3770
box -8 -3 46 105
use FILL  FILL_2174
timestamp 1677677812
transform 1 0 4296 0 1 3770
box -8 -3 16 105
use FILL  FILL_2182
timestamp 1677677812
transform 1 0 4304 0 1 3770
box -8 -3 16 105
use FILL  FILL_2184
timestamp 1677677812
transform 1 0 4312 0 1 3770
box -8 -3 16 105
use FILL  FILL_2186
timestamp 1677677812
transform 1 0 4320 0 1 3770
box -8 -3 16 105
use NAND3X1  NAND3X1_10
timestamp 1677677812
transform -1 0 4360 0 1 3770
box -8 -3 40 105
use FILL  FILL_2187
timestamp 1677677812
transform 1 0 4360 0 1 3770
box -8 -3 16 105
use FILL  FILL_2194
timestamp 1677677812
transform 1 0 4368 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_155
timestamp 1677677812
transform 1 0 4376 0 1 3770
box -8 -3 104 105
use FILL  FILL_2196
timestamp 1677677812
transform 1 0 4472 0 1 3770
box -8 -3 16 105
use FILL  FILL_2206
timestamp 1677677812
transform 1 0 4480 0 1 3770
box -8 -3 16 105
use FILL  FILL_2207
timestamp 1677677812
transform 1 0 4488 0 1 3770
box -8 -3 16 105
use FILL  FILL_2208
timestamp 1677677812
transform 1 0 4496 0 1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1703
timestamp 1677677812
transform 1 0 4532 0 1 3775
box -3 -3 3 3
use M3_M2  M3_M2_1704
timestamp 1677677812
transform 1 0 4580 0 1 3775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_156
timestamp 1677677812
transform 1 0 4504 0 1 3770
box -8 -3 104 105
use FILL  FILL_2209
timestamp 1677677812
transform 1 0 4600 0 1 3770
box -8 -3 16 105
use FILL  FILL_2210
timestamp 1677677812
transform 1 0 4608 0 1 3770
box -8 -3 16 105
use FILL  FILL_2211
timestamp 1677677812
transform 1 0 4616 0 1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_97
timestamp 1677677812
transform 1 0 4624 0 1 3770
box -8 -3 46 105
use FILL  FILL_2212
timestamp 1677677812
transform 1 0 4664 0 1 3770
box -8 -3 16 105
use FILL  FILL_2213
timestamp 1677677812
transform 1 0 4672 0 1 3770
box -8 -3 16 105
use FILL  FILL_2214
timestamp 1677677812
transform 1 0 4680 0 1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_157
timestamp 1677677812
transform 1 0 4688 0 1 3770
box -8 -3 104 105
use FILL  FILL_2215
timestamp 1677677812
transform 1 0 4784 0 1 3770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_19
timestamp 1677677812
transform 1 0 4819 0 1 3770
box -10 -3 10 3
use M3_M2  M3_M2_1723
timestamp 1677677812
transform 1 0 92 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2042
timestamp 1677677812
transform 1 0 92 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1813
timestamp 1677677812
transform 1 0 92 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2129
timestamp 1677677812
transform 1 0 108 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2130
timestamp 1677677812
transform 1 0 124 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1747
timestamp 1677677812
transform 1 0 172 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1774
timestamp 1677677812
transform 1 0 164 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2043
timestamp 1677677812
transform 1 0 172 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2044
timestamp 1677677812
transform 1 0 180 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2045
timestamp 1677677812
transform 1 0 196 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2131
timestamp 1677677812
transform 1 0 164 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2132
timestamp 1677677812
transform 1 0 188 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1793
timestamp 1677677812
transform 1 0 196 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1814
timestamp 1677677812
transform 1 0 188 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1748
timestamp 1677677812
transform 1 0 212 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2046
timestamp 1677677812
transform 1 0 220 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1775
timestamp 1677677812
transform 1 0 228 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2234
timestamp 1677677812
transform 1 0 220 0 1 3705
box -2 -2 2 2
use M2_M1  M2_M1_2047
timestamp 1677677812
transform 1 0 260 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2048
timestamp 1677677812
transform 1 0 276 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2133
timestamp 1677677812
transform 1 0 244 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2134
timestamp 1677677812
transform 1 0 252 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2135
timestamp 1677677812
transform 1 0 268 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1705
timestamp 1677677812
transform 1 0 332 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1724
timestamp 1677677812
transform 1 0 308 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1725
timestamp 1677677812
transform 1 0 340 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1749
timestamp 1677677812
transform 1 0 388 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2049
timestamp 1677677812
transform 1 0 308 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2136
timestamp 1677677812
transform 1 0 356 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2137
timestamp 1677677812
transform 1 0 388 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2138
timestamp 1677677812
transform 1 0 396 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1815
timestamp 1677677812
transform 1 0 356 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1816
timestamp 1677677812
transform 1 0 396 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2139
timestamp 1677677812
transform 1 0 428 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1706
timestamp 1677677812
transform 1 0 444 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1750
timestamp 1677677812
transform 1 0 468 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2050
timestamp 1677677812
transform 1 0 444 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2051
timestamp 1677677812
transform 1 0 452 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2052
timestamp 1677677812
transform 1 0 468 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1794
timestamp 1677677812
transform 1 0 452 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2140
timestamp 1677677812
transform 1 0 460 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1776
timestamp 1677677812
transform 1 0 492 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2141
timestamp 1677677812
transform 1 0 492 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1817
timestamp 1677677812
transform 1 0 492 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1707
timestamp 1677677812
transform 1 0 588 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1726
timestamp 1677677812
transform 1 0 516 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1727
timestamp 1677677812
transform 1 0 588 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2053
timestamp 1677677812
transform 1 0 516 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2142
timestamp 1677677812
transform 1 0 556 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2143
timestamp 1677677812
transform 1 0 604 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1728
timestamp 1677677812
transform 1 0 652 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1729
timestamp 1677677812
transform 1 0 668 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2054
timestamp 1677677812
transform 1 0 644 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2055
timestamp 1677677812
transform 1 0 668 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2056
timestamp 1677677812
transform 1 0 676 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2144
timestamp 1677677812
transform 1 0 636 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1795
timestamp 1677677812
transform 1 0 644 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2145
timestamp 1677677812
transform 1 0 652 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1796
timestamp 1677677812
transform 1 0 660 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2146
timestamp 1677677812
transform 1 0 668 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1797
timestamp 1677677812
transform 1 0 676 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1818
timestamp 1677677812
transform 1 0 668 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2147
timestamp 1677677812
transform 1 0 692 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1819
timestamp 1677677812
transform 1 0 684 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1730
timestamp 1677677812
transform 1 0 740 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2057
timestamp 1677677812
transform 1 0 740 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2148
timestamp 1677677812
transform 1 0 740 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2149
timestamp 1677677812
transform 1 0 772 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1798
timestamp 1677677812
transform 1 0 780 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1731
timestamp 1677677812
transform 1 0 876 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2058
timestamp 1677677812
transform 1 0 796 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1777
timestamp 1677677812
transform 1 0 844 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1799
timestamp 1677677812
transform 1 0 796 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1800
timestamp 1677677812
transform 1 0 820 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2059
timestamp 1677677812
transform 1 0 892 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2150
timestamp 1677677812
transform 1 0 836 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2151
timestamp 1677677812
transform 1 0 876 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2152
timestamp 1677677812
transform 1 0 892 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1820
timestamp 1677677812
transform 1 0 796 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1821
timestamp 1677677812
transform 1 0 884 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1856
timestamp 1677677812
transform 1 0 836 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1857
timestamp 1677677812
transform 1 0 892 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1732
timestamp 1677677812
transform 1 0 908 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2038
timestamp 1677677812
transform 1 0 924 0 1 3745
box -2 -2 2 2
use M3_M2  M3_M2_1733
timestamp 1677677812
transform 1 0 972 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1751
timestamp 1677677812
transform 1 0 964 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2060
timestamp 1677677812
transform 1 0 956 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2061
timestamp 1677677812
transform 1 0 972 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2153
timestamp 1677677812
transform 1 0 964 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2154
timestamp 1677677812
transform 1 0 972 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1822
timestamp 1677677812
transform 1 0 972 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1708
timestamp 1677677812
transform 1 0 1004 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1752
timestamp 1677677812
transform 1 0 1004 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2062
timestamp 1677677812
transform 1 0 1004 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2039
timestamp 1677677812
transform 1 0 1012 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2227
timestamp 1677677812
transform 1 0 1036 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1874
timestamp 1677677812
transform 1 0 1036 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1709
timestamp 1677677812
transform 1 0 1052 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2063
timestamp 1677677812
transform 1 0 1052 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1734
timestamp 1677677812
transform 1 0 1100 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2228
timestamp 1677677812
transform 1 0 1100 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2064
timestamp 1677677812
transform 1 0 1132 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2155
timestamp 1677677812
transform 1 0 1148 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1823
timestamp 1677677812
transform 1 0 1164 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1710
timestamp 1677677812
transform 1 0 1220 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2065
timestamp 1677677812
transform 1 0 1204 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2066
timestamp 1677677812
transform 1 0 1212 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2156
timestamp 1677677812
transform 1 0 1180 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2157
timestamp 1677677812
transform 1 0 1196 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1753
timestamp 1677677812
transform 1 0 1228 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2067
timestamp 1677677812
transform 1 0 1228 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2068
timestamp 1677677812
transform 1 0 1260 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1801
timestamp 1677677812
transform 1 0 1252 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1875
timestamp 1677677812
transform 1 0 1260 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2158
timestamp 1677677812
transform 1 0 1268 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1802
timestamp 1677677812
transform 1 0 1284 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2229
timestamp 1677677812
transform 1 0 1284 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1858
timestamp 1677677812
transform 1 0 1284 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1754
timestamp 1677677812
transform 1 0 1308 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1755
timestamp 1677677812
transform 1 0 1332 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1735
timestamp 1677677812
transform 1 0 1348 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2069
timestamp 1677677812
transform 1 0 1324 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2070
timestamp 1677677812
transform 1 0 1340 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2071
timestamp 1677677812
transform 1 0 1348 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2159
timestamp 1677677812
transform 1 0 1316 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1803
timestamp 1677677812
transform 1 0 1324 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2160
timestamp 1677677812
transform 1 0 1332 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1824
timestamp 1677677812
transform 1 0 1316 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1825
timestamp 1677677812
transform 1 0 1340 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2230
timestamp 1677677812
transform 1 0 1348 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1859
timestamp 1677677812
transform 1 0 1348 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2161
timestamp 1677677812
transform 1 0 1388 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1826
timestamp 1677677812
transform 1 0 1388 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2072
timestamp 1677677812
transform 1 0 1428 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1827
timestamp 1677677812
transform 1 0 1428 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1736
timestamp 1677677812
transform 1 0 1460 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1737
timestamp 1677677812
transform 1 0 1508 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1756
timestamp 1677677812
transform 1 0 1484 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2073
timestamp 1677677812
transform 1 0 1444 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2162
timestamp 1677677812
transform 1 0 1492 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1804
timestamp 1677677812
transform 1 0 1524 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1882
timestamp 1677677812
transform 1 0 1476 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1883
timestamp 1677677812
transform 1 0 1500 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1805
timestamp 1677677812
transform 1 0 1548 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1757
timestamp 1677677812
transform 1 0 1564 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2074
timestamp 1677677812
transform 1 0 1564 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2163
timestamp 1677677812
transform 1 0 1556 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1860
timestamp 1677677812
transform 1 0 1540 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2075
timestamp 1677677812
transform 1 0 1612 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2076
timestamp 1677677812
transform 1 0 1628 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2164
timestamp 1677677812
transform 1 0 1620 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2165
timestamp 1677677812
transform 1 0 1636 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1828
timestamp 1677677812
transform 1 0 1620 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1861
timestamp 1677677812
transform 1 0 1636 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1884
timestamp 1677677812
transform 1 0 1620 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2077
timestamp 1677677812
transform 1 0 1668 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1829
timestamp 1677677812
transform 1 0 1668 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1758
timestamp 1677677812
transform 1 0 1700 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1759
timestamp 1677677812
transform 1 0 1764 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2078
timestamp 1677677812
transform 1 0 1700 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1738
timestamp 1677677812
transform 1 0 1796 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2079
timestamp 1677677812
transform 1 0 1796 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2166
timestamp 1677677812
transform 1 0 1748 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2167
timestamp 1677677812
transform 1 0 1780 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2168
timestamp 1677677812
transform 1 0 1788 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1830
timestamp 1677677812
transform 1 0 1788 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2169
timestamp 1677677812
transform 1 0 1804 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1711
timestamp 1677677812
transform 1 0 1892 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1760
timestamp 1677677812
transform 1 0 1908 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2080
timestamp 1677677812
transform 1 0 1908 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2170
timestamp 1677677812
transform 1 0 1876 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1876
timestamp 1677677812
transform 1 0 1884 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1885
timestamp 1677677812
transform 1 0 1900 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2171
timestamp 1677677812
transform 1 0 1940 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2172
timestamp 1677677812
transform 1 0 1948 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1862
timestamp 1677677812
transform 1 0 1972 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1712
timestamp 1677677812
transform 1 0 1996 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1713
timestamp 1677677812
transform 1 0 2020 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1739
timestamp 1677677812
transform 1 0 2020 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1740
timestamp 1677677812
transform 1 0 2036 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1741
timestamp 1677677812
transform 1 0 2068 0 1 3755
box -3 -3 3 3
use M2_M1  M2_M1_2081
timestamp 1677677812
transform 1 0 1988 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2082
timestamp 1677677812
transform 1 0 1996 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2173
timestamp 1677677812
transform 1 0 1980 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1778
timestamp 1677677812
transform 1 0 2004 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1761
timestamp 1677677812
transform 1 0 2052 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1762
timestamp 1677677812
transform 1 0 2084 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2083
timestamp 1677677812
transform 1 0 2012 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2084
timestamp 1677677812
transform 1 0 2020 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2085
timestamp 1677677812
transform 1 0 2028 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2086
timestamp 1677677812
transform 1 0 2052 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1763
timestamp 1677677812
transform 1 0 2156 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1764
timestamp 1677677812
transform 1 0 2180 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2087
timestamp 1677677812
transform 1 0 2148 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2088
timestamp 1677677812
transform 1 0 2156 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2089
timestamp 1677677812
transform 1 0 2164 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2090
timestamp 1677677812
transform 1 0 2180 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2174
timestamp 1677677812
transform 1 0 2004 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2175
timestamp 1677677812
transform 1 0 2028 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2176
timestamp 1677677812
transform 1 0 2036 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2177
timestamp 1677677812
transform 1 0 2100 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2178
timestamp 1677677812
transform 1 0 2132 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2179
timestamp 1677677812
transform 1 0 2140 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1863
timestamp 1677677812
transform 1 0 1996 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1864
timestamp 1677677812
transform 1 0 2020 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1886
timestamp 1677677812
transform 1 0 2100 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1887
timestamp 1677677812
transform 1 0 2140 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1779
timestamp 1677677812
transform 1 0 2188 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2180
timestamp 1677677812
transform 1 0 2172 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2181
timestamp 1677677812
transform 1 0 2188 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1831
timestamp 1677677812
transform 1 0 2172 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1832
timestamp 1677677812
transform 1 0 2196 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1877
timestamp 1677677812
transform 1 0 2188 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2091
timestamp 1677677812
transform 1 0 2236 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1765
timestamp 1677677812
transform 1 0 2252 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2092
timestamp 1677677812
transform 1 0 2252 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2182
timestamp 1677677812
transform 1 0 2244 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1833
timestamp 1677677812
transform 1 0 2236 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1878
timestamp 1677677812
transform 1 0 2252 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2183
timestamp 1677677812
transform 1 0 2260 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2184
timestamp 1677677812
transform 1 0 2276 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1766
timestamp 1677677812
transform 1 0 2308 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2093
timestamp 1677677812
transform 1 0 2308 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2185
timestamp 1677677812
transform 1 0 2316 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2094
timestamp 1677677812
transform 1 0 2332 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1780
timestamp 1677677812
transform 1 0 2356 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1834
timestamp 1677677812
transform 1 0 2356 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1781
timestamp 1677677812
transform 1 0 2404 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2095
timestamp 1677677812
transform 1 0 2452 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2186
timestamp 1677677812
transform 1 0 2404 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1865
timestamp 1677677812
transform 1 0 2428 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1879
timestamp 1677677812
transform 1 0 2452 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2187
timestamp 1677677812
transform 1 0 2468 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1866
timestamp 1677677812
transform 1 0 2468 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2096
timestamp 1677677812
transform 1 0 2532 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1782
timestamp 1677677812
transform 1 0 2548 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2097
timestamp 1677677812
transform 1 0 2564 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1783
timestamp 1677677812
transform 1 0 2572 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2098
timestamp 1677677812
transform 1 0 2580 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2188
timestamp 1677677812
transform 1 0 2572 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1835
timestamp 1677677812
transform 1 0 2572 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1867
timestamp 1677677812
transform 1 0 2580 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1888
timestamp 1677677812
transform 1 0 2572 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2099
timestamp 1677677812
transform 1 0 2596 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1784
timestamp 1677677812
transform 1 0 2604 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2189
timestamp 1677677812
transform 1 0 2604 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1836
timestamp 1677677812
transform 1 0 2596 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2190
timestamp 1677677812
transform 1 0 2644 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1837
timestamp 1677677812
transform 1 0 2644 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2100
timestamp 1677677812
transform 1 0 2660 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1714
timestamp 1677677812
transform 1 0 2748 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2040
timestamp 1677677812
transform 1 0 2748 0 1 3745
box -2 -2 2 2
use M2_M1  M2_M1_2191
timestamp 1677677812
transform 1 0 2684 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2192
timestamp 1677677812
transform 1 0 2740 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1838
timestamp 1677677812
transform 1 0 2684 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1868
timestamp 1677677812
transform 1 0 2740 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1869
timestamp 1677677812
transform 1 0 2780 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2193
timestamp 1677677812
transform 1 0 2812 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2041
timestamp 1677677812
transform 1 0 2828 0 1 3745
box -2 -2 2 2
use M3_M2  M3_M2_1785
timestamp 1677677812
transform 1 0 2828 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1767
timestamp 1677677812
transform 1 0 2844 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2101
timestamp 1677677812
transform 1 0 2844 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1839
timestamp 1677677812
transform 1 0 2844 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1880
timestamp 1677677812
transform 1 0 2844 0 1 3695
box -3 -3 3 3
use M3_M2  M3_M2_1768
timestamp 1677677812
transform 1 0 2868 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2194
timestamp 1677677812
transform 1 0 2860 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2102
timestamp 1677677812
transform 1 0 2876 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1870
timestamp 1677677812
transform 1 0 2876 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1881
timestamp 1677677812
transform 1 0 2868 0 1 3695
box -3 -3 3 3
use M2_M1  M2_M1_2103
timestamp 1677677812
transform 1 0 2892 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2195
timestamp 1677677812
transform 1 0 2908 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2104
timestamp 1677677812
transform 1 0 2948 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1889
timestamp 1677677812
transform 1 0 2948 0 1 3685
box -3 -3 3 3
use M2_M1  M2_M1_2231
timestamp 1677677812
transform 1 0 2956 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2105
timestamp 1677677812
transform 1 0 2996 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2196
timestamp 1677677812
transform 1 0 2972 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2197
timestamp 1677677812
transform 1 0 2988 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2198
timestamp 1677677812
transform 1 0 3020 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2106
timestamp 1677677812
transform 1 0 3052 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2107
timestamp 1677677812
transform 1 0 3076 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2199
timestamp 1677677812
transform 1 0 3068 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1806
timestamp 1677677812
transform 1 0 3148 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2108
timestamp 1677677812
transform 1 0 3172 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2200
timestamp 1677677812
transform 1 0 3196 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2201
timestamp 1677677812
transform 1 0 3252 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1840
timestamp 1677677812
transform 1 0 3284 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2232
timestamp 1677677812
transform 1 0 3332 0 1 3715
box -2 -2 2 2
use M2_M1  M2_M1_2202
timestamp 1677677812
transform 1 0 3364 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2235
timestamp 1677677812
transform 1 0 3372 0 1 3705
box -2 -2 2 2
use M3_M2  M3_M2_1786
timestamp 1677677812
transform 1 0 3388 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1807
timestamp 1677677812
transform 1 0 3412 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2233
timestamp 1677677812
transform 1 0 3412 0 1 3715
box -2 -2 2 2
use M3_M2  M3_M2_1841
timestamp 1677677812
transform 1 0 3420 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1715
timestamp 1677677812
transform 1 0 3468 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1769
timestamp 1677677812
transform 1 0 3452 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1770
timestamp 1677677812
transform 1 0 3476 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2109
timestamp 1677677812
transform 1 0 3436 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1787
timestamp 1677677812
transform 1 0 3516 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2203
timestamp 1677677812
transform 1 0 3460 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2204
timestamp 1677677812
transform 1 0 3516 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2205
timestamp 1677677812
transform 1 0 3532 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1842
timestamp 1677677812
transform 1 0 3532 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1716
timestamp 1677677812
transform 1 0 3652 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1742
timestamp 1677677812
transform 1 0 3652 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1743
timestamp 1677677812
transform 1 0 3700 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1744
timestamp 1677677812
transform 1 0 3716 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1788
timestamp 1677677812
transform 1 0 3636 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1789
timestamp 1677677812
transform 1 0 3668 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2110
timestamp 1677677812
transform 1 0 3716 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1843
timestamp 1677677812
transform 1 0 3628 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2206
timestamp 1677677812
transform 1 0 3668 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1844
timestamp 1677677812
transform 1 0 3644 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1845
timestamp 1677677812
transform 1 0 3716 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2111
timestamp 1677677812
transform 1 0 3740 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2112
timestamp 1677677812
transform 1 0 3788 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2207
timestamp 1677677812
transform 1 0 3780 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2208
timestamp 1677677812
transform 1 0 3788 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2113
timestamp 1677677812
transform 1 0 3820 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1846
timestamp 1677677812
transform 1 0 3820 0 1 3715
box -3 -3 3 3
use M2_M1  M2_M1_2209
timestamp 1677677812
transform 1 0 3828 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1717
timestamp 1677677812
transform 1 0 3868 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2114
timestamp 1677677812
transform 1 0 3852 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2115
timestamp 1677677812
transform 1 0 3868 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2210
timestamp 1677677812
transform 1 0 3844 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2211
timestamp 1677677812
transform 1 0 3860 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1847
timestamp 1677677812
transform 1 0 3852 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1890
timestamp 1677677812
transform 1 0 3868 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1848
timestamp 1677677812
transform 1 0 3892 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1808
timestamp 1677677812
transform 1 0 3908 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2212
timestamp 1677677812
transform 1 0 3916 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2116
timestamp 1677677812
transform 1 0 4044 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2213
timestamp 1677677812
transform 1 0 3996 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1849
timestamp 1677677812
transform 1 0 3972 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1850
timestamp 1677677812
transform 1 0 3996 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1891
timestamp 1677677812
transform 1 0 3988 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1871
timestamp 1677677812
transform 1 0 4092 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1790
timestamp 1677677812
transform 1 0 4132 0 1 3735
box -3 -3 3 3
use M3_M2  M3_M2_1791
timestamp 1677677812
transform 1 0 4148 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2117
timestamp 1677677812
transform 1 0 4172 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2118
timestamp 1677677812
transform 1 0 4244 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2214
timestamp 1677677812
transform 1 0 4276 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1745
timestamp 1677677812
transform 1 0 4348 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1792
timestamp 1677677812
transform 1 0 4348 0 1 3735
box -3 -3 3 3
use M2_M1  M2_M1_2215
timestamp 1677677812
transform 1 0 4372 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1718
timestamp 1677677812
transform 1 0 4420 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2119
timestamp 1677677812
transform 1 0 4444 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2120
timestamp 1677677812
transform 1 0 4452 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1809
timestamp 1677677812
transform 1 0 4444 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2121
timestamp 1677677812
transform 1 0 4476 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1810
timestamp 1677677812
transform 1 0 4476 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1719
timestamp 1677677812
transform 1 0 4500 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2122
timestamp 1677677812
transform 1 0 4500 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2216
timestamp 1677677812
transform 1 0 4484 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2217
timestamp 1677677812
transform 1 0 4492 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2218
timestamp 1677677812
transform 1 0 4508 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1851
timestamp 1677677812
transform 1 0 4484 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1852
timestamp 1677677812
transform 1 0 4508 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1872
timestamp 1677677812
transform 1 0 4516 0 1 3705
box -3 -3 3 3
use M2_M1  M2_M1_2123
timestamp 1677677812
transform 1 0 4532 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1720
timestamp 1677677812
transform 1 0 4580 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1721
timestamp 1677677812
transform 1 0 4652 0 1 3765
box -3 -3 3 3
use M3_M2  M3_M2_1746
timestamp 1677677812
transform 1 0 4564 0 1 3755
box -3 -3 3 3
use M3_M2  M3_M2_1771
timestamp 1677677812
transform 1 0 4548 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2124
timestamp 1677677812
transform 1 0 4540 0 1 3735
box -2 -2 2 2
use M3_M2  M3_M2_1772
timestamp 1677677812
transform 1 0 4628 0 1 3745
box -3 -3 3 3
use M3_M2  M3_M2_1773
timestamp 1677677812
transform 1 0 4644 0 1 3745
box -3 -3 3 3
use M2_M1  M2_M1_2125
timestamp 1677677812
transform 1 0 4580 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2126
timestamp 1677677812
transform 1 0 4596 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2219
timestamp 1677677812
transform 1 0 4548 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2220
timestamp 1677677812
transform 1 0 4564 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2221
timestamp 1677677812
transform 1 0 4580 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2222
timestamp 1677677812
transform 1 0 4620 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1853
timestamp 1677677812
transform 1 0 4540 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1892
timestamp 1677677812
transform 1 0 4548 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1811
timestamp 1677677812
transform 1 0 4668 0 1 3725
box -3 -3 3 3
use M3_M2  M3_M2_1722
timestamp 1677677812
transform 1 0 4788 0 1 3765
box -3 -3 3 3
use M2_M1  M2_M1_2127
timestamp 1677677812
transform 1 0 4692 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2128
timestamp 1677677812
transform 1 0 4780 0 1 3735
box -2 -2 2 2
use M2_M1  M2_M1_2223
timestamp 1677677812
transform 1 0 4676 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2224
timestamp 1677677812
transform 1 0 4716 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1854
timestamp 1677677812
transform 1 0 4668 0 1 3715
box -3 -3 3 3
use M3_M2  M3_M2_1873
timestamp 1677677812
transform 1 0 4620 0 1 3705
box -3 -3 3 3
use M3_M2  M3_M2_1893
timestamp 1677677812
transform 1 0 4604 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1894
timestamp 1677677812
transform 1 0 4628 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1895
timestamp 1677677812
transform 1 0 4644 0 1 3685
box -3 -3 3 3
use M3_M2  M3_M2_1812
timestamp 1677677812
transform 1 0 4740 0 1 3725
box -3 -3 3 3
use M2_M1  M2_M1_2225
timestamp 1677677812
transform 1 0 4772 0 1 3725
box -2 -2 2 2
use M2_M1  M2_M1_2226
timestamp 1677677812
transform 1 0 4788 0 1 3725
box -2 -2 2 2
use M3_M2  M3_M2_1855
timestamp 1677677812
transform 1 0 4716 0 1 3715
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_20
timestamp 1677677812
transform 1 0 24 0 1 3670
box -10 -3 10 3
use FILL  FILL_1706
timestamp 1677677812
transform 1 0 72 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1710
timestamp 1677677812
transform 1 0 80 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_149
timestamp 1677677812
transform 1 0 88 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1711
timestamp 1677677812
transform 1 0 104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1712
timestamp 1677677812
transform 1 0 112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1713
timestamp 1677677812
transform 1 0 120 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_150
timestamp 1677677812
transform -1 0 144 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1714
timestamp 1677677812
transform 1 0 144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1715
timestamp 1677677812
transform 1 0 152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1716
timestamp 1677677812
transform 1 0 160 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_85
timestamp 1677677812
transform -1 0 208 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1717
timestamp 1677677812
transform 1 0 208 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1718
timestamp 1677677812
transform 1 0 216 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1719
timestamp 1677677812
transform 1 0 224 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1720
timestamp 1677677812
transform 1 0 232 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_85
timestamp 1677677812
transform 1 0 240 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1737
timestamp 1677677812
transform 1 0 280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1738
timestamp 1677677812
transform 1 0 288 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_134
timestamp 1677677812
transform 1 0 296 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1739
timestamp 1677677812
transform 1 0 392 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_153
timestamp 1677677812
transform -1 0 416 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1740
timestamp 1677677812
transform 1 0 416 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1741
timestamp 1677677812
transform 1 0 424 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1742
timestamp 1677677812
transform 1 0 432 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_88
timestamp 1677677812
transform 1 0 440 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1743
timestamp 1677677812
transform 1 0 480 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1744
timestamp 1677677812
transform 1 0 488 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1745
timestamp 1677677812
transform 1 0 496 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_135
timestamp 1677677812
transform 1 0 504 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1746
timestamp 1677677812
transform 1 0 600 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1747
timestamp 1677677812
transform 1 0 608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1749
timestamp 1677677812
transform 1 0 616 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1751
timestamp 1677677812
transform 1 0 624 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_90
timestamp 1677677812
transform 1 0 632 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1755
timestamp 1677677812
transform 1 0 672 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1756
timestamp 1677677812
transform 1 0 680 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1757
timestamp 1677677812
transform 1 0 688 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1759
timestamp 1677677812
transform 1 0 696 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1761
timestamp 1677677812
transform 1 0 704 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1763
timestamp 1677677812
transform 1 0 712 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_154
timestamp 1677677812
transform 1 0 720 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_155
timestamp 1677677812
transform 1 0 736 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1772
timestamp 1677677812
transform 1 0 752 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1773
timestamp 1677677812
transform 1 0 760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1774
timestamp 1677677812
transform 1 0 768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1775
timestamp 1677677812
transform 1 0 776 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_137
timestamp 1677677812
transform 1 0 784 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_156
timestamp 1677677812
transform -1 0 896 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1776
timestamp 1677677812
transform 1 0 896 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1777
timestamp 1677677812
transform 1 0 904 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1778
timestamp 1677677812
transform 1 0 912 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1780
timestamp 1677677812
transform 1 0 920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1782
timestamp 1677677812
transform 1 0 928 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1784
timestamp 1677677812
transform 1 0 936 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1896
timestamp 1677677812
transform 1 0 964 0 1 3675
box -3 -3 3 3
use NOR2X1  NOR2X1_20
timestamp 1677677812
transform 1 0 944 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1791
timestamp 1677677812
transform 1 0 968 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_41
timestamp 1677677812
transform 1 0 976 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1792
timestamp 1677677812
transform 1 0 1008 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1794
timestamp 1677677812
transform 1 0 1016 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1795
timestamp 1677677812
transform 1 0 1024 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1796
timestamp 1677677812
transform 1 0 1032 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1797
timestamp 1677677812
transform 1 0 1040 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1799
timestamp 1677677812
transform 1 0 1048 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_22
timestamp 1677677812
transform 1 0 1056 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1807
timestamp 1677677812
transform 1 0 1080 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1808
timestamp 1677677812
transform 1 0 1088 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1809
timestamp 1677677812
transform 1 0 1096 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_43
timestamp 1677677812
transform -1 0 1136 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1810
timestamp 1677677812
transform 1 0 1136 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1812
timestamp 1677677812
transform 1 0 1144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1814
timestamp 1677677812
transform 1 0 1152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1816
timestamp 1677677812
transform 1 0 1160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1822
timestamp 1677677812
transform 1 0 1168 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_92
timestamp 1677677812
transform -1 0 1216 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1823
timestamp 1677677812
transform 1 0 1216 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1825
timestamp 1677677812
transform 1 0 1224 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1827
timestamp 1677677812
transform 1 0 1232 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_158
timestamp 1677677812
transform 1 0 1240 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1830
timestamp 1677677812
transform 1 0 1256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1831
timestamp 1677677812
transform 1 0 1264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1832
timestamp 1677677812
transform 1 0 1272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1833
timestamp 1677677812
transform 1 0 1280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1838
timestamp 1677677812
transform 1 0 1288 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_45
timestamp 1677677812
transform -1 0 1328 0 -1 3770
box -8 -3 34 105
use INVX2  INVX2_159
timestamp 1677677812
transform -1 0 1344 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1839
timestamp 1677677812
transform 1 0 1344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1840
timestamp 1677677812
transform 1 0 1352 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1841
timestamp 1677677812
transform 1 0 1360 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_46
timestamp 1677677812
transform -1 0 1400 0 -1 3770
box -8 -3 34 105
use FILL  FILL_1842
timestamp 1677677812
transform 1 0 1400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1843
timestamp 1677677812
transform 1 0 1408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1845
timestamp 1677677812
transform 1 0 1416 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1847
timestamp 1677677812
transform 1 0 1424 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_139
timestamp 1677677812
transform 1 0 1432 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1855
timestamp 1677677812
transform 1 0 1528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1856
timestamp 1677677812
transform 1 0 1536 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_161
timestamp 1677677812
transform 1 0 1544 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1860
timestamp 1677677812
transform 1 0 1560 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1862
timestamp 1677677812
transform 1 0 1568 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1864
timestamp 1677677812
transform 1 0 1576 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1866
timestamp 1677677812
transform 1 0 1584 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1868
timestamp 1677677812
transform 1 0 1592 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1874
timestamp 1677677812
transform 1 0 1600 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_87
timestamp 1677677812
transform -1 0 1648 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1875
timestamp 1677677812
transform 1 0 1648 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1877
timestamp 1677677812
transform 1 0 1656 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1879
timestamp 1677677812
transform 1 0 1664 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1889
timestamp 1677677812
transform 1 0 1672 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1890
timestamp 1677677812
transform 1 0 1680 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_140
timestamp 1677677812
transform 1 0 1688 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_164
timestamp 1677677812
transform -1 0 1800 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1891
timestamp 1677677812
transform 1 0 1800 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1893
timestamp 1677677812
transform 1 0 1808 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1908
timestamp 1677677812
transform 1 0 1816 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1897
timestamp 1677677812
transform 1 0 1836 0 1 3675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_143
timestamp 1677677812
transform -1 0 1920 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1909
timestamp 1677677812
transform 1 0 1920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1910
timestamp 1677677812
transform 1 0 1928 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_165
timestamp 1677677812
transform -1 0 1952 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1911
timestamp 1677677812
transform 1 0 1952 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1912
timestamp 1677677812
transform 1 0 1960 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1913
timestamp 1677677812
transform 1 0 1968 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1914
timestamp 1677677812
transform 1 0 1976 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_94
timestamp 1677677812
transform -1 0 2024 0 -1 3770
box -8 -3 46 105
use INVX2  INVX2_166
timestamp 1677677812
transform 1 0 2024 0 -1 3770
box -9 -3 26 105
use M3_M2  M3_M2_1898
timestamp 1677677812
transform 1 0 2068 0 1 3675
box -3 -3 3 3
use M3_M2  M3_M2_1899
timestamp 1677677812
transform 1 0 2084 0 1 3675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_144
timestamp 1677677812
transform 1 0 2040 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_167
timestamp 1677677812
transform -1 0 2152 0 -1 3770
box -9 -3 26 105
use AOI22X1  AOI22X1_95
timestamp 1677677812
transform 1 0 2152 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1915
timestamp 1677677812
transform 1 0 2192 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1917
timestamp 1677677812
transform 1 0 2200 0 -1 3770
box -8 -3 16 105
use M3_M2  M3_M2_1900
timestamp 1677677812
transform 1 0 2220 0 1 3675
box -3 -3 3 3
use FILL  FILL_1919
timestamp 1677677812
transform 1 0 2208 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1921
timestamp 1677677812
transform 1 0 2216 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1923
timestamp 1677677812
transform 1 0 2224 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_168
timestamp 1677677812
transform 1 0 2232 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1927
timestamp 1677677812
transform 1 0 2248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1929
timestamp 1677677812
transform 1 0 2256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1931
timestamp 1677677812
transform 1 0 2264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1933
timestamp 1677677812
transform 1 0 2272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1935
timestamp 1677677812
transform 1 0 2280 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_89
timestamp 1677677812
transform 1 0 2288 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1937
timestamp 1677677812
transform 1 0 2328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1939
timestamp 1677677812
transform 1 0 2336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1941
timestamp 1677677812
transform 1 0 2344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1944
timestamp 1677677812
transform 1 0 2352 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1945
timestamp 1677677812
transform 1 0 2360 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_146
timestamp 1677677812
transform -1 0 2464 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1946
timestamp 1677677812
transform 1 0 2464 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1947
timestamp 1677677812
transform 1 0 2472 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1948
timestamp 1677677812
transform 1 0 2480 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1949
timestamp 1677677812
transform 1 0 2488 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1950
timestamp 1677677812
transform 1 0 2496 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1952
timestamp 1677677812
transform 1 0 2504 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1954
timestamp 1677677812
transform 1 0 2512 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1958
timestamp 1677677812
transform 1 0 2520 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1959
timestamp 1677677812
transform 1 0 2528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1960
timestamp 1677677812
transform 1 0 2536 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1961
timestamp 1677677812
transform 1 0 2544 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_98
timestamp 1677677812
transform 1 0 2552 0 -1 3770
box -8 -3 46 105
use FILL  FILL_1962
timestamp 1677677812
transform 1 0 2592 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1964
timestamp 1677677812
transform 1 0 2600 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_171
timestamp 1677677812
transform 1 0 2608 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1971
timestamp 1677677812
transform 1 0 2624 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1972
timestamp 1677677812
transform 1 0 2632 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1973
timestamp 1677677812
transform 1 0 2640 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_148
timestamp 1677677812
transform 1 0 2648 0 -1 3770
box -8 -3 104 105
use FILL  FILL_1974
timestamp 1677677812
transform 1 0 2744 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1975
timestamp 1677677812
transform 1 0 2752 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1976
timestamp 1677677812
transform 1 0 2760 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1977
timestamp 1677677812
transform 1 0 2768 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1978
timestamp 1677677812
transform 1 0 2776 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1980
timestamp 1677677812
transform 1 0 2784 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_24
timestamp 1677677812
transform 1 0 2792 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1982
timestamp 1677677812
transform 1 0 2816 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1984
timestamp 1677677812
transform 1 0 2824 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1986
timestamp 1677677812
transform 1 0 2832 0 -1 3770
box -8 -3 16 105
use NOR2X1  NOR2X1_25
timestamp 1677677812
transform 1 0 2840 0 -1 3770
box -8 -3 32 105
use FILL  FILL_1987
timestamp 1677677812
transform 1 0 2864 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1989
timestamp 1677677812
transform 1 0 2872 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1992
timestamp 1677677812
transform 1 0 2880 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_172
timestamp 1677677812
transform 1 0 2888 0 -1 3770
box -9 -3 26 105
use FILL  FILL_1993
timestamp 1677677812
transform 1 0 2904 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1994
timestamp 1677677812
transform 1 0 2912 0 -1 3770
box -8 -3 16 105
use FILL  FILL_1995
timestamp 1677677812
transform 1 0 2920 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_173
timestamp 1677677812
transform 1 0 2928 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2012
timestamp 1677677812
transform 1 0 2944 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2013
timestamp 1677677812
transform 1 0 2952 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2014
timestamp 1677677812
transform 1 0 2960 0 -1 3770
box -8 -3 16 105
use OAI21X1  OAI21X1_51
timestamp 1677677812
transform -1 0 3000 0 -1 3770
box -8 -3 34 105
use FILL  FILL_2015
timestamp 1677677812
transform 1 0 3000 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2016
timestamp 1677677812
transform 1 0 3008 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2017
timestamp 1677677812
transform 1 0 3016 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2018
timestamp 1677677812
transform 1 0 3024 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2019
timestamp 1677677812
transform 1 0 3032 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_174
timestamp 1677677812
transform -1 0 3056 0 -1 3770
box -9 -3 26 105
use INVX2  INVX2_175
timestamp 1677677812
transform -1 0 3072 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2020
timestamp 1677677812
transform 1 0 3072 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2021
timestamp 1677677812
transform 1 0 3080 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2022
timestamp 1677677812
transform 1 0 3088 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2023
timestamp 1677677812
transform 1 0 3096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2024
timestamp 1677677812
transform 1 0 3104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2025
timestamp 1677677812
transform 1 0 3112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2026
timestamp 1677677812
transform 1 0 3120 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2027
timestamp 1677677812
transform 1 0 3128 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2028
timestamp 1677677812
transform 1 0 3136 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2029
timestamp 1677677812
transform 1 0 3144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2030
timestamp 1677677812
transform 1 0 3152 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_150
timestamp 1677677812
transform 1 0 3160 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2031
timestamp 1677677812
transform 1 0 3256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2033
timestamp 1677677812
transform 1 0 3264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2035
timestamp 1677677812
transform 1 0 3272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2038
timestamp 1677677812
transform 1 0 3280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2039
timestamp 1677677812
transform 1 0 3288 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2040
timestamp 1677677812
transform 1 0 3296 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2041
timestamp 1677677812
transform 1 0 3304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2043
timestamp 1677677812
transform 1 0 3312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2045
timestamp 1677677812
transform 1 0 3320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2047
timestamp 1677677812
transform 1 0 3328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2052
timestamp 1677677812
transform 1 0 3336 0 -1 3770
box -8 -3 16 105
use NAND3X1  NAND3X1_9
timestamp 1677677812
transform -1 0 3376 0 -1 3770
box -8 -3 40 105
use FILL  FILL_2053
timestamp 1677677812
transform 1 0 3376 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2055
timestamp 1677677812
transform 1 0 3384 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2057
timestamp 1677677812
transform 1 0 3392 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2059
timestamp 1677677812
transform 1 0 3400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2061
timestamp 1677677812
transform 1 0 3408 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2063
timestamp 1677677812
transform 1 0 3416 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_151
timestamp 1677677812
transform 1 0 3424 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2072
timestamp 1677677812
transform 1 0 3520 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2074
timestamp 1677677812
transform 1 0 3528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2076
timestamp 1677677812
transform 1 0 3536 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2078
timestamp 1677677812
transform 1 0 3544 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2082
timestamp 1677677812
transform 1 0 3552 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2083
timestamp 1677677812
transform 1 0 3560 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_179
timestamp 1677677812
transform -1 0 3584 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2084
timestamp 1677677812
transform 1 0 3584 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2086
timestamp 1677677812
transform 1 0 3592 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2088
timestamp 1677677812
transform 1 0 3600 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2100
timestamp 1677677812
transform 1 0 3608 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2101
timestamp 1677677812
transform 1 0 3616 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2102
timestamp 1677677812
transform 1 0 3624 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_152
timestamp 1677677812
transform -1 0 3728 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2103
timestamp 1677677812
transform 1 0 3728 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2105
timestamp 1677677812
transform 1 0 3736 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2107
timestamp 1677677812
transform 1 0 3744 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2112
timestamp 1677677812
transform 1 0 3752 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2113
timestamp 1677677812
transform 1 0 3760 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_180
timestamp 1677677812
transform 1 0 3768 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2114
timestamp 1677677812
transform 1 0 3784 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_181
timestamp 1677677812
transform 1 0 3792 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2115
timestamp 1677677812
transform 1 0 3808 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2116
timestamp 1677677812
transform 1 0 3816 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2117
timestamp 1677677812
transform 1 0 3824 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_93
timestamp 1677677812
transform -1 0 3872 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2118
timestamp 1677677812
transform 1 0 3872 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2121
timestamp 1677677812
transform 1 0 3880 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2122
timestamp 1677677812
transform 1 0 3888 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2123
timestamp 1677677812
transform 1 0 3896 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2124
timestamp 1677677812
transform 1 0 3904 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2125
timestamp 1677677812
transform 1 0 3912 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2126
timestamp 1677677812
transform 1 0 3920 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2127
timestamp 1677677812
transform 1 0 3928 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2135
timestamp 1677677812
transform 1 0 3936 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2136
timestamp 1677677812
transform 1 0 3944 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2137
timestamp 1677677812
transform 1 0 3952 0 -1 3770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_154
timestamp 1677677812
transform -1 0 4056 0 -1 3770
box -8 -3 104 105
use FILL  FILL_2138
timestamp 1677677812
transform 1 0 4056 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2139
timestamp 1677677812
transform 1 0 4064 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2140
timestamp 1677677812
transform 1 0 4072 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2141
timestamp 1677677812
transform 1 0 4080 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2143
timestamp 1677677812
transform 1 0 4088 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2145
timestamp 1677677812
transform 1 0 4096 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2146
timestamp 1677677812
transform 1 0 4104 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2147
timestamp 1677677812
transform 1 0 4112 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2149
timestamp 1677677812
transform 1 0 4120 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2151
timestamp 1677677812
transform 1 0 4128 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2153
timestamp 1677677812
transform 1 0 4136 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2155
timestamp 1677677812
transform 1 0 4144 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2156
timestamp 1677677812
transform 1 0 4152 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2157
timestamp 1677677812
transform 1 0 4160 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2158
timestamp 1677677812
transform 1 0 4168 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2159
timestamp 1677677812
transform 1 0 4176 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2160
timestamp 1677677812
transform 1 0 4184 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2162
timestamp 1677677812
transform 1 0 4192 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2164
timestamp 1677677812
transform 1 0 4200 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2166
timestamp 1677677812
transform 1 0 4208 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2171
timestamp 1677677812
transform 1 0 4216 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_184
timestamp 1677677812
transform -1 0 4240 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2172
timestamp 1677677812
transform 1 0 4240 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2175
timestamp 1677677812
transform 1 0 4248 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2176
timestamp 1677677812
transform 1 0 4256 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2177
timestamp 1677677812
transform 1 0 4264 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2178
timestamp 1677677812
transform 1 0 4272 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2179
timestamp 1677677812
transform 1 0 4280 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2180
timestamp 1677677812
transform 1 0 4288 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2181
timestamp 1677677812
transform 1 0 4296 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2183
timestamp 1677677812
transform 1 0 4304 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2185
timestamp 1677677812
transform 1 0 4312 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2188
timestamp 1677677812
transform 1 0 4320 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2189
timestamp 1677677812
transform 1 0 4328 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2190
timestamp 1677677812
transform 1 0 4336 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2191
timestamp 1677677812
transform 1 0 4344 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2192
timestamp 1677677812
transform 1 0 4352 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2193
timestamp 1677677812
transform 1 0 4360 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2195
timestamp 1677677812
transform 1 0 4368 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2197
timestamp 1677677812
transform 1 0 4376 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2198
timestamp 1677677812
transform 1 0 4384 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2199
timestamp 1677677812
transform 1 0 4392 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2200
timestamp 1677677812
transform 1 0 4400 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2201
timestamp 1677677812
transform 1 0 4408 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_185
timestamp 1677677812
transform -1 0 4432 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2202
timestamp 1677677812
transform 1 0 4432 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2203
timestamp 1677677812
transform 1 0 4440 0 -1 3770
box -8 -3 16 105
use INVX2  INVX2_186
timestamp 1677677812
transform 1 0 4448 0 -1 3770
box -9 -3 26 105
use FILL  FILL_2204
timestamp 1677677812
transform 1 0 4464 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2205
timestamp 1677677812
transform 1 0 4472 0 -1 3770
box -8 -3 16 105
use OAI22X1  OAI22X1_98
timestamp 1677677812
transform 1 0 4480 0 -1 3770
box -8 -3 46 105
use FILL  FILL_2216
timestamp 1677677812
transform 1 0 4520 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2217
timestamp 1677677812
transform 1 0 4528 0 -1 3770
box -8 -3 16 105
use FILL  FILL_2218
timestamp 1677677812
transform 1 0 4536 0 -1 3770
box -8 -3 16 105
use AOI22X1  AOI22X1_102
timestamp 1677677812
transform -1 0 4584 0 -1 3770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_158
timestamp 1677677812
transform 1 0 4584 0 -1 3770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_159
timestamp 1677677812
transform 1 0 4680 0 -1 3770
box -8 -3 104 105
use INVX2  INVX2_187
timestamp 1677677812
transform 1 0 4776 0 -1 3770
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_21
timestamp 1677677812
transform 1 0 4843 0 1 3670
box -10 -3 10 3
use M2_M1  M2_M1_2247
timestamp 1677677812
transform 1 0 108 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2355
timestamp 1677677812
transform 1 0 84 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2248
timestamp 1677677812
transform 1 0 180 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1939
timestamp 1677677812
transform 1 0 236 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1983
timestamp 1677677812
transform 1 0 308 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2006
timestamp 1677677812
transform 1 0 428 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1905
timestamp 1677677812
transform 1 0 484 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2356
timestamp 1677677812
transform 1 0 500 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2249
timestamp 1677677812
transform 1 0 556 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1906
timestamp 1677677812
transform 1 0 612 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1907
timestamp 1677677812
transform 1 0 636 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1984
timestamp 1677677812
transform 1 0 716 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2250
timestamp 1677677812
transform 1 0 740 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2251
timestamp 1677677812
transform 1 0 796 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2357
timestamp 1677677812
transform 1 0 716 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1985
timestamp 1677677812
transform 1 0 812 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2252
timestamp 1677677812
transform 1 0 836 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2253
timestamp 1677677812
transform 1 0 892 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2358
timestamp 1677677812
transform 1 0 812 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1950
timestamp 1677677812
transform 1 0 924 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1951
timestamp 1677677812
transform 1 0 948 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2254
timestamp 1677677812
transform 1 0 916 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2255
timestamp 1677677812
transform 1 0 932 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2029
timestamp 1677677812
transform 1 0 948 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1940
timestamp 1677677812
transform 1 0 964 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2256
timestamp 1677677812
transform 1 0 964 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1941
timestamp 1677677812
transform 1 0 980 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1986
timestamp 1677677812
transform 1 0 980 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2359
timestamp 1677677812
transform 1 0 972 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2050
timestamp 1677677812
transform 1 0 972 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2030
timestamp 1677677812
transform 1 0 988 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1921
timestamp 1677677812
transform 1 0 1020 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1942
timestamp 1677677812
transform 1 0 1012 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2257
timestamp 1677677812
transform 1 0 1004 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1952
timestamp 1677677812
transform 1 0 1020 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2258
timestamp 1677677812
transform 1 0 1020 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1953
timestamp 1677677812
transform 1 0 1036 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2360
timestamp 1677677812
transform 1 0 1036 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1943
timestamp 1677677812
transform 1 0 1092 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1954
timestamp 1677677812
transform 1 0 1068 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1955
timestamp 1677677812
transform 1 0 1084 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2259
timestamp 1677677812
transform 1 0 1068 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2260
timestamp 1677677812
transform 1 0 1092 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2361
timestamp 1677677812
transform 1 0 1060 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2362
timestamp 1677677812
transform 1 0 1076 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2363
timestamp 1677677812
transform 1 0 1084 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2031
timestamp 1677677812
transform 1 0 1076 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2007
timestamp 1677677812
transform 1 0 1092 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1987
timestamp 1677677812
transform 1 0 1108 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2364
timestamp 1677677812
transform 1 0 1100 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2261
timestamp 1677677812
transform 1 0 1132 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2262
timestamp 1677677812
transform 1 0 1140 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1988
timestamp 1677677812
transform 1 0 1148 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1908
timestamp 1677677812
transform 1 0 1164 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1909
timestamp 1677677812
transform 1 0 1204 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1922
timestamp 1677677812
transform 1 0 1180 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1923
timestamp 1677677812
transform 1 0 1196 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1956
timestamp 1677677812
transform 1 0 1172 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1957
timestamp 1677677812
transform 1 0 1204 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2263
timestamp 1677677812
transform 1 0 1164 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2264
timestamp 1677677812
transform 1 0 1180 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2265
timestamp 1677677812
transform 1 0 1196 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2365
timestamp 1677677812
transform 1 0 1164 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2366
timestamp 1677677812
transform 1 0 1172 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2367
timestamp 1677677812
transform 1 0 1196 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2032
timestamp 1677677812
transform 1 0 1196 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2238
timestamp 1677677812
transform 1 0 1236 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2368
timestamp 1677677812
transform 1 0 1236 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2266
timestamp 1677677812
transform 1 0 1276 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2267
timestamp 1677677812
transform 1 0 1284 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2369
timestamp 1677677812
transform 1 0 1268 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2033
timestamp 1677677812
transform 1 0 1268 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2370
timestamp 1677677812
transform 1 0 1308 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1910
timestamp 1677677812
transform 1 0 1356 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2239
timestamp 1677677812
transform 1 0 1348 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_2034
timestamp 1677677812
transform 1 0 1348 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1924
timestamp 1677677812
transform 1 0 1460 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2268
timestamp 1677677812
transform 1 0 1380 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2269
timestamp 1677677812
transform 1 0 1428 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2371
timestamp 1677677812
transform 1 0 1460 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2372
timestamp 1677677812
transform 1 0 1484 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2008
timestamp 1677677812
transform 1 0 1492 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2270
timestamp 1677677812
transform 1 0 1524 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2271
timestamp 1677677812
transform 1 0 1540 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2373
timestamp 1677677812
transform 1 0 1516 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2009
timestamp 1677677812
transform 1 0 1524 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2374
timestamp 1677677812
transform 1 0 1532 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2272
timestamp 1677677812
transform 1 0 1556 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2273
timestamp 1677677812
transform 1 0 1580 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1911
timestamp 1677677812
transform 1 0 1604 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1901
timestamp 1677677812
transform 1 0 1620 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2274
timestamp 1677677812
transform 1 0 1612 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2375
timestamp 1677677812
transform 1 0 1604 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1925
timestamp 1677677812
transform 1 0 1636 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2275
timestamp 1677677812
transform 1 0 1660 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2376
timestamp 1677677812
transform 1 0 1620 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2377
timestamp 1677677812
transform 1 0 1636 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1926
timestamp 1677677812
transform 1 0 1724 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2276
timestamp 1677677812
transform 1 0 1748 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2277
timestamp 1677677812
transform 1 0 1772 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2051
timestamp 1677677812
transform 1 0 1764 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1927
timestamp 1677677812
transform 1 0 1796 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1902
timestamp 1677677812
transform 1 0 1812 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1958
timestamp 1677677812
transform 1 0 1804 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2052
timestamp 1677677812
transform 1 0 1804 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2378
timestamp 1677677812
transform 1 0 1820 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1928
timestamp 1677677812
transform 1 0 1844 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2278
timestamp 1677677812
transform 1 0 1844 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1903
timestamp 1677677812
transform 1 0 1892 0 1 3665
box -3 -3 3 3
use M3_M2  M3_M2_1929
timestamp 1677677812
transform 1 0 1876 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1959
timestamp 1677677812
transform 1 0 1876 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2279
timestamp 1677677812
transform 1 0 1868 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2280
timestamp 1677677812
transform 1 0 1884 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2281
timestamp 1677677812
transform 1 0 1900 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2379
timestamp 1677677812
transform 1 0 1868 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2380
timestamp 1677677812
transform 1 0 1876 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2381
timestamp 1677677812
transform 1 0 1892 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1930
timestamp 1677677812
transform 1 0 1980 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1944
timestamp 1677677812
transform 1 0 1988 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2282
timestamp 1677677812
transform 1 0 1964 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2283
timestamp 1677677812
transform 1 0 1980 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2284
timestamp 1677677812
transform 1 0 1988 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2382
timestamp 1677677812
transform 1 0 1948 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2383
timestamp 1677677812
transform 1 0 1956 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2384
timestamp 1677677812
transform 1 0 1972 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2053
timestamp 1677677812
transform 1 0 1956 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2385
timestamp 1677677812
transform 1 0 1988 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2054
timestamp 1677677812
transform 1 0 1988 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2386
timestamp 1677677812
transform 1 0 2012 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1912
timestamp 1677677812
transform 1 0 2028 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1931
timestamp 1677677812
transform 1 0 2060 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2285
timestamp 1677677812
transform 1 0 2028 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2286
timestamp 1677677812
transform 1 0 2044 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2287
timestamp 1677677812
transform 1 0 2060 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2387
timestamp 1677677812
transform 1 0 2068 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1913
timestamp 1677677812
transform 1 0 2076 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1932
timestamp 1677677812
transform 1 0 2076 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1914
timestamp 1677677812
transform 1 0 2108 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1945
timestamp 1677677812
transform 1 0 2116 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2288
timestamp 1677677812
transform 1 0 2108 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2289
timestamp 1677677812
transform 1 0 2124 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2388
timestamp 1677677812
transform 1 0 2116 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2290
timestamp 1677677812
transform 1 0 2140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2389
timestamp 1677677812
transform 1 0 2148 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2055
timestamp 1677677812
transform 1 0 2148 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1904
timestamp 1677677812
transform 1 0 2164 0 1 3665
box -3 -3 3 3
use M2_M1  M2_M1_2390
timestamp 1677677812
transform 1 0 2164 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1933
timestamp 1677677812
transform 1 0 2188 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2391
timestamp 1677677812
transform 1 0 2188 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2291
timestamp 1677677812
transform 1 0 2244 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2392
timestamp 1677677812
transform 1 0 2220 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2010
timestamp 1677677812
transform 1 0 2244 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2011
timestamp 1677677812
transform 1 0 2268 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2012
timestamp 1677677812
transform 1 0 2292 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1915
timestamp 1677677812
transform 1 0 2324 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1989
timestamp 1677677812
transform 1 0 2316 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1934
timestamp 1677677812
transform 1 0 2340 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2292
timestamp 1677677812
transform 1 0 2340 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1916
timestamp 1677677812
transform 1 0 2380 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2293
timestamp 1677677812
transform 1 0 2364 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2294
timestamp 1677677812
transform 1 0 2380 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2393
timestamp 1677677812
transform 1 0 2348 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2394
timestamp 1677677812
transform 1 0 2372 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2013
timestamp 1677677812
transform 1 0 2388 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1935
timestamp 1677677812
transform 1 0 2420 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1960
timestamp 1677677812
transform 1 0 2428 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1961
timestamp 1677677812
transform 1 0 2468 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1962
timestamp 1677677812
transform 1 0 2492 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1963
timestamp 1677677812
transform 1 0 2532 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1990
timestamp 1677677812
transform 1 0 2420 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2295
timestamp 1677677812
transform 1 0 2428 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2296
timestamp 1677677812
transform 1 0 2436 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1991
timestamp 1677677812
transform 1 0 2452 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2297
timestamp 1677677812
transform 1 0 2468 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1992
timestamp 1677677812
transform 1 0 2476 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1993
timestamp 1677677812
transform 1 0 2516 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2298
timestamp 1677677812
transform 1 0 2532 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2395
timestamp 1677677812
transform 1 0 2420 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2014
timestamp 1677677812
transform 1 0 2436 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2015
timestamp 1677677812
transform 1 0 2476 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2396
timestamp 1677677812
transform 1 0 2516 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2397
timestamp 1677677812
transform 1 0 2532 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2056
timestamp 1677677812
transform 1 0 2436 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2057
timestamp 1677677812
transform 1 0 2484 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2058
timestamp 1677677812
transform 1 0 2500 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2016
timestamp 1677677812
transform 1 0 2540 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2398
timestamp 1677677812
transform 1 0 2556 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2240
timestamp 1677677812
transform 1 0 2572 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1964
timestamp 1677677812
transform 1 0 2588 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1965
timestamp 1677677812
transform 1 0 2620 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1994
timestamp 1677677812
transform 1 0 2588 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2299
timestamp 1677677812
transform 1 0 2612 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1995
timestamp 1677677812
transform 1 0 2660 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2300
timestamp 1677677812
transform 1 0 2668 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2399
timestamp 1677677812
transform 1 0 2588 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2059
timestamp 1677677812
transform 1 0 2588 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_2060
timestamp 1677677812
transform 1 0 2620 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2301
timestamp 1677677812
transform 1 0 2684 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2302
timestamp 1677677812
transform 1 0 2740 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1996
timestamp 1677677812
transform 1 0 2764 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2400
timestamp 1677677812
transform 1 0 2764 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1936
timestamp 1677677812
transform 1 0 2788 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2303
timestamp 1677677812
transform 1 0 2788 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2401
timestamp 1677677812
transform 1 0 2780 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2402
timestamp 1677677812
transform 1 0 2812 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2241
timestamp 1677677812
transform 1 0 2828 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1997
timestamp 1677677812
transform 1 0 2828 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2017
timestamp 1677677812
transform 1 0 2828 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2450
timestamp 1677677812
transform 1 0 2828 0 1 3595
box -2 -2 2 2
use M2_M1  M2_M1_2242
timestamp 1677677812
transform 1 0 2868 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2304
timestamp 1677677812
transform 1 0 2860 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2035
timestamp 1677677812
transform 1 0 2868 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2305
timestamp 1677677812
transform 1 0 2884 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1998
timestamp 1677677812
transform 1 0 2916 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2306
timestamp 1677677812
transform 1 0 2932 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2403
timestamp 1677677812
transform 1 0 2892 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2404
timestamp 1677677812
transform 1 0 2908 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2405
timestamp 1677677812
transform 1 0 2916 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2307
timestamp 1677677812
transform 1 0 2948 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1999
timestamp 1677677812
transform 1 0 2964 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_1966
timestamp 1677677812
transform 1 0 2980 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2406
timestamp 1677677812
transform 1 0 2980 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1967
timestamp 1677677812
transform 1 0 3068 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2000
timestamp 1677677812
transform 1 0 2996 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2308
timestamp 1677677812
transform 1 0 3044 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2309
timestamp 1677677812
transform 1 0 3076 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2310
timestamp 1677677812
transform 1 0 3084 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2407
timestamp 1677677812
transform 1 0 2996 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2036
timestamp 1677677812
transform 1 0 3044 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2408
timestamp 1677677812
transform 1 0 3084 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2311
timestamp 1677677812
transform 1 0 3100 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1968
timestamp 1677677812
transform 1 0 3124 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2312
timestamp 1677677812
transform 1 0 3124 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2313
timestamp 1677677812
transform 1 0 3140 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2314
timestamp 1677677812
transform 1 0 3156 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2409
timestamp 1677677812
transform 1 0 3132 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2410
timestamp 1677677812
transform 1 0 3148 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2037
timestamp 1677677812
transform 1 0 3132 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2411
timestamp 1677677812
transform 1 0 3172 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2412
timestamp 1677677812
transform 1 0 3196 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2038
timestamp 1677677812
transform 1 0 3196 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2413
timestamp 1677677812
transform 1 0 3252 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2236
timestamp 1677677812
transform 1 0 3284 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_2243
timestamp 1677677812
transform 1 0 3276 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1969
timestamp 1677677812
transform 1 0 3292 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2315
timestamp 1677677812
transform 1 0 3292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2316
timestamp 1677677812
transform 1 0 3324 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1946
timestamp 1677677812
transform 1 0 3348 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2244
timestamp 1677677812
transform 1 0 3348 0 1 3625
box -2 -2 2 2
use M3_M2  M3_M2_1970
timestamp 1677677812
transform 1 0 3372 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2317
timestamp 1677677812
transform 1 0 3372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2318
timestamp 1677677812
transform 1 0 3388 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2414
timestamp 1677677812
transform 1 0 3364 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2018
timestamp 1677677812
transform 1 0 3372 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1971
timestamp 1677677812
transform 1 0 3412 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1972
timestamp 1677677812
transform 1 0 3436 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2001
timestamp 1677677812
transform 1 0 3428 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2319
timestamp 1677677812
transform 1 0 3436 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2415
timestamp 1677677812
transform 1 0 3420 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2416
timestamp 1677677812
transform 1 0 3428 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2019
timestamp 1677677812
transform 1 0 3436 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2417
timestamp 1677677812
transform 1 0 3444 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2418
timestamp 1677677812
transform 1 0 3460 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2039
timestamp 1677677812
transform 1 0 3460 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2320
timestamp 1677677812
transform 1 0 3484 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2040
timestamp 1677677812
transform 1 0 3484 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2321
timestamp 1677677812
transform 1 0 3500 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2020
timestamp 1677677812
transform 1 0 3500 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2419
timestamp 1677677812
transform 1 0 3516 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2002
timestamp 1677677812
transform 1 0 3532 0 1 3615
box -3 -3 3 3
use M3_M2  M3_M2_2021
timestamp 1677677812
transform 1 0 3556 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2041
timestamp 1677677812
transform 1 0 3556 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2022
timestamp 1677677812
transform 1 0 3596 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2322
timestamp 1677677812
transform 1 0 3700 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2420
timestamp 1677677812
transform 1 0 3652 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2323
timestamp 1677677812
transform 1 0 3740 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1947
timestamp 1677677812
transform 1 0 3772 0 1 3635
box -3 -3 3 3
use M2_M1  M2_M1_2324
timestamp 1677677812
transform 1 0 3772 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2421
timestamp 1677677812
transform 1 0 3756 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2422
timestamp 1677677812
transform 1 0 3764 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2023
timestamp 1677677812
transform 1 0 3772 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2423
timestamp 1677677812
transform 1 0 3788 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2424
timestamp 1677677812
transform 1 0 3796 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2042
timestamp 1677677812
transform 1 0 3764 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1973
timestamp 1677677812
transform 1 0 3876 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2325
timestamp 1677677812
transform 1 0 3876 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2326
timestamp 1677677812
transform 1 0 3884 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2043
timestamp 1677677812
transform 1 0 3884 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1917
timestamp 1677677812
transform 1 0 3900 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2425
timestamp 1677677812
transform 1 0 3916 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2327
timestamp 1677677812
transform 1 0 3948 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2328
timestamp 1677677812
transform 1 0 3964 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2426
timestamp 1677677812
transform 1 0 3956 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2427
timestamp 1677677812
transform 1 0 3972 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2428
timestamp 1677677812
transform 1 0 3988 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2429
timestamp 1677677812
transform 1 0 3996 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2061
timestamp 1677677812
transform 1 0 3956 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2329
timestamp 1677677812
transform 1 0 4012 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2330
timestamp 1677677812
transform 1 0 4028 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2331
timestamp 1677677812
transform 1 0 4060 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2430
timestamp 1677677812
transform 1 0 4052 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2024
timestamp 1677677812
transform 1 0 4060 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2431
timestamp 1677677812
transform 1 0 4068 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2044
timestamp 1677677812
transform 1 0 4044 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2062
timestamp 1677677812
transform 1 0 4068 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1918
timestamp 1677677812
transform 1 0 4108 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1937
timestamp 1677677812
transform 1 0 4100 0 1 3645
box -3 -3 3 3
use M2_M1  M2_M1_2237
timestamp 1677677812
transform 1 0 4092 0 1 3635
box -2 -2 2 2
use M2_M1  M2_M1_2245
timestamp 1677677812
transform 1 0 4084 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2332
timestamp 1677677812
transform 1 0 4100 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2045
timestamp 1677677812
transform 1 0 4092 0 1 3595
box -3 -3 3 3
use M2_M1  M2_M1_2246
timestamp 1677677812
transform 1 0 4116 0 1 3625
box -2 -2 2 2
use M2_M1  M2_M1_2333
timestamp 1677677812
transform 1 0 4124 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_2025
timestamp 1677677812
transform 1 0 4124 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_2063
timestamp 1677677812
transform 1 0 4116 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2432
timestamp 1677677812
transform 1 0 4140 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2046
timestamp 1677677812
transform 1 0 4140 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1919
timestamp 1677677812
transform 1 0 4156 0 1 3655
box -3 -3 3 3
use M3_M2  M3_M2_1920
timestamp 1677677812
transform 1 0 4188 0 1 3655
box -3 -3 3 3
use M2_M1  M2_M1_2334
timestamp 1677677812
transform 1 0 4180 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2433
timestamp 1677677812
transform 1 0 4156 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2047
timestamp 1677677812
transform 1 0 4172 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_1974
timestamp 1677677812
transform 1 0 4252 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2335
timestamp 1677677812
transform 1 0 4244 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2336
timestamp 1677677812
transform 1 0 4252 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1975
timestamp 1677677812
transform 1 0 4292 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2337
timestamp 1677677812
transform 1 0 4292 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2338
timestamp 1677677812
transform 1 0 4308 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2434
timestamp 1677677812
transform 1 0 4276 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2064
timestamp 1677677812
transform 1 0 4292 0 1 3585
box -3 -3 3 3
use M2_M1  M2_M1_2339
timestamp 1677677812
transform 1 0 4324 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1976
timestamp 1677677812
transform 1 0 4364 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2003
timestamp 1677677812
transform 1 0 4348 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2340
timestamp 1677677812
transform 1 0 4356 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2341
timestamp 1677677812
transform 1 0 4372 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2435
timestamp 1677677812
transform 1 0 4340 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2436
timestamp 1677677812
transform 1 0 4348 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2048
timestamp 1677677812
transform 1 0 4340 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2026
timestamp 1677677812
transform 1 0 4356 0 1 3605
box -3 -3 3 3
use M3_M2  M3_M2_1977
timestamp 1677677812
transform 1 0 4420 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2342
timestamp 1677677812
transform 1 0 4420 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2343
timestamp 1677677812
transform 1 0 4476 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2437
timestamp 1677677812
transform 1 0 4364 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2438
timestamp 1677677812
transform 1 0 4380 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2439
timestamp 1677677812
transform 1 0 4396 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2049
timestamp 1677677812
transform 1 0 4372 0 1 3595
box -3 -3 3 3
use M3_M2  M3_M2_2004
timestamp 1677677812
transform 1 0 4484 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2344
timestamp 1677677812
transform 1 0 4492 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2440
timestamp 1677677812
transform 1 0 4484 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2065
timestamp 1677677812
transform 1 0 4492 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1978
timestamp 1677677812
transform 1 0 4524 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2345
timestamp 1677677812
transform 1 0 4524 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2346
timestamp 1677677812
transform 1 0 4540 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2441
timestamp 1677677812
transform 1 0 4516 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2442
timestamp 1677677812
transform 1 0 4532 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2066
timestamp 1677677812
transform 1 0 4524 0 1 3585
box -3 -3 3 3
use M3_M2  M3_M2_1948
timestamp 1677677812
transform 1 0 4564 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1938
timestamp 1677677812
transform 1 0 4588 0 1 3645
box -3 -3 3 3
use M3_M2  M3_M2_1949
timestamp 1677677812
transform 1 0 4596 0 1 3635
box -3 -3 3 3
use M3_M2  M3_M2_1979
timestamp 1677677812
transform 1 0 4596 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_1980
timestamp 1677677812
transform 1 0 4612 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2347
timestamp 1677677812
transform 1 0 4572 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2348
timestamp 1677677812
transform 1 0 4588 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2349
timestamp 1677677812
transform 1 0 4604 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2350
timestamp 1677677812
transform 1 0 4612 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2443
timestamp 1677677812
transform 1 0 4580 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2027
timestamp 1677677812
transform 1 0 4588 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2444
timestamp 1677677812
transform 1 0 4596 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_1981
timestamp 1677677812
transform 1 0 4644 0 1 3625
box -3 -3 3 3
use M2_M1  M2_M1_2351
timestamp 1677677812
transform 1 0 4636 0 1 3615
box -2 -2 2 2
use M3_M2  M3_M2_1982
timestamp 1677677812
transform 1 0 4676 0 1 3625
box -3 -3 3 3
use M3_M2  M3_M2_2005
timestamp 1677677812
transform 1 0 4652 0 1 3615
box -3 -3 3 3
use M2_M1  M2_M1_2352
timestamp 1677677812
transform 1 0 4660 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2353
timestamp 1677677812
transform 1 0 4676 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2445
timestamp 1677677812
transform 1 0 4644 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2446
timestamp 1677677812
transform 1 0 4652 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2447
timestamp 1677677812
transform 1 0 4668 0 1 3605
box -2 -2 2 2
use M3_M2  M3_M2_2028
timestamp 1677677812
transform 1 0 4676 0 1 3605
box -3 -3 3 3
use M2_M1  M2_M1_2354
timestamp 1677677812
transform 1 0 4692 0 1 3615
box -2 -2 2 2
use M2_M1  M2_M1_2448
timestamp 1677677812
transform 1 0 4740 0 1 3605
box -2 -2 2 2
use M2_M1  M2_M1_2449
timestamp 1677677812
transform 1 0 4772 0 1 3605
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_22
timestamp 1677677812
transform 1 0 48 0 1 3570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_160
timestamp 1677677812
transform 1 0 72 0 1 3570
box -8 -3 104 105
use FILL  FILL_2219
timestamp 1677677812
transform 1 0 168 0 1 3570
box -8 -3 16 105
use FILL  FILL_2231
timestamp 1677677812
transform 1 0 176 0 1 3570
box -8 -3 16 105
use FILL  FILL_2232
timestamp 1677677812
transform 1 0 184 0 1 3570
box -8 -3 16 105
use FILL  FILL_2233
timestamp 1677677812
transform 1 0 192 0 1 3570
box -8 -3 16 105
use FILL  FILL_2234
timestamp 1677677812
transform 1 0 200 0 1 3570
box -8 -3 16 105
use FILL  FILL_2235
timestamp 1677677812
transform 1 0 208 0 1 3570
box -8 -3 16 105
use FILL  FILL_2236
timestamp 1677677812
transform 1 0 216 0 1 3570
box -8 -3 16 105
use FILL  FILL_2237
timestamp 1677677812
transform 1 0 224 0 1 3570
box -8 -3 16 105
use FILL  FILL_2240
timestamp 1677677812
transform 1 0 232 0 1 3570
box -8 -3 16 105
use FILL  FILL_2241
timestamp 1677677812
transform 1 0 240 0 1 3570
box -8 -3 16 105
use FILL  FILL_2242
timestamp 1677677812
transform 1 0 248 0 1 3570
box -8 -3 16 105
use FILL  FILL_2243
timestamp 1677677812
transform 1 0 256 0 1 3570
box -8 -3 16 105
use FILL  FILL_2244
timestamp 1677677812
transform 1 0 264 0 1 3570
box -8 -3 16 105
use FILL  FILL_2245
timestamp 1677677812
transform 1 0 272 0 1 3570
box -8 -3 16 105
use FILL  FILL_2246
timestamp 1677677812
transform 1 0 280 0 1 3570
box -8 -3 16 105
use FILL  FILL_2247
timestamp 1677677812
transform 1 0 288 0 1 3570
box -8 -3 16 105
use FILL  FILL_2248
timestamp 1677677812
transform 1 0 296 0 1 3570
box -8 -3 16 105
use FILL  FILL_2249
timestamp 1677677812
transform 1 0 304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2250
timestamp 1677677812
transform 1 0 312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2251
timestamp 1677677812
transform 1 0 320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2252
timestamp 1677677812
transform 1 0 328 0 1 3570
box -8 -3 16 105
use FILL  FILL_2253
timestamp 1677677812
transform 1 0 336 0 1 3570
box -8 -3 16 105
use FILL  FILL_2254
timestamp 1677677812
transform 1 0 344 0 1 3570
box -8 -3 16 105
use FILL  FILL_2256
timestamp 1677677812
transform 1 0 352 0 1 3570
box -8 -3 16 105
use FILL  FILL_2258
timestamp 1677677812
transform 1 0 360 0 1 3570
box -8 -3 16 105
use FILL  FILL_2260
timestamp 1677677812
transform 1 0 368 0 1 3570
box -8 -3 16 105
use FILL  FILL_2262
timestamp 1677677812
transform 1 0 376 0 1 3570
box -8 -3 16 105
use FILL  FILL_2263
timestamp 1677677812
transform 1 0 384 0 1 3570
box -8 -3 16 105
use FILL  FILL_2264
timestamp 1677677812
transform 1 0 392 0 1 3570
box -8 -3 16 105
use FILL  FILL_2265
timestamp 1677677812
transform 1 0 400 0 1 3570
box -8 -3 16 105
use FILL  FILL_2266
timestamp 1677677812
transform 1 0 408 0 1 3570
box -8 -3 16 105
use FILL  FILL_2267
timestamp 1677677812
transform 1 0 416 0 1 3570
box -8 -3 16 105
use FILL  FILL_2268
timestamp 1677677812
transform 1 0 424 0 1 3570
box -8 -3 16 105
use FILL  FILL_2271
timestamp 1677677812
transform 1 0 432 0 1 3570
box -8 -3 16 105
use FILL  FILL_2273
timestamp 1677677812
transform 1 0 440 0 1 3570
box -8 -3 16 105
use FILL  FILL_2275
timestamp 1677677812
transform 1 0 448 0 1 3570
box -8 -3 16 105
use FILL  FILL_2277
timestamp 1677677812
transform 1 0 456 0 1 3570
box -8 -3 16 105
use FILL  FILL_2279
timestamp 1677677812
transform 1 0 464 0 1 3570
box -8 -3 16 105
use FILL  FILL_2281
timestamp 1677677812
transform 1 0 472 0 1 3570
box -8 -3 16 105
use FILL  FILL_2283
timestamp 1677677812
transform 1 0 480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2284
timestamp 1677677812
transform 1 0 488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2285
timestamp 1677677812
transform 1 0 496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2286
timestamp 1677677812
transform 1 0 504 0 1 3570
box -8 -3 16 105
use FILL  FILL_2287
timestamp 1677677812
transform 1 0 512 0 1 3570
box -8 -3 16 105
use FILL  FILL_2288
timestamp 1677677812
transform 1 0 520 0 1 3570
box -8 -3 16 105
use FILL  FILL_2290
timestamp 1677677812
transform 1 0 528 0 1 3570
box -8 -3 16 105
use FILL  FILL_2292
timestamp 1677677812
transform 1 0 536 0 1 3570
box -8 -3 16 105
use FILL  FILL_2294
timestamp 1677677812
transform 1 0 544 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_190
timestamp 1677677812
transform 1 0 552 0 1 3570
box -9 -3 26 105
use FILL  FILL_2296
timestamp 1677677812
transform 1 0 568 0 1 3570
box -8 -3 16 105
use FILL  FILL_2300
timestamp 1677677812
transform 1 0 576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2302
timestamp 1677677812
transform 1 0 584 0 1 3570
box -8 -3 16 105
use FILL  FILL_2304
timestamp 1677677812
transform 1 0 592 0 1 3570
box -8 -3 16 105
use FILL  FILL_2306
timestamp 1677677812
transform 1 0 600 0 1 3570
box -8 -3 16 105
use FILL  FILL_2307
timestamp 1677677812
transform 1 0 608 0 1 3570
box -8 -3 16 105
use FILL  FILL_2308
timestamp 1677677812
transform 1 0 616 0 1 3570
box -8 -3 16 105
use FILL  FILL_2309
timestamp 1677677812
transform 1 0 624 0 1 3570
box -8 -3 16 105
use FILL  FILL_2310
timestamp 1677677812
transform 1 0 632 0 1 3570
box -8 -3 16 105
use FILL  FILL_2311
timestamp 1677677812
transform 1 0 640 0 1 3570
box -8 -3 16 105
use FILL  FILL_2314
timestamp 1677677812
transform 1 0 648 0 1 3570
box -8 -3 16 105
use FILL  FILL_2316
timestamp 1677677812
transform 1 0 656 0 1 3570
box -8 -3 16 105
use FILL  FILL_2317
timestamp 1677677812
transform 1 0 664 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2067
timestamp 1677677812
transform 1 0 684 0 1 3575
box -3 -3 3 3
use FILL  FILL_2318
timestamp 1677677812
transform 1 0 672 0 1 3570
box -8 -3 16 105
use FILL  FILL_2319
timestamp 1677677812
transform 1 0 680 0 1 3570
box -8 -3 16 105
use FILL  FILL_2320
timestamp 1677677812
transform 1 0 688 0 1 3570
box -8 -3 16 105
use FILL  FILL_2321
timestamp 1677677812
transform 1 0 696 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_162
timestamp 1677677812
transform 1 0 704 0 1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_163
timestamp 1677677812
transform 1 0 800 0 1 3570
box -8 -3 104 105
use FILL  FILL_2324
timestamp 1677677812
transform 1 0 896 0 1 3570
box -8 -3 16 105
use FILL  FILL_2325
timestamp 1677677812
transform 1 0 904 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_106
timestamp 1677677812
transform -1 0 952 0 1 3570
box -8 -3 46 105
use FILL  FILL_2326
timestamp 1677677812
transform 1 0 952 0 1 3570
box -8 -3 16 105
use FILL  FILL_2348
timestamp 1677677812
transform 1 0 960 0 1 3570
box -8 -3 16 105
use FILL  FILL_2350
timestamp 1677677812
transform 1 0 968 0 1 3570
box -8 -3 16 105
use FILL  FILL_2351
timestamp 1677677812
transform 1 0 976 0 1 3570
box -8 -3 16 105
use FILL  FILL_2352
timestamp 1677677812
transform 1 0 984 0 1 3570
box -8 -3 16 105
use FILL  FILL_2353
timestamp 1677677812
transform 1 0 992 0 1 3570
box -8 -3 16 105
use FILL  FILL_2354
timestamp 1677677812
transform 1 0 1000 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_192
timestamp 1677677812
transform -1 0 1024 0 1 3570
box -9 -3 26 105
use FILL  FILL_2355
timestamp 1677677812
transform 1 0 1024 0 1 3570
box -8 -3 16 105
use FILL  FILL_2356
timestamp 1677677812
transform 1 0 1032 0 1 3570
box -8 -3 16 105
use FILL  FILL_2357
timestamp 1677677812
transform 1 0 1040 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_107
timestamp 1677677812
transform -1 0 1088 0 1 3570
box -8 -3 46 105
use FILL  FILL_2358
timestamp 1677677812
transform 1 0 1088 0 1 3570
box -8 -3 16 105
use FILL  FILL_2363
timestamp 1677677812
transform 1 0 1096 0 1 3570
box -8 -3 16 105
use FILL  FILL_2364
timestamp 1677677812
transform 1 0 1104 0 1 3570
box -8 -3 16 105
use FILL  FILL_2365
timestamp 1677677812
transform 1 0 1112 0 1 3570
box -8 -3 16 105
use FILL  FILL_2366
timestamp 1677677812
transform 1 0 1120 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_193
timestamp 1677677812
transform -1 0 1144 0 1 3570
box -9 -3 26 105
use FILL  FILL_2367
timestamp 1677677812
transform 1 0 1144 0 1 3570
box -8 -3 16 105
use FILL  FILL_2368
timestamp 1677677812
transform 1 0 1152 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_108
timestamp 1677677812
transform 1 0 1160 0 1 3570
box -8 -3 46 105
use FILL  FILL_2369
timestamp 1677677812
transform 1 0 1200 0 1 3570
box -8 -3 16 105
use FILL  FILL_2372
timestamp 1677677812
transform 1 0 1208 0 1 3570
box -8 -3 16 105
use FILL  FILL_2374
timestamp 1677677812
transform 1 0 1216 0 1 3570
box -8 -3 16 105
use FILL  FILL_2375
timestamp 1677677812
transform 1 0 1224 0 1 3570
box -8 -3 16 105
use FILL  FILL_2376
timestamp 1677677812
transform 1 0 1232 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_53
timestamp 1677677812
transform -1 0 1272 0 1 3570
box -8 -3 34 105
use FILL  FILL_2377
timestamp 1677677812
transform 1 0 1272 0 1 3570
box -8 -3 16 105
use FILL  FILL_2378
timestamp 1677677812
transform 1 0 1280 0 1 3570
box -8 -3 16 105
use FILL  FILL_2379
timestamp 1677677812
transform 1 0 1288 0 1 3570
box -8 -3 16 105
use FILL  FILL_2380
timestamp 1677677812
transform 1 0 1296 0 1 3570
box -8 -3 16 105
use FILL  FILL_2381
timestamp 1677677812
transform 1 0 1304 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1677677812
transform 1 0 1312 0 1 3570
box -8 -3 32 105
use FILL  FILL_2382
timestamp 1677677812
transform 1 0 1336 0 1 3570
box -8 -3 16 105
use FILL  FILL_2392
timestamp 1677677812
transform 1 0 1344 0 1 3570
box -8 -3 16 105
use FILL  FILL_2393
timestamp 1677677812
transform 1 0 1352 0 1 3570
box -8 -3 16 105
use FILL  FILL_2394
timestamp 1677677812
transform 1 0 1360 0 1 3570
box -8 -3 16 105
use FILL  FILL_2395
timestamp 1677677812
transform 1 0 1368 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_166
timestamp 1677677812
transform -1 0 1472 0 1 3570
box -8 -3 104 105
use FILL  FILL_2396
timestamp 1677677812
transform 1 0 1472 0 1 3570
box -8 -3 16 105
use FILL  FILL_2408
timestamp 1677677812
transform 1 0 1480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2410
timestamp 1677677812
transform 1 0 1488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2412
timestamp 1677677812
transform 1 0 1496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2414
timestamp 1677677812
transform 1 0 1504 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_100
timestamp 1677677812
transform -1 0 1552 0 1 3570
box -8 -3 46 105
use FILL  FILL_2415
timestamp 1677677812
transform 1 0 1552 0 1 3570
box -8 -3 16 105
use FILL  FILL_2416
timestamp 1677677812
transform 1 0 1560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2417
timestamp 1677677812
transform 1 0 1568 0 1 3570
box -8 -3 16 105
use FILL  FILL_2422
timestamp 1677677812
transform 1 0 1576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2424
timestamp 1677677812
transform 1 0 1584 0 1 3570
box -8 -3 16 105
use FILL  FILL_2426
timestamp 1677677812
transform 1 0 1592 0 1 3570
box -8 -3 16 105
use FILL  FILL_2428
timestamp 1677677812
transform 1 0 1600 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_195
timestamp 1677677812
transform -1 0 1624 0 1 3570
box -9 -3 26 105
use M3_M2  M3_M2_2068
timestamp 1677677812
transform 1 0 1692 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2069
timestamp 1677677812
transform 1 0 1724 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_167
timestamp 1677677812
transform 1 0 1624 0 1 3570
box -8 -3 104 105
use FILL  FILL_2429
timestamp 1677677812
transform 1 0 1720 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_196
timestamp 1677677812
transform 1 0 1728 0 1 3570
box -9 -3 26 105
use FILL  FILL_2430
timestamp 1677677812
transform 1 0 1744 0 1 3570
box -8 -3 16 105
use FILL  FILL_2441
timestamp 1677677812
transform 1 0 1752 0 1 3570
box -8 -3 16 105
use FILL  FILL_2443
timestamp 1677677812
transform 1 0 1760 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2070
timestamp 1677677812
transform 1 0 1780 0 1 3575
box -3 -3 3 3
use FILL  FILL_2444
timestamp 1677677812
transform 1 0 1768 0 1 3570
box -8 -3 16 105
use BUFX2  BUFX2_15
timestamp 1677677812
transform 1 0 1776 0 1 3570
box -5 -3 28 105
use FILL  FILL_2445
timestamp 1677677812
transform 1 0 1800 0 1 3570
box -8 -3 16 105
use FILL  FILL_2447
timestamp 1677677812
transform 1 0 1808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2449
timestamp 1677677812
transform 1 0 1816 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_197
timestamp 1677677812
transform -1 0 1840 0 1 3570
box -9 -3 26 105
use FILL  FILL_2450
timestamp 1677677812
transform 1 0 1840 0 1 3570
box -8 -3 16 105
use FILL  FILL_2451
timestamp 1677677812
transform 1 0 1848 0 1 3570
box -8 -3 16 105
use FILL  FILL_2452
timestamp 1677677812
transform 1 0 1856 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_109
timestamp 1677677812
transform -1 0 1904 0 1 3570
box -8 -3 46 105
use FILL  FILL_2453
timestamp 1677677812
transform 1 0 1904 0 1 3570
box -8 -3 16 105
use FILL  FILL_2454
timestamp 1677677812
transform 1 0 1912 0 1 3570
box -8 -3 16 105
use FILL  FILL_2455
timestamp 1677677812
transform 1 0 1920 0 1 3570
box -8 -3 16 105
use FILL  FILL_2456
timestamp 1677677812
transform 1 0 1928 0 1 3570
box -8 -3 16 105
use FILL  FILL_2457
timestamp 1677677812
transform 1 0 1936 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_110
timestamp 1677677812
transform 1 0 1944 0 1 3570
box -8 -3 46 105
use FILL  FILL_2458
timestamp 1677677812
transform 1 0 1984 0 1 3570
box -8 -3 16 105
use FILL  FILL_2467
timestamp 1677677812
transform 1 0 1992 0 1 3570
box -8 -3 16 105
use FILL  FILL_2468
timestamp 1677677812
transform 1 0 2000 0 1 3570
box -8 -3 16 105
use FILL  FILL_2469
timestamp 1677677812
transform 1 0 2008 0 1 3570
box -8 -3 16 105
use FILL  FILL_2471
timestamp 1677677812
transform 1 0 2016 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_111
timestamp 1677677812
transform 1 0 2024 0 1 3570
box -8 -3 46 105
use FILL  FILL_2473
timestamp 1677677812
transform 1 0 2064 0 1 3570
box -8 -3 16 105
use FILL  FILL_2474
timestamp 1677677812
transform 1 0 2072 0 1 3570
box -8 -3 16 105
use FILL  FILL_2475
timestamp 1677677812
transform 1 0 2080 0 1 3570
box -8 -3 16 105
use FILL  FILL_2476
timestamp 1677677812
transform 1 0 2088 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_104
timestamp 1677677812
transform -1 0 2136 0 1 3570
box -8 -3 46 105
use FILL  FILL_2477
timestamp 1677677812
transform 1 0 2136 0 1 3570
box -8 -3 16 105
use FILL  FILL_2478
timestamp 1677677812
transform 1 0 2144 0 1 3570
box -8 -3 16 105
use FILL  FILL_2479
timestamp 1677677812
transform 1 0 2152 0 1 3570
box -8 -3 16 105
use FILL  FILL_2480
timestamp 1677677812
transform 1 0 2160 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_200
timestamp 1677677812
transform -1 0 2184 0 1 3570
box -9 -3 26 105
use FILL  FILL_2481
timestamp 1677677812
transform 1 0 2184 0 1 3570
box -8 -3 16 105
use FILL  FILL_2482
timestamp 1677677812
transform 1 0 2192 0 1 3570
box -8 -3 16 105
use FILL  FILL_2483
timestamp 1677677812
transform 1 0 2200 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_169
timestamp 1677677812
transform 1 0 2208 0 1 3570
box -8 -3 104 105
use FILL  FILL_2484
timestamp 1677677812
transform 1 0 2304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2485
timestamp 1677677812
transform 1 0 2312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2486
timestamp 1677677812
transform 1 0 2320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2487
timestamp 1677677812
transform 1 0 2328 0 1 3570
box -8 -3 16 105
use FILL  FILL_2488
timestamp 1677677812
transform 1 0 2336 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_112
timestamp 1677677812
transform -1 0 2384 0 1 3570
box -8 -3 46 105
use FILL  FILL_2489
timestamp 1677677812
transform 1 0 2384 0 1 3570
box -8 -3 16 105
use FILL  FILL_2490
timestamp 1677677812
transform 1 0 2392 0 1 3570
box -8 -3 16 105
use FILL  FILL_2491
timestamp 1677677812
transform 1 0 2400 0 1 3570
box -8 -3 16 105
use FILL  FILL_2492
timestamp 1677677812
transform 1 0 2408 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2071
timestamp 1677677812
transform 1 0 2428 0 1 3575
box -3 -3 3 3
use M3_M2  M3_M2_2072
timestamp 1677677812
transform 1 0 2444 0 1 3575
box -3 -3 3 3
use INVX2  INVX2_201
timestamp 1677677812
transform 1 0 2416 0 1 3570
box -9 -3 26 105
use M3_M2  M3_M2_2073
timestamp 1677677812
transform 1 0 2484 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_170
timestamp 1677677812
transform -1 0 2528 0 1 3570
box -8 -3 104 105
use OAI21X1  OAI21X1_56
timestamp 1677677812
transform 1 0 2528 0 1 3570
box -8 -3 34 105
use FILL  FILL_2493
timestamp 1677677812
transform 1 0 2560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2513
timestamp 1677677812
transform 1 0 2568 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_173
timestamp 1677677812
transform 1 0 2576 0 1 3570
box -8 -3 104 105
use FILL  FILL_2515
timestamp 1677677812
transform 1 0 2672 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_174
timestamp 1677677812
transform -1 0 2776 0 1 3570
box -8 -3 104 105
use FILL  FILL_2516
timestamp 1677677812
transform 1 0 2776 0 1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_57
timestamp 1677677812
transform 1 0 2784 0 1 3570
box -8 -3 34 105
use FILL  FILL_2531
timestamp 1677677812
transform 1 0 2816 0 1 3570
box -8 -3 16 105
use FILL  FILL_2533
timestamp 1677677812
transform 1 0 2824 0 1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_27
timestamp 1677677812
transform 1 0 2832 0 1 3570
box -8 -3 32 105
use FILL  FILL_2535
timestamp 1677677812
transform 1 0 2856 0 1 3570
box -8 -3 16 105
use FILL  FILL_2540
timestamp 1677677812
transform 1 0 2864 0 1 3570
box -8 -3 16 105
use FILL  FILL_2542
timestamp 1677677812
transform 1 0 2872 0 1 3570
box -8 -3 16 105
use FILL  FILL_2543
timestamp 1677677812
transform 1 0 2880 0 1 3570
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1677677812
transform -1 0 2912 0 1 3570
box -8 -3 32 105
use OAI21X1  OAI21X1_59
timestamp 1677677812
transform -1 0 2944 0 1 3570
box -8 -3 34 105
use FILL  FILL_2544
timestamp 1677677812
transform 1 0 2944 0 1 3570
box -8 -3 16 105
use FILL  FILL_2545
timestamp 1677677812
transform 1 0 2952 0 1 3570
box -8 -3 16 105
use FILL  FILL_2546
timestamp 1677677812
transform 1 0 2960 0 1 3570
box -8 -3 16 105
use FILL  FILL_2547
timestamp 1677677812
transform 1 0 2968 0 1 3570
box -8 -3 16 105
use FILL  FILL_2548
timestamp 1677677812
transform 1 0 2976 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2074
timestamp 1677677812
transform 1 0 3084 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_175
timestamp 1677677812
transform 1 0 2984 0 1 3570
box -8 -3 104 105
use FILL  FILL_2549
timestamp 1677677812
transform 1 0 3080 0 1 3570
box -8 -3 16 105
use FILL  FILL_2560
timestamp 1677677812
transform 1 0 3088 0 1 3570
box -8 -3 16 105
use FILL  FILL_2562
timestamp 1677677812
transform 1 0 3096 0 1 3570
box -8 -3 16 105
use FILL  FILL_2564
timestamp 1677677812
transform 1 0 3104 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_106
timestamp 1677677812
transform -1 0 3152 0 1 3570
box -8 -3 46 105
use FILL  FILL_2565
timestamp 1677677812
transform 1 0 3152 0 1 3570
box -8 -3 16 105
use FILL  FILL_2571
timestamp 1677677812
transform 1 0 3160 0 1 3570
box -8 -3 16 105
use FILL  FILL_2572
timestamp 1677677812
transform 1 0 3168 0 1 3570
box -8 -3 16 105
use FILL  FILL_2573
timestamp 1677677812
transform 1 0 3176 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2075
timestamp 1677677812
transform 1 0 3196 0 1 3575
box -3 -3 3 3
use FILL  FILL_2574
timestamp 1677677812
transform 1 0 3184 0 1 3570
box -8 -3 16 105
use FILL  FILL_2575
timestamp 1677677812
transform 1 0 3192 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_207
timestamp 1677677812
transform -1 0 3216 0 1 3570
box -9 -3 26 105
use FILL  FILL_2576
timestamp 1677677812
transform 1 0 3216 0 1 3570
box -8 -3 16 105
use FILL  FILL_2580
timestamp 1677677812
transform 1 0 3224 0 1 3570
box -8 -3 16 105
use FILL  FILL_2582
timestamp 1677677812
transform 1 0 3232 0 1 3570
box -8 -3 16 105
use FILL  FILL_2583
timestamp 1677677812
transform 1 0 3240 0 1 3570
box -8 -3 16 105
use FILL  FILL_2584
timestamp 1677677812
transform 1 0 3248 0 1 3570
box -8 -3 16 105
use FILL  FILL_2585
timestamp 1677677812
transform 1 0 3256 0 1 3570
box -8 -3 16 105
use FILL  FILL_2586
timestamp 1677677812
transform 1 0 3264 0 1 3570
box -8 -3 16 105
use NAND3X1  NAND3X1_11
timestamp 1677677812
transform -1 0 3304 0 1 3570
box -8 -3 40 105
use FILL  FILL_2587
timestamp 1677677812
transform 1 0 3304 0 1 3570
box -8 -3 16 105
use FILL  FILL_2594
timestamp 1677677812
transform 1 0 3312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2596
timestamp 1677677812
transform 1 0 3320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2598
timestamp 1677677812
transform 1 0 3328 0 1 3570
box -8 -3 16 105
use FILL  FILL_2599
timestamp 1677677812
transform 1 0 3336 0 1 3570
box -8 -3 16 105
use FILL  FILL_2600
timestamp 1677677812
transform 1 0 3344 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_118
timestamp 1677677812
transform 1 0 3352 0 1 3570
box -8 -3 46 105
use FILL  FILL_2601
timestamp 1677677812
transform 1 0 3392 0 1 3570
box -8 -3 16 105
use FILL  FILL_2606
timestamp 1677677812
transform 1 0 3400 0 1 3570
box -8 -3 16 105
use FILL  FILL_2608
timestamp 1677677812
transform 1 0 3408 0 1 3570
box -8 -3 16 105
use FILL  FILL_2610
timestamp 1677677812
transform 1 0 3416 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_108
timestamp 1677677812
transform -1 0 3464 0 1 3570
box -8 -3 46 105
use FILL  FILL_2611
timestamp 1677677812
transform 1 0 3464 0 1 3570
box -8 -3 16 105
use FILL  FILL_2612
timestamp 1677677812
transform 1 0 3472 0 1 3570
box -8 -3 16 105
use FILL  FILL_2613
timestamp 1677677812
transform 1 0 3480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2614
timestamp 1677677812
transform 1 0 3488 0 1 3570
box -8 -3 16 105
use FILL  FILL_2615
timestamp 1677677812
transform 1 0 3496 0 1 3570
box -8 -3 16 105
use FILL  FILL_2616
timestamp 1677677812
transform 1 0 3504 0 1 3570
box -8 -3 16 105
use FILL  FILL_2617
timestamp 1677677812
transform 1 0 3512 0 1 3570
box -8 -3 16 105
use FILL  FILL_2619
timestamp 1677677812
transform 1 0 3520 0 1 3570
box -8 -3 16 105
use FILL  FILL_2620
timestamp 1677677812
transform 1 0 3528 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_208
timestamp 1677677812
transform 1 0 3536 0 1 3570
box -9 -3 26 105
use FILL  FILL_2621
timestamp 1677677812
transform 1 0 3552 0 1 3570
box -8 -3 16 105
use FILL  FILL_2622
timestamp 1677677812
transform 1 0 3560 0 1 3570
box -8 -3 16 105
use FILL  FILL_2623
timestamp 1677677812
transform 1 0 3568 0 1 3570
box -8 -3 16 105
use FILL  FILL_2626
timestamp 1677677812
transform 1 0 3576 0 1 3570
box -8 -3 16 105
use FILL  FILL_2628
timestamp 1677677812
transform 1 0 3584 0 1 3570
box -8 -3 16 105
use FILL  FILL_2630
timestamp 1677677812
transform 1 0 3592 0 1 3570
box -8 -3 16 105
use FILL  FILL_2632
timestamp 1677677812
transform 1 0 3600 0 1 3570
box -8 -3 16 105
use FILL  FILL_2634
timestamp 1677677812
transform 1 0 3608 0 1 3570
box -8 -3 16 105
use FILL  FILL_2635
timestamp 1677677812
transform 1 0 3616 0 1 3570
box -8 -3 16 105
use FILL  FILL_2636
timestamp 1677677812
transform 1 0 3624 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2076
timestamp 1677677812
transform 1 0 3644 0 1 3575
box -3 -3 3 3
use FILL  FILL_2638
timestamp 1677677812
transform 1 0 3632 0 1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_177
timestamp 1677677812
transform 1 0 3640 0 1 3570
box -8 -3 104 105
use FILL  FILL_2640
timestamp 1677677812
transform 1 0 3736 0 1 3570
box -8 -3 16 105
use FILL  FILL_2649
timestamp 1677677812
transform 1 0 3744 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_120
timestamp 1677677812
transform 1 0 3752 0 1 3570
box -8 -3 46 105
use FILL  FILL_2651
timestamp 1677677812
transform 1 0 3792 0 1 3570
box -8 -3 16 105
use FILL  FILL_2652
timestamp 1677677812
transform 1 0 3800 0 1 3570
box -8 -3 16 105
use FILL  FILL_2655
timestamp 1677677812
transform 1 0 3808 0 1 3570
box -8 -3 16 105
use FILL  FILL_2657
timestamp 1677677812
transform 1 0 3816 0 1 3570
box -8 -3 16 105
use FILL  FILL_2658
timestamp 1677677812
transform 1 0 3824 0 1 3570
box -8 -3 16 105
use FILL  FILL_2659
timestamp 1677677812
transform 1 0 3832 0 1 3570
box -8 -3 16 105
use FILL  FILL_2660
timestamp 1677677812
transform 1 0 3840 0 1 3570
box -8 -3 16 105
use FILL  FILL_2661
timestamp 1677677812
transform 1 0 3848 0 1 3570
box -8 -3 16 105
use FILL  FILL_2662
timestamp 1677677812
transform 1 0 3856 0 1 3570
box -8 -3 16 105
use FILL  FILL_2664
timestamp 1677677812
transform 1 0 3864 0 1 3570
box -8 -3 16 105
use FILL  FILL_2666
timestamp 1677677812
transform 1 0 3872 0 1 3570
box -8 -3 16 105
use FILL  FILL_2668
timestamp 1677677812
transform 1 0 3880 0 1 3570
box -8 -3 16 105
use FILL  FILL_2670
timestamp 1677677812
transform 1 0 3888 0 1 3570
box -8 -3 16 105
use FILL  FILL_2671
timestamp 1677677812
transform 1 0 3896 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_210
timestamp 1677677812
transform -1 0 3920 0 1 3570
box -9 -3 26 105
use FILL  FILL_2672
timestamp 1677677812
transform 1 0 3920 0 1 3570
box -8 -3 16 105
use FILL  FILL_2673
timestamp 1677677812
transform 1 0 3928 0 1 3570
box -8 -3 16 105
use FILL  FILL_2674
timestamp 1677677812
transform 1 0 3936 0 1 3570
box -8 -3 16 105
use FILL  FILL_2675
timestamp 1677677812
transform 1 0 3944 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_112
timestamp 1677677812
transform -1 0 3992 0 1 3570
box -8 -3 46 105
use FILL  FILL_2676
timestamp 1677677812
transform 1 0 3992 0 1 3570
box -8 -3 16 105
use FILL  FILL_2677
timestamp 1677677812
transform 1 0 4000 0 1 3570
box -8 -3 16 105
use FILL  FILL_2679
timestamp 1677677812
transform 1 0 4008 0 1 3570
box -8 -3 16 105
use FILL  FILL_2681
timestamp 1677677812
transform 1 0 4016 0 1 3570
box -8 -3 16 105
use FILL  FILL_2683
timestamp 1677677812
transform 1 0 4024 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_113
timestamp 1677677812
transform 1 0 4032 0 1 3570
box -8 -3 46 105
use M3_M2  M3_M2_2077
timestamp 1677677812
transform 1 0 4084 0 1 3575
box -3 -3 3 3
use FILL  FILL_2685
timestamp 1677677812
transform 1 0 4072 0 1 3570
box -8 -3 16 105
use NAND3X1  NAND3X1_13
timestamp 1677677812
transform -1 0 4112 0 1 3570
box -8 -3 40 105
use FILL  FILL_2686
timestamp 1677677812
transform 1 0 4112 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2078
timestamp 1677677812
transform 1 0 4140 0 1 3575
box -3 -3 3 3
use INVX2  INVX2_212
timestamp 1677677812
transform -1 0 4136 0 1 3570
box -9 -3 26 105
use FILL  FILL_2687
timestamp 1677677812
transform 1 0 4136 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2079
timestamp 1677677812
transform 1 0 4196 0 1 3575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_179
timestamp 1677677812
transform 1 0 4144 0 1 3570
box -8 -3 104 105
use FILL  FILL_2688
timestamp 1677677812
transform 1 0 4240 0 1 3570
box -8 -3 16 105
use FILL  FILL_2689
timestamp 1677677812
transform 1 0 4248 0 1 3570
box -8 -3 16 105
use FILL  FILL_2690
timestamp 1677677812
transform 1 0 4256 0 1 3570
box -8 -3 16 105
use FILL  FILL_2691
timestamp 1677677812
transform 1 0 4264 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_122
timestamp 1677677812
transform -1 0 4312 0 1 3570
box -8 -3 46 105
use FILL  FILL_2692
timestamp 1677677812
transform 1 0 4312 0 1 3570
box -8 -3 16 105
use FILL  FILL_2693
timestamp 1677677812
transform 1 0 4320 0 1 3570
box -8 -3 16 105
use FILL  FILL_2694
timestamp 1677677812
transform 1 0 4328 0 1 3570
box -8 -3 16 105
use FILL  FILL_2695
timestamp 1677677812
transform 1 0 4336 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_114
timestamp 1677677812
transform 1 0 4344 0 1 3570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_180
timestamp 1677677812
transform 1 0 4384 0 1 3570
box -8 -3 104 105
use M3_M2  M3_M2_2080
timestamp 1677677812
transform 1 0 4492 0 1 3575
box -3 -3 3 3
use FILL  FILL_2696
timestamp 1677677812
transform 1 0 4480 0 1 3570
box -8 -3 16 105
use FILL  FILL_2711
timestamp 1677677812
transform 1 0 4488 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_116
timestamp 1677677812
transform 1 0 4496 0 1 3570
box -8 -3 46 105
use FILL  FILL_2712
timestamp 1677677812
transform 1 0 4536 0 1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2081
timestamp 1677677812
transform 1 0 4556 0 1 3575
box -3 -3 3 3
use FILL  FILL_2715
timestamp 1677677812
transform 1 0 4544 0 1 3570
box -8 -3 16 105
use FILL  FILL_2717
timestamp 1677677812
transform 1 0 4552 0 1 3570
box -8 -3 16 105
use FILL  FILL_2719
timestamp 1677677812
transform 1 0 4560 0 1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_123
timestamp 1677677812
transform 1 0 4568 0 1 3570
box -8 -3 46 105
use INVX2  INVX2_214
timestamp 1677677812
transform -1 0 4624 0 1 3570
box -9 -3 26 105
use FILL  FILL_2720
timestamp 1677677812
transform 1 0 4624 0 1 3570
box -8 -3 16 105
use FILL  FILL_2721
timestamp 1677677812
transform 1 0 4632 0 1 3570
box -8 -3 16 105
use FILL  FILL_2722
timestamp 1677677812
transform 1 0 4640 0 1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_118
timestamp 1677677812
transform 1 0 4648 0 1 3570
box -8 -3 46 105
use FILL  FILL_2723
timestamp 1677677812
transform 1 0 4688 0 1 3570
box -8 -3 16 105
use FILL  FILL_2724
timestamp 1677677812
transform 1 0 4696 0 1 3570
box -8 -3 16 105
use FILL  FILL_2725
timestamp 1677677812
transform 1 0 4704 0 1 3570
box -8 -3 16 105
use FILL  FILL_2726
timestamp 1677677812
transform 1 0 4712 0 1 3570
box -8 -3 16 105
use FILL  FILL_2727
timestamp 1677677812
transform 1 0 4720 0 1 3570
box -8 -3 16 105
use FILL  FILL_2728
timestamp 1677677812
transform 1 0 4728 0 1 3570
box -8 -3 16 105
use FILL  FILL_2729
timestamp 1677677812
transform 1 0 4736 0 1 3570
box -8 -3 16 105
use INVX2  INVX2_215
timestamp 1677677812
transform -1 0 4760 0 1 3570
box -9 -3 26 105
use FILL  FILL_2730
timestamp 1677677812
transform 1 0 4760 0 1 3570
box -8 -3 16 105
use FILL  FILL_2731
timestamp 1677677812
transform 1 0 4768 0 1 3570
box -8 -3 16 105
use FILL  FILL_2732
timestamp 1677677812
transform 1 0 4776 0 1 3570
box -8 -3 16 105
use FILL  FILL_2733
timestamp 1677677812
transform 1 0 4784 0 1 3570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_23
timestamp 1677677812
transform 1 0 4819 0 1 3570
box -10 -3 10 3
use M2_M1  M2_M1_2550
timestamp 1677677812
transform 1 0 124 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2452
timestamp 1677677812
transform 1 0 188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2453
timestamp 1677677812
transform 1 0 196 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2121
timestamp 1677677812
transform 1 0 228 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2454
timestamp 1677677812
transform 1 0 228 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2551
timestamp 1677677812
transform 1 0 188 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2552
timestamp 1677677812
transform 1 0 204 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2553
timestamp 1677677812
transform 1 0 220 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2210
timestamp 1677677812
transform 1 0 188 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2177
timestamp 1677677812
transform 1 0 228 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2082
timestamp 1677677812
transform 1 0 244 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2101
timestamp 1677677812
transform 1 0 244 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2102
timestamp 1677677812
transform 1 0 340 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2122
timestamp 1677677812
transform 1 0 332 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2455
timestamp 1677677812
transform 1 0 244 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2160
timestamp 1677677812
transform 1 0 268 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2161
timestamp 1677677812
transform 1 0 332 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2554
timestamp 1677677812
transform 1 0 268 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2178
timestamp 1677677812
transform 1 0 316 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2555
timestamp 1677677812
transform 1 0 324 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2556
timestamp 1677677812
transform 1 0 332 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2557
timestamp 1677677812
transform 1 0 340 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2211
timestamp 1677677812
transform 1 0 340 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2123
timestamp 1677677812
transform 1 0 412 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2456
timestamp 1677677812
transform 1 0 388 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2457
timestamp 1677677812
transform 1 0 396 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2458
timestamp 1677677812
transform 1 0 412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2558
timestamp 1677677812
transform 1 0 388 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2179
timestamp 1677677812
transform 1 0 396 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2559
timestamp 1677677812
transform 1 0 404 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2180
timestamp 1677677812
transform 1 0 412 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2237
timestamp 1677677812
transform 1 0 388 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2560
timestamp 1677677812
transform 1 0 428 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2561
timestamp 1677677812
transform 1 0 444 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2083
timestamp 1677677812
transform 1 0 460 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2562
timestamp 1677677812
transform 1 0 460 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2212
timestamp 1677677812
transform 1 0 468 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2124
timestamp 1677677812
transform 1 0 492 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2459
timestamp 1677677812
transform 1 0 492 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2125
timestamp 1677677812
transform 1 0 524 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2563
timestamp 1677677812
transform 1 0 500 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2564
timestamp 1677677812
transform 1 0 516 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2565
timestamp 1677677812
transform 1 0 524 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2213
timestamp 1677677812
transform 1 0 492 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2238
timestamp 1677677812
transform 1 0 516 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2126
timestamp 1677677812
transform 1 0 604 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2460
timestamp 1677677812
transform 1 0 604 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2084
timestamp 1677677812
transform 1 0 636 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2103
timestamp 1677677812
transform 1 0 636 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2566
timestamp 1677677812
transform 1 0 628 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2567
timestamp 1677677812
transform 1 0 644 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2461
timestamp 1677677812
transform 1 0 660 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2462
timestamp 1677677812
transform 1 0 692 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2568
timestamp 1677677812
transform 1 0 684 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2127
timestamp 1677677812
transform 1 0 708 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2463
timestamp 1677677812
transform 1 0 708 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2181
timestamp 1677677812
transform 1 0 740 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2464
timestamp 1677677812
transform 1 0 780 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2162
timestamp 1677677812
transform 1 0 788 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2465
timestamp 1677677812
transform 1 0 796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2569
timestamp 1677677812
transform 1 0 772 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2570
timestamp 1677677812
transform 1 0 796 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2264
timestamp 1677677812
transform 1 0 796 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2571
timestamp 1677677812
transform 1 0 836 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2128
timestamp 1677677812
transform 1 0 868 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2466
timestamp 1677677812
transform 1 0 868 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2467
timestamp 1677677812
transform 1 0 892 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2572
timestamp 1677677812
transform 1 0 884 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2129
timestamp 1677677812
transform 1 0 932 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2468
timestamp 1677677812
transform 1 0 924 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2182
timestamp 1677677812
transform 1 0 924 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2183
timestamp 1677677812
transform 1 0 964 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2663
timestamp 1677677812
transform 1 0 964 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2130
timestamp 1677677812
transform 1 0 996 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2131
timestamp 1677677812
transform 1 0 1020 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2469
timestamp 1677677812
transform 1 0 980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2573
timestamp 1677677812
transform 1 0 1004 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2574
timestamp 1677677812
transform 1 0 1060 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2470
timestamp 1677677812
transform 1 0 1108 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2575
timestamp 1677677812
transform 1 0 1132 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2451
timestamp 1677677812
transform 1 0 1212 0 1 3545
box -2 -2 2 2
use M2_M1  M2_M1_2471
timestamp 1677677812
transform 1 0 1204 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2576
timestamp 1677677812
transform 1 0 1196 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2163
timestamp 1677677812
transform 1 0 1212 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2577
timestamp 1677677812
transform 1 0 1236 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2472
timestamp 1677677812
transform 1 0 1260 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2664
timestamp 1677677812
transform 1 0 1284 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2239
timestamp 1677677812
transform 1 0 1284 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2132
timestamp 1677677812
transform 1 0 1308 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2473
timestamp 1677677812
transform 1 0 1308 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2474
timestamp 1677677812
transform 1 0 1316 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2184
timestamp 1677677812
transform 1 0 1316 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2578
timestamp 1677677812
transform 1 0 1324 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2665
timestamp 1677677812
transform 1 0 1316 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2240
timestamp 1677677812
transform 1 0 1316 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2185
timestamp 1677677812
transform 1 0 1332 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2164
timestamp 1677677812
transform 1 0 1372 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2475
timestamp 1677677812
transform 1 0 1388 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2579
timestamp 1677677812
transform 1 0 1372 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2186
timestamp 1677677812
transform 1 0 1380 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2214
timestamp 1677677812
transform 1 0 1372 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2133
timestamp 1677677812
transform 1 0 1428 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2580
timestamp 1677677812
transform 1 0 1444 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2241
timestamp 1677677812
transform 1 0 1444 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2476
timestamp 1677677812
transform 1 0 1516 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2187
timestamp 1677677812
transform 1 0 1516 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2134
timestamp 1677677812
transform 1 0 1548 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2477
timestamp 1677677812
transform 1 0 1548 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2581
timestamp 1677677812
transform 1 0 1540 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2582
timestamp 1677677812
transform 1 0 1556 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2242
timestamp 1677677812
transform 1 0 1540 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2135
timestamp 1677677812
transform 1 0 1628 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2478
timestamp 1677677812
transform 1 0 1604 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2479
timestamp 1677677812
transform 1 0 1612 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2480
timestamp 1677677812
transform 1 0 1628 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2165
timestamp 1677677812
transform 1 0 1636 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2481
timestamp 1677677812
transform 1 0 1644 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2583
timestamp 1677677812
transform 1 0 1636 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2243
timestamp 1677677812
transform 1 0 1612 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2188
timestamp 1677677812
transform 1 0 1644 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2584
timestamp 1677677812
transform 1 0 1652 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2136
timestamp 1677677812
transform 1 0 1660 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2482
timestamp 1677677812
transform 1 0 1724 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2585
timestamp 1677677812
transform 1 0 1716 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2189
timestamp 1677677812
transform 1 0 1748 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2483
timestamp 1677677812
transform 1 0 1764 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2484
timestamp 1677677812
transform 1 0 1780 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2586
timestamp 1677677812
transform 1 0 1756 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2265
timestamp 1677677812
transform 1 0 1756 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2190
timestamp 1677677812
transform 1 0 1780 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2587
timestamp 1677677812
transform 1 0 1788 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2266
timestamp 1677677812
transform 1 0 1780 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2191
timestamp 1677677812
transform 1 0 1804 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2588
timestamp 1677677812
transform 1 0 1812 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2192
timestamp 1677677812
transform 1 0 1820 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2485
timestamp 1677677812
transform 1 0 1836 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2486
timestamp 1677677812
transform 1 0 1852 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2193
timestamp 1677677812
transform 1 0 1844 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2589
timestamp 1677677812
transform 1 0 1852 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2085
timestamp 1677677812
transform 1 0 1964 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2137
timestamp 1677677812
transform 1 0 1892 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2138
timestamp 1677677812
transform 1 0 1972 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2166
timestamp 1677677812
transform 1 0 1924 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2487
timestamp 1677677812
transform 1 0 1972 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2590
timestamp 1677677812
transform 1 0 1892 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2591
timestamp 1677677812
transform 1 0 1940 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2194
timestamp 1677677812
transform 1 0 1972 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2244
timestamp 1677677812
transform 1 0 1924 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2245
timestamp 1677677812
transform 1 0 1940 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2267
timestamp 1677677812
transform 1 0 1932 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2268
timestamp 1677677812
transform 1 0 1956 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2086
timestamp 1677677812
transform 1 0 1988 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2488
timestamp 1677677812
transform 1 0 1988 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2592
timestamp 1677677812
transform 1 0 1988 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2195
timestamp 1677677812
transform 1 0 1996 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2246
timestamp 1677677812
transform 1 0 1988 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2139
timestamp 1677677812
transform 1 0 2028 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2489
timestamp 1677677812
transform 1 0 2044 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2087
timestamp 1677677812
transform 1 0 2156 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2140
timestamp 1677677812
transform 1 0 2148 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2490
timestamp 1677677812
transform 1 0 2148 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2593
timestamp 1677677812
transform 1 0 2060 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2594
timestamp 1677677812
transform 1 0 2068 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2595
timestamp 1677677812
transform 1 0 2100 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2196
timestamp 1677677812
transform 1 0 2148 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2247
timestamp 1677677812
transform 1 0 2060 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2248
timestamp 1677677812
transform 1 0 2100 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2491
timestamp 1677677812
transform 1 0 2164 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2088
timestamp 1677677812
transform 1 0 2204 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2141
timestamp 1677677812
transform 1 0 2212 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2492
timestamp 1677677812
transform 1 0 2204 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2493
timestamp 1677677812
transform 1 0 2212 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2596
timestamp 1677677812
transform 1 0 2180 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2597
timestamp 1677677812
transform 1 0 2196 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2598
timestamp 1677677812
transform 1 0 2236 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2249
timestamp 1677677812
transform 1 0 2228 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2494
timestamp 1677677812
transform 1 0 2252 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2197
timestamp 1677677812
transform 1 0 2252 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2599
timestamp 1677677812
transform 1 0 2292 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2198
timestamp 1677677812
transform 1 0 2324 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2600
timestamp 1677677812
transform 1 0 2332 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2601
timestamp 1677677812
transform 1 0 2340 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2215
timestamp 1677677812
transform 1 0 2292 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2216
timestamp 1677677812
transform 1 0 2340 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2250
timestamp 1677677812
transform 1 0 2244 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2251
timestamp 1677677812
transform 1 0 2332 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2269
timestamp 1677677812
transform 1 0 2276 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2270
timestamp 1677677812
transform 1 0 2324 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2273
timestamp 1677677812
transform 1 0 2284 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2089
timestamp 1677677812
transform 1 0 2372 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2090
timestamp 1677677812
transform 1 0 2420 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2104
timestamp 1677677812
transform 1 0 2412 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2495
timestamp 1677677812
transform 1 0 2356 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2496
timestamp 1677677812
transform 1 0 2364 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2497
timestamp 1677677812
transform 1 0 2388 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2498
timestamp 1677677812
transform 1 0 2420 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2602
timestamp 1677677812
transform 1 0 2356 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2603
timestamp 1677677812
transform 1 0 2372 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2604
timestamp 1677677812
transform 1 0 2388 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2605
timestamp 1677677812
transform 1 0 2396 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2606
timestamp 1677677812
transform 1 0 2412 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2217
timestamp 1677677812
transform 1 0 2388 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2252
timestamp 1677677812
transform 1 0 2364 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2274
timestamp 1677677812
transform 1 0 2356 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2253
timestamp 1677677812
transform 1 0 2404 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2275
timestamp 1677677812
transform 1 0 2412 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2091
timestamp 1677677812
transform 1 0 2468 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2105
timestamp 1677677812
transform 1 0 2452 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2142
timestamp 1677677812
transform 1 0 2436 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2499
timestamp 1677677812
transform 1 0 2436 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2167
timestamp 1677677812
transform 1 0 2444 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2500
timestamp 1677677812
transform 1 0 2460 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2501
timestamp 1677677812
transform 1 0 2476 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2607
timestamp 1677677812
transform 1 0 2444 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2608
timestamp 1677677812
transform 1 0 2452 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2199
timestamp 1677677812
transform 1 0 2460 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2609
timestamp 1677677812
transform 1 0 2468 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2218
timestamp 1677677812
transform 1 0 2452 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2106
timestamp 1677677812
transform 1 0 2508 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2502
timestamp 1677677812
transform 1 0 2524 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2200
timestamp 1677677812
transform 1 0 2524 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2219
timestamp 1677677812
transform 1 0 2516 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2254
timestamp 1677677812
transform 1 0 2508 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2610
timestamp 1677677812
transform 1 0 2548 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2220
timestamp 1677677812
transform 1 0 2548 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2143
timestamp 1677677812
transform 1 0 2572 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2503
timestamp 1677677812
transform 1 0 2564 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2611
timestamp 1677677812
transform 1 0 2572 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2144
timestamp 1677677812
transform 1 0 2604 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2504
timestamp 1677677812
transform 1 0 2604 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2612
timestamp 1677677812
transform 1 0 2620 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2613
timestamp 1677677812
transform 1 0 2636 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2614
timestamp 1677677812
transform 1 0 2644 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2221
timestamp 1677677812
transform 1 0 2636 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2255
timestamp 1677677812
transform 1 0 2644 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2107
timestamp 1677677812
transform 1 0 2668 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2145
timestamp 1677677812
transform 1 0 2676 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2146
timestamp 1677677812
transform 1 0 2692 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2147
timestamp 1677677812
transform 1 0 2708 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2505
timestamp 1677677812
transform 1 0 2668 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2506
timestamp 1677677812
transform 1 0 2676 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2507
timestamp 1677677812
transform 1 0 2700 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2508
timestamp 1677677812
transform 1 0 2708 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2615
timestamp 1677677812
transform 1 0 2692 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2616
timestamp 1677677812
transform 1 0 2708 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2256
timestamp 1677677812
transform 1 0 2676 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2222
timestamp 1677677812
transform 1 0 2708 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2257
timestamp 1677677812
transform 1 0 2708 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2617
timestamp 1677677812
transform 1 0 2740 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2108
timestamp 1677677812
transform 1 0 2756 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2509
timestamp 1677677812
transform 1 0 2756 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2618
timestamp 1677677812
transform 1 0 2788 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2510
timestamp 1677677812
transform 1 0 2860 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2511
timestamp 1677677812
transform 1 0 2876 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2201
timestamp 1677677812
transform 1 0 2868 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2666
timestamp 1677677812
transform 1 0 2868 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2092
timestamp 1677677812
transform 1 0 2892 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2667
timestamp 1677677812
transform 1 0 2884 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2109
timestamp 1677677812
transform 1 0 2908 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2512
timestamp 1677677812
transform 1 0 2908 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2513
timestamp 1677677812
transform 1 0 2916 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2202
timestamp 1677677812
transform 1 0 2916 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2668
timestamp 1677677812
transform 1 0 2916 0 1 3515
box -2 -2 2 2
use M2_M1  M2_M1_2514
timestamp 1677677812
transform 1 0 2972 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2515
timestamp 1677677812
transform 1 0 2980 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2619
timestamp 1677677812
transform 1 0 2948 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2620
timestamp 1677677812
transform 1 0 2964 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2621
timestamp 1677677812
transform 1 0 2988 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2203
timestamp 1677677812
transform 1 0 2996 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2622
timestamp 1677677812
transform 1 0 3004 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2223
timestamp 1677677812
transform 1 0 2972 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2271
timestamp 1677677812
transform 1 0 2988 0 1 3495
box -3 -3 3 3
use M3_M2  M3_M2_2276
timestamp 1677677812
transform 1 0 2972 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2277
timestamp 1677677812
transform 1 0 3004 0 1 3485
box -3 -3 3 3
use M3_M2  M3_M2_2148
timestamp 1677677812
transform 1 0 3028 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2516
timestamp 1677677812
transform 1 0 3028 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2204
timestamp 1677677812
transform 1 0 3020 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2517
timestamp 1677677812
transform 1 0 3060 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2518
timestamp 1677677812
transform 1 0 3076 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2623
timestamp 1677677812
transform 1 0 3052 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2624
timestamp 1677677812
transform 1 0 3068 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2205
timestamp 1677677812
transform 1 0 3076 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2625
timestamp 1677677812
transform 1 0 3084 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2224
timestamp 1677677812
transform 1 0 3068 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2258
timestamp 1677677812
transform 1 0 3052 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2225
timestamp 1677677812
transform 1 0 3084 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2519
timestamp 1677677812
transform 1 0 3108 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2626
timestamp 1677677812
transform 1 0 3124 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2259
timestamp 1677677812
transform 1 0 3124 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2627
timestamp 1677677812
transform 1 0 3140 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2110
timestamp 1677677812
transform 1 0 3156 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2520
timestamp 1677677812
transform 1 0 3164 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2521
timestamp 1677677812
transform 1 0 3180 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2522
timestamp 1677677812
transform 1 0 3196 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2206
timestamp 1677677812
transform 1 0 3156 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2628
timestamp 1677677812
transform 1 0 3188 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2207
timestamp 1677677812
transform 1 0 3196 0 1 3525
box -3 -3 3 3
use M3_M2  M3_M2_2226
timestamp 1677677812
transform 1 0 3188 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2278
timestamp 1677677812
transform 1 0 3164 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2669
timestamp 1677677812
transform 1 0 3204 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2227
timestamp 1677677812
transform 1 0 3212 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2093
timestamp 1677677812
transform 1 0 3252 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2629
timestamp 1677677812
transform 1 0 3260 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2228
timestamp 1677677812
transform 1 0 3260 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2671
timestamp 1677677812
transform 1 0 3252 0 1 3505
box -2 -2 2 2
use M2_M1  M2_M1_2630
timestamp 1677677812
transform 1 0 3324 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2670
timestamp 1677677812
transform 1 0 3324 0 1 3515
box -2 -2 2 2
use M3_M2  M3_M2_2260
timestamp 1677677812
transform 1 0 3324 0 1 3505
box -3 -3 3 3
use M2_M1  M2_M1_2523
timestamp 1677677812
transform 1 0 3340 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2208
timestamp 1677677812
transform 1 0 3340 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2631
timestamp 1677677812
transform 1 0 3348 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2229
timestamp 1677677812
transform 1 0 3348 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2272
timestamp 1677677812
transform 1 0 3348 0 1 3495
box -3 -3 3 3
use M2_M1  M2_M1_2632
timestamp 1677677812
transform 1 0 3388 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2111
timestamp 1677677812
transform 1 0 3412 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2524
timestamp 1677677812
transform 1 0 3412 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2525
timestamp 1677677812
transform 1 0 3428 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2168
timestamp 1677677812
transform 1 0 3468 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2633
timestamp 1677677812
transform 1 0 3468 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2634
timestamp 1677677812
transform 1 0 3516 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2230
timestamp 1677677812
transform 1 0 3516 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2672
timestamp 1677677812
transform 1 0 3516 0 1 3505
box -2 -2 2 2
use M3_M2  M3_M2_2094
timestamp 1677677812
transform 1 0 3548 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2095
timestamp 1677677812
transform 1 0 3572 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2149
timestamp 1677677812
transform 1 0 3564 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2526
timestamp 1677677812
transform 1 0 3532 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2169
timestamp 1677677812
transform 1 0 3540 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2527
timestamp 1677677812
transform 1 0 3548 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2528
timestamp 1677677812
transform 1 0 3564 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2209
timestamp 1677677812
transform 1 0 3532 0 1 3525
box -3 -3 3 3
use M2_M1  M2_M1_2635
timestamp 1677677812
transform 1 0 3540 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2636
timestamp 1677677812
transform 1 0 3556 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2279
timestamp 1677677812
transform 1 0 3564 0 1 3485
box -3 -3 3 3
use M2_M1  M2_M1_2529
timestamp 1677677812
transform 1 0 3604 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2231
timestamp 1677677812
transform 1 0 3604 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2530
timestamp 1677677812
transform 1 0 3628 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2637
timestamp 1677677812
transform 1 0 3620 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2232
timestamp 1677677812
transform 1 0 3620 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2112
timestamp 1677677812
transform 1 0 3700 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2150
timestamp 1677677812
transform 1 0 3724 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2531
timestamp 1677677812
transform 1 0 3708 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2532
timestamp 1677677812
transform 1 0 3724 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2638
timestamp 1677677812
transform 1 0 3700 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2639
timestamp 1677677812
transform 1 0 3716 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2640
timestamp 1677677812
transform 1 0 3756 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2113
timestamp 1677677812
transform 1 0 3780 0 1 3555
box -3 -3 3 3
use M2_M1  M2_M1_2533
timestamp 1677677812
transform 1 0 3772 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2170
timestamp 1677677812
transform 1 0 3780 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2534
timestamp 1677677812
transform 1 0 3788 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2535
timestamp 1677677812
transform 1 0 3796 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2641
timestamp 1677677812
transform 1 0 3780 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2642
timestamp 1677677812
transform 1 0 3796 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2261
timestamp 1677677812
transform 1 0 3780 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2096
timestamp 1677677812
transform 1 0 3828 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2114
timestamp 1677677812
transform 1 0 3820 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2151
timestamp 1677677812
transform 1 0 3820 0 1 3545
box -3 -3 3 3
use M3_M2  M3_M2_2152
timestamp 1677677812
transform 1 0 3836 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2536
timestamp 1677677812
transform 1 0 3820 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2537
timestamp 1677677812
transform 1 0 3836 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2171
timestamp 1677677812
transform 1 0 3844 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2097
timestamp 1677677812
transform 1 0 3860 0 1 3565
box -3 -3 3 3
use M2_M1  M2_M1_2538
timestamp 1677677812
transform 1 0 3852 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2643
timestamp 1677677812
transform 1 0 3828 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2644
timestamp 1677677812
transform 1 0 3844 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2153
timestamp 1677677812
transform 1 0 3924 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2539
timestamp 1677677812
transform 1 0 3900 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2645
timestamp 1677677812
transform 1 0 3924 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2115
timestamp 1677677812
transform 1 0 3996 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2172
timestamp 1677677812
transform 1 0 3996 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2646
timestamp 1677677812
transform 1 0 3996 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2233
timestamp 1677677812
transform 1 0 4028 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2173
timestamp 1677677812
transform 1 0 4052 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2098
timestamp 1677677812
transform 1 0 4068 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2116
timestamp 1677677812
transform 1 0 4092 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2154
timestamp 1677677812
transform 1 0 4164 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2540
timestamp 1677677812
transform 1 0 4092 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2174
timestamp 1677677812
transform 1 0 4116 0 1 3535
box -3 -3 3 3
use M3_M2  M3_M2_2155
timestamp 1677677812
transform 1 0 4204 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2541
timestamp 1677677812
transform 1 0 4188 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2647
timestamp 1677677812
transform 1 0 4116 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2648
timestamp 1677677812
transform 1 0 4172 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2649
timestamp 1677677812
transform 1 0 4228 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2542
timestamp 1677677812
transform 1 0 4292 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2650
timestamp 1677677812
transform 1 0 4284 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2651
timestamp 1677677812
transform 1 0 4292 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2234
timestamp 1677677812
transform 1 0 4292 0 1 3515
box -3 -3 3 3
use M3_M2  M3_M2_2099
timestamp 1677677812
transform 1 0 4348 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2156
timestamp 1677677812
transform 1 0 4332 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2543
timestamp 1677677812
transform 1 0 4332 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2175
timestamp 1677677812
transform 1 0 4340 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2544
timestamp 1677677812
transform 1 0 4348 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2652
timestamp 1677677812
transform 1 0 4324 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2653
timestamp 1677677812
transform 1 0 4340 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2262
timestamp 1677677812
transform 1 0 4340 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2100
timestamp 1677677812
transform 1 0 4380 0 1 3565
box -3 -3 3 3
use M3_M2  M3_M2_2117
timestamp 1677677812
transform 1 0 4380 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2118
timestamp 1677677812
transform 1 0 4396 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2157
timestamp 1677677812
transform 1 0 4428 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2545
timestamp 1677677812
transform 1 0 4380 0 1 3535
box -2 -2 2 2
use M3_M2  M3_M2_2176
timestamp 1677677812
transform 1 0 4404 0 1 3535
box -3 -3 3 3
use M2_M1  M2_M1_2654
timestamp 1677677812
transform 1 0 4404 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2655
timestamp 1677677812
transform 1 0 4460 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2263
timestamp 1677677812
transform 1 0 4372 0 1 3505
box -3 -3 3 3
use M3_M2  M3_M2_2119
timestamp 1677677812
transform 1 0 4500 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2120
timestamp 1677677812
transform 1 0 4532 0 1 3555
box -3 -3 3 3
use M3_M2  M3_M2_2158
timestamp 1677677812
transform 1 0 4516 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2546
timestamp 1677677812
transform 1 0 4500 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2547
timestamp 1677677812
transform 1 0 4516 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2656
timestamp 1677677812
transform 1 0 4508 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2657
timestamp 1677677812
transform 1 0 4524 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2658
timestamp 1677677812
transform 1 0 4532 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2159
timestamp 1677677812
transform 1 0 4596 0 1 3545
box -3 -3 3 3
use M2_M1  M2_M1_2548
timestamp 1677677812
transform 1 0 4572 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2659
timestamp 1677677812
transform 1 0 4596 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2660
timestamp 1677677812
transform 1 0 4652 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2235
timestamp 1677677812
transform 1 0 4684 0 1 3515
box -3 -3 3 3
use M2_M1  M2_M1_2549
timestamp 1677677812
transform 1 0 4700 0 1 3535
box -2 -2 2 2
use M2_M1  M2_M1_2661
timestamp 1677677812
transform 1 0 4724 0 1 3525
box -2 -2 2 2
use M2_M1  M2_M1_2662
timestamp 1677677812
transform 1 0 4780 0 1 3525
box -2 -2 2 2
use M3_M2  M3_M2_2236
timestamp 1677677812
transform 1 0 4724 0 1 3515
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_24
timestamp 1677677812
transform 1 0 24 0 1 3470
box -10 -3 10 3
use FILL  FILL_2220
timestamp 1677677812
transform 1 0 72 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2221
timestamp 1677677812
transform 1 0 80 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2222
timestamp 1677677812
transform 1 0 88 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2223
timestamp 1677677812
transform 1 0 96 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2224
timestamp 1677677812
transform 1 0 104 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2225
timestamp 1677677812
transform 1 0 112 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2226
timestamp 1677677812
transform 1 0 120 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2227
timestamp 1677677812
transform 1 0 128 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_188
timestamp 1677677812
transform -1 0 152 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2228
timestamp 1677677812
transform 1 0 152 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2229
timestamp 1677677812
transform 1 0 160 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2230
timestamp 1677677812
transform 1 0 168 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2238
timestamp 1677677812
transform 1 0 176 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_103
timestamp 1677677812
transform -1 0 224 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2239
timestamp 1677677812
transform 1 0 224 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_161
timestamp 1677677812
transform 1 0 232 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_189
timestamp 1677677812
transform -1 0 344 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2255
timestamp 1677677812
transform 1 0 344 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2257
timestamp 1677677812
transform 1 0 352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2259
timestamp 1677677812
transform 1 0 360 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2261
timestamp 1677677812
transform 1 0 368 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2269
timestamp 1677677812
transform 1 0 376 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_104
timestamp 1677677812
transform -1 0 424 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2270
timestamp 1677677812
transform 1 0 424 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2272
timestamp 1677677812
transform 1 0 432 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2274
timestamp 1677677812
transform 1 0 440 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2276
timestamp 1677677812
transform 1 0 448 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2278
timestamp 1677677812
transform 1 0 456 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2280
timestamp 1677677812
transform 1 0 464 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2282
timestamp 1677677812
transform 1 0 472 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_105
timestamp 1677677812
transform 1 0 480 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2289
timestamp 1677677812
transform 1 0 520 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2291
timestamp 1677677812
transform 1 0 528 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2293
timestamp 1677677812
transform 1 0 536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2295
timestamp 1677677812
transform 1 0 544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2297
timestamp 1677677812
transform 1 0 552 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2298
timestamp 1677677812
transform 1 0 560 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2299
timestamp 1677677812
transform 1 0 568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2301
timestamp 1677677812
transform 1 0 576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2303
timestamp 1677677812
transform 1 0 584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2305
timestamp 1677677812
transform 1 0 592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2312
timestamp 1677677812
transform 1 0 600 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1677677812
transform -1 0 640 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2313
timestamp 1677677812
transform 1 0 640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2315
timestamp 1677677812
transform 1 0 648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2322
timestamp 1677677812
transform 1 0 656 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_1
timestamp 1677677812
transform -1 0 696 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2323
timestamp 1677677812
transform 1 0 696 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2327
timestamp 1677677812
transform 1 0 704 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2328
timestamp 1677677812
transform 1 0 712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2329
timestamp 1677677812
transform 1 0 720 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2330
timestamp 1677677812
transform 1 0 728 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2331
timestamp 1677677812
transform 1 0 736 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2332
timestamp 1677677812
transform 1 0 744 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2333
timestamp 1677677812
transform 1 0 752 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_99
timestamp 1677677812
transform -1 0 800 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2334
timestamp 1677677812
transform 1 0 800 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2335
timestamp 1677677812
transform 1 0 808 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2336
timestamp 1677677812
transform 1 0 816 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2337
timestamp 1677677812
transform 1 0 824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2338
timestamp 1677677812
transform 1 0 832 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_191
timestamp 1677677812
transform -1 0 856 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2339
timestamp 1677677812
transform 1 0 856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2340
timestamp 1677677812
transform 1 0 864 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2341
timestamp 1677677812
transform 1 0 872 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2342
timestamp 1677677812
transform 1 0 880 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_52
timestamp 1677677812
transform 1 0 888 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2343
timestamp 1677677812
transform 1 0 920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2344
timestamp 1677677812
transform 1 0 928 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2345
timestamp 1677677812
transform 1 0 936 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2346
timestamp 1677677812
transform 1 0 944 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2347
timestamp 1677677812
transform 1 0 952 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2349
timestamp 1677677812
transform 1 0 960 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2280
timestamp 1677677812
transform 1 0 1036 0 1 3475
box -3 -3 3 3
use M3_M2  M3_M2_2281
timestamp 1677677812
transform 1 0 1060 0 1 3475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_164
timestamp 1677677812
transform 1 0 968 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2359
timestamp 1677677812
transform 1 0 1064 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2360
timestamp 1677677812
transform 1 0 1072 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2361
timestamp 1677677812
transform 1 0 1080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2362
timestamp 1677677812
transform 1 0 1088 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2282
timestamp 1677677812
transform 1 0 1108 0 1 3475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_165
timestamp 1677677812
transform 1 0 1096 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2370
timestamp 1677677812
transform 1 0 1192 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2371
timestamp 1677677812
transform 1 0 1200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2373
timestamp 1677677812
transform 1 0 1208 0 -1 3570
box -8 -3 16 105
use NOR2X1  NOR2X1_26
timestamp 1677677812
transform 1 0 1216 0 -1 3570
box -8 -3 32 105
use FILL  FILL_2383
timestamp 1677677812
transform 1 0 1240 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2384
timestamp 1677677812
transform 1 0 1248 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2385
timestamp 1677677812
transform 1 0 1256 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2386
timestamp 1677677812
transform 1 0 1264 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2387
timestamp 1677677812
transform 1 0 1272 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_54
timestamp 1677677812
transform -1 0 1312 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2388
timestamp 1677677812
transform 1 0 1312 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2389
timestamp 1677677812
transform 1 0 1320 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2283
timestamp 1677677812
transform 1 0 1340 0 1 3475
box -3 -3 3 3
use FILL  FILL_2390
timestamp 1677677812
transform 1 0 1328 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2391
timestamp 1677677812
transform 1 0 1336 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2397
timestamp 1677677812
transform 1 0 1344 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_55
timestamp 1677677812
transform -1 0 1384 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2398
timestamp 1677677812
transform 1 0 1384 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2399
timestamp 1677677812
transform 1 0 1392 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2400
timestamp 1677677812
transform 1 0 1400 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2401
timestamp 1677677812
transform 1 0 1408 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2402
timestamp 1677677812
transform 1 0 1416 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2403
timestamp 1677677812
transform 1 0 1424 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_194
timestamp 1677677812
transform 1 0 1432 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2404
timestamp 1677677812
transform 1 0 1448 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2405
timestamp 1677677812
transform 1 0 1456 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2406
timestamp 1677677812
transform 1 0 1464 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2407
timestamp 1677677812
transform 1 0 1472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2409
timestamp 1677677812
transform 1 0 1480 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2284
timestamp 1677677812
transform 1 0 1500 0 1 3475
box -3 -3 3 3
use FILL  FILL_2411
timestamp 1677677812
transform 1 0 1488 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2413
timestamp 1677677812
transform 1 0 1496 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2418
timestamp 1677677812
transform 1 0 1504 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2419
timestamp 1677677812
transform 1 0 1512 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2285
timestamp 1677677812
transform 1 0 1532 0 1 3475
box -3 -3 3 3
use FILL  FILL_2420
timestamp 1677677812
transform 1 0 1520 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_101
timestamp 1677677812
transform -1 0 1568 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2421
timestamp 1677677812
transform 1 0 1568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2423
timestamp 1677677812
transform 1 0 1576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2425
timestamp 1677677812
transform 1 0 1584 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2286
timestamp 1677677812
transform 1 0 1604 0 1 3475
box -3 -3 3 3
use FILL  FILL_2427
timestamp 1677677812
transform 1 0 1592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2431
timestamp 1677677812
transform 1 0 1600 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_102
timestamp 1677677812
transform 1 0 1608 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2432
timestamp 1677677812
transform 1 0 1648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2433
timestamp 1677677812
transform 1 0 1656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2434
timestamp 1677677812
transform 1 0 1664 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2435
timestamp 1677677812
transform 1 0 1672 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2436
timestamp 1677677812
transform 1 0 1680 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2437
timestamp 1677677812
transform 1 0 1688 0 -1 3570
box -8 -3 16 105
use AND2X2  AND2X2_2
timestamp 1677677812
transform -1 0 1728 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2438
timestamp 1677677812
transform 1 0 1728 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2439
timestamp 1677677812
transform 1 0 1736 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2440
timestamp 1677677812
transform 1 0 1744 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2442
timestamp 1677677812
transform 1 0 1752 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_103
timestamp 1677677812
transform 1 0 1760 0 -1 3570
box -8 -3 46 105
use M3_M2  M3_M2_2287
timestamp 1677677812
transform 1 0 1812 0 1 3475
box -3 -3 3 3
use FILL  FILL_2446
timestamp 1677677812
transform 1 0 1800 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2448
timestamp 1677677812
transform 1 0 1808 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2459
timestamp 1677677812
transform 1 0 1816 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2460
timestamp 1677677812
transform 1 0 1824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2461
timestamp 1677677812
transform 1 0 1832 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_198
timestamp 1677677812
transform -1 0 1856 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2462
timestamp 1677677812
transform 1 0 1856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2463
timestamp 1677677812
transform 1 0 1864 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2464
timestamp 1677677812
transform 1 0 1872 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2465
timestamp 1677677812
transform 1 0 1880 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_168
timestamp 1677677812
transform -1 0 1984 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2466
timestamp 1677677812
transform 1 0 1984 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_199
timestamp 1677677812
transform 1 0 1992 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2470
timestamp 1677677812
transform 1 0 2008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2472
timestamp 1677677812
transform 1 0 2016 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2494
timestamp 1677677812
transform 1 0 2024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2495
timestamp 1677677812
transform 1 0 2032 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2496
timestamp 1677677812
transform 1 0 2040 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_202
timestamp 1677677812
transform 1 0 2048 0 -1 3570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_171
timestamp 1677677812
transform -1 0 2160 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2497
timestamp 1677677812
transform 1 0 2160 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2498
timestamp 1677677812
transform 1 0 2168 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_113
timestamp 1677677812
transform -1 0 2216 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2499
timestamp 1677677812
transform 1 0 2216 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2500
timestamp 1677677812
transform 1 0 2224 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2501
timestamp 1677677812
transform 1 0 2232 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_172
timestamp 1677677812
transform 1 0 2240 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_203
timestamp 1677677812
transform -1 0 2352 0 -1 3570
box -9 -3 26 105
use AOI22X1  AOI22X1_114
timestamp 1677677812
transform -1 0 2392 0 -1 3570
box -8 -3 46 105
use M3_M2  M3_M2_2288
timestamp 1677677812
transform 1 0 2420 0 1 3475
box -3 -3 3 3
use AND2X2  AND2X2_3
timestamp 1677677812
transform -1 0 2424 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2502
timestamp 1677677812
transform 1 0 2424 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_204
timestamp 1677677812
transform 1 0 2432 0 -1 3570
box -9 -3 26 105
use AOI22X1  AOI22X1_115
timestamp 1677677812
transform 1 0 2448 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2503
timestamp 1677677812
transform 1 0 2488 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2504
timestamp 1677677812
transform 1 0 2496 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2505
timestamp 1677677812
transform 1 0 2504 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2506
timestamp 1677677812
transform 1 0 2512 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2507
timestamp 1677677812
transform 1 0 2520 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2508
timestamp 1677677812
transform 1 0 2528 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2509
timestamp 1677677812
transform 1 0 2536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2510
timestamp 1677677812
transform 1 0 2544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2511
timestamp 1677677812
transform 1 0 2552 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2512
timestamp 1677677812
transform 1 0 2560 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2514
timestamp 1677677812
transform 1 0 2568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2517
timestamp 1677677812
transform 1 0 2576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2518
timestamp 1677677812
transform 1 0 2584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2519
timestamp 1677677812
transform 1 0 2592 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_116
timestamp 1677677812
transform 1 0 2600 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2520
timestamp 1677677812
transform 1 0 2640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2521
timestamp 1677677812
transform 1 0 2648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2522
timestamp 1677677812
transform 1 0 2656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2523
timestamp 1677677812
transform 1 0 2664 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_117
timestamp 1677677812
transform 1 0 2672 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2524
timestamp 1677677812
transform 1 0 2712 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2525
timestamp 1677677812
transform 1 0 2720 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_205
timestamp 1677677812
transform 1 0 2728 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2526
timestamp 1677677812
transform 1 0 2744 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2527
timestamp 1677677812
transform 1 0 2752 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2528
timestamp 1677677812
transform 1 0 2760 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2529
timestamp 1677677812
transform 1 0 2768 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2530
timestamp 1677677812
transform 1 0 2776 0 -1 3570
box -8 -3 16 105
use OAI21X1  OAI21X1_58
timestamp 1677677812
transform 1 0 2784 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2532
timestamp 1677677812
transform 1 0 2816 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2534
timestamp 1677677812
transform 1 0 2824 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2536
timestamp 1677677812
transform 1 0 2832 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2537
timestamp 1677677812
transform 1 0 2840 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2538
timestamp 1677677812
transform 1 0 2848 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2539
timestamp 1677677812
transform 1 0 2856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2541
timestamp 1677677812
transform 1 0 2864 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2550
timestamp 1677677812
transform 1 0 2872 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2289
timestamp 1677677812
transform 1 0 2892 0 1 3475
box -3 -3 3 3
use OAI21X1  OAI21X1_60
timestamp 1677677812
transform -1 0 2912 0 -1 3570
box -8 -3 34 105
use FILL  FILL_2551
timestamp 1677677812
transform 1 0 2912 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2552
timestamp 1677677812
transform 1 0 2920 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2553
timestamp 1677677812
transform 1 0 2928 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2554
timestamp 1677677812
transform 1 0 2936 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2290
timestamp 1677677812
transform 1 0 2980 0 1 3475
box -3 -3 3 3
use OAI21X1  OAI21X1_61
timestamp 1677677812
transform -1 0 2976 0 -1 3570
box -8 -3 34 105
use M3_M2  M3_M2_2291
timestamp 1677677812
transform 1 0 2996 0 1 3475
box -3 -3 3 3
use AND2X2  AND2X2_4
timestamp 1677677812
transform 1 0 2976 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2555
timestamp 1677677812
transform 1 0 3008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2556
timestamp 1677677812
transform 1 0 3016 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2557
timestamp 1677677812
transform 1 0 3024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2558
timestamp 1677677812
transform 1 0 3032 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_105
timestamp 1677677812
transform 1 0 3040 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2559
timestamp 1677677812
transform 1 0 3080 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2561
timestamp 1677677812
transform 1 0 3088 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2563
timestamp 1677677812
transform 1 0 3096 0 -1 3570
box -8 -3 16 105
use INVX2  INVX2_206
timestamp 1677677812
transform 1 0 3104 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2566
timestamp 1677677812
transform 1 0 3120 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2567
timestamp 1677677812
transform 1 0 3128 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2568
timestamp 1677677812
transform 1 0 3136 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2569
timestamp 1677677812
transform 1 0 3144 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2570
timestamp 1677677812
transform 1 0 3152 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_107
timestamp 1677677812
transform 1 0 3160 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2577
timestamp 1677677812
transform 1 0 3200 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2578
timestamp 1677677812
transform 1 0 3208 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2579
timestamp 1677677812
transform 1 0 3216 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2581
timestamp 1677677812
transform 1 0 3224 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2588
timestamp 1677677812
transform 1 0 3232 0 -1 3570
box -8 -3 16 105
use NAND3X1  NAND3X1_12
timestamp 1677677812
transform -1 0 3272 0 -1 3570
box -8 -3 40 105
use FILL  FILL_2589
timestamp 1677677812
transform 1 0 3272 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2590
timestamp 1677677812
transform 1 0 3280 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2591
timestamp 1677677812
transform 1 0 3288 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2592
timestamp 1677677812
transform 1 0 3296 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2593
timestamp 1677677812
transform 1 0 3304 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2595
timestamp 1677677812
transform 1 0 3312 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2597
timestamp 1677677812
transform 1 0 3320 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_119
timestamp 1677677812
transform 1 0 3328 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2602
timestamp 1677677812
transform 1 0 3368 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2603
timestamp 1677677812
transform 1 0 3376 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2604
timestamp 1677677812
transform 1 0 3384 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2605
timestamp 1677677812
transform 1 0 3392 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2607
timestamp 1677677812
transform 1 0 3400 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2609
timestamp 1677677812
transform 1 0 3408 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_176
timestamp 1677677812
transform 1 0 3416 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2618
timestamp 1677677812
transform 1 0 3512 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2624
timestamp 1677677812
transform 1 0 3520 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_109
timestamp 1677677812
transform -1 0 3568 0 -1 3570
box -8 -3 46 105
use M3_M2  M3_M2_2292
timestamp 1677677812
transform 1 0 3580 0 1 3475
box -3 -3 3 3
use FILL  FILL_2625
timestamp 1677677812
transform 1 0 3568 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2627
timestamp 1677677812
transform 1 0 3576 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2629
timestamp 1677677812
transform 1 0 3584 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2631
timestamp 1677677812
transform 1 0 3592 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2633
timestamp 1677677812
transform 1 0 3600 0 -1 3570
box -8 -3 16 105
use M3_M2  M3_M2_2293
timestamp 1677677812
transform 1 0 3628 0 1 3475
box -3 -3 3 3
use INVX2  INVX2_209
timestamp 1677677812
transform 1 0 3608 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2637
timestamp 1677677812
transform 1 0 3624 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2639
timestamp 1677677812
transform 1 0 3632 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2641
timestamp 1677677812
transform 1 0 3640 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2642
timestamp 1677677812
transform 1 0 3648 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2643
timestamp 1677677812
transform 1 0 3656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2644
timestamp 1677677812
transform 1 0 3664 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2645
timestamp 1677677812
transform 1 0 3672 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2646
timestamp 1677677812
transform 1 0 3680 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_110
timestamp 1677677812
transform -1 0 3728 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2647
timestamp 1677677812
transform 1 0 3728 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2648
timestamp 1677677812
transform 1 0 3736 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2650
timestamp 1677677812
transform 1 0 3744 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2653
timestamp 1677677812
transform 1 0 3752 0 -1 3570
box -8 -3 16 105
use AOI22X1  AOI22X1_121
timestamp 1677677812
transform 1 0 3760 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2654
timestamp 1677677812
transform 1 0 3800 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2656
timestamp 1677677812
transform 1 0 3808 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_111
timestamp 1677677812
transform 1 0 3816 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2663
timestamp 1677677812
transform 1 0 3856 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2665
timestamp 1677677812
transform 1 0 3864 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2667
timestamp 1677677812
transform 1 0 3872 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2669
timestamp 1677677812
transform 1 0 3880 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_178
timestamp 1677677812
transform 1 0 3888 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_211
timestamp 1677677812
transform 1 0 3984 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2678
timestamp 1677677812
transform 1 0 4000 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2680
timestamp 1677677812
transform 1 0 4008 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2682
timestamp 1677677812
transform 1 0 4016 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2684
timestamp 1677677812
transform 1 0 4024 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2697
timestamp 1677677812
transform 1 0 4032 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2698
timestamp 1677677812
transform 1 0 4040 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2699
timestamp 1677677812
transform 1 0 4048 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2700
timestamp 1677677812
transform 1 0 4056 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2701
timestamp 1677677812
transform 1 0 4064 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2702
timestamp 1677677812
transform 1 0 4072 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_181
timestamp 1677677812
transform 1 0 4080 0 -1 3570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_182
timestamp 1677677812
transform 1 0 4176 0 -1 3570
box -8 -3 104 105
use INVX2  INVX2_213
timestamp 1677677812
transform 1 0 4272 0 -1 3570
box -9 -3 26 105
use FILL  FILL_2703
timestamp 1677677812
transform 1 0 4288 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2704
timestamp 1677677812
transform 1 0 4296 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2705
timestamp 1677677812
transform 1 0 4304 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_115
timestamp 1677677812
transform 1 0 4312 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2706
timestamp 1677677812
transform 1 0 4352 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2707
timestamp 1677677812
transform 1 0 4360 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_183
timestamp 1677677812
transform 1 0 4368 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2708
timestamp 1677677812
transform 1 0 4464 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2709
timestamp 1677677812
transform 1 0 4472 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2710
timestamp 1677677812
transform 1 0 4480 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2713
timestamp 1677677812
transform 1 0 4488 0 -1 3570
box -8 -3 16 105
use OAI22X1  OAI22X1_117
timestamp 1677677812
transform -1 0 4536 0 -1 3570
box -8 -3 46 105
use FILL  FILL_2714
timestamp 1677677812
transform 1 0 4536 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2716
timestamp 1677677812
transform 1 0 4544 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2718
timestamp 1677677812
transform 1 0 4552 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_184
timestamp 1677677812
transform 1 0 4560 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2734
timestamp 1677677812
transform 1 0 4656 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2735
timestamp 1677677812
transform 1 0 4664 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2736
timestamp 1677677812
transform 1 0 4672 0 -1 3570
box -8 -3 16 105
use FILL  FILL_2737
timestamp 1677677812
transform 1 0 4680 0 -1 3570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_185
timestamp 1677677812
transform 1 0 4688 0 -1 3570
box -8 -3 104 105
use FILL  FILL_2738
timestamp 1677677812
transform 1 0 4784 0 -1 3570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_25
timestamp 1677677812
transform 1 0 4843 0 1 3470
box -10 -3 10 3
use M3_M2  M3_M2_2338
timestamp 1677677812
transform 1 0 92 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2679
timestamp 1677677812
transform 1 0 124 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2780
timestamp 1677677812
transform 1 0 92 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2781
timestamp 1677677812
transform 1 0 180 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2680
timestamp 1677677812
transform 1 0 196 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2412
timestamp 1677677812
transform 1 0 196 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2339
timestamp 1677677812
transform 1 0 244 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2681
timestamp 1677677812
transform 1 0 228 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2682
timestamp 1677677812
transform 1 0 244 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2782
timestamp 1677677812
transform 1 0 236 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2783
timestamp 1677677812
transform 1 0 252 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2413
timestamp 1677677812
transform 1 0 252 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2434
timestamp 1677677812
transform 1 0 236 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2294
timestamp 1677677812
transform 1 0 292 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2295
timestamp 1677677812
transform 1 0 324 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2340
timestamp 1677677812
transform 1 0 340 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2341
timestamp 1677677812
transform 1 0 380 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2683
timestamp 1677677812
transform 1 0 340 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2684
timestamp 1677677812
transform 1 0 372 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2685
timestamp 1677677812
transform 1 0 380 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2784
timestamp 1677677812
transform 1 0 292 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2414
timestamp 1677677812
transform 1 0 292 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2373
timestamp 1677677812
transform 1 0 404 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2785
timestamp 1677677812
transform 1 0 396 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2415
timestamp 1677677812
transform 1 0 388 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2786
timestamp 1677677812
transform 1 0 412 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2862
timestamp 1677677812
transform 1 0 412 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_2391
timestamp 1677677812
transform 1 0 428 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2863
timestamp 1677677812
transform 1 0 436 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_2313
timestamp 1677677812
transform 1 0 452 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2342
timestamp 1677677812
transform 1 0 476 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2686
timestamp 1677677812
transform 1 0 452 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2687
timestamp 1677677812
transform 1 0 476 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2392
timestamp 1677677812
transform 1 0 452 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2787
timestamp 1677677812
transform 1 0 460 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2393
timestamp 1677677812
transform 1 0 468 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2688
timestamp 1677677812
transform 1 0 492 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2788
timestamp 1677677812
transform 1 0 492 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2330
timestamp 1677677812
transform 1 0 532 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2343
timestamp 1677677812
transform 1 0 524 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2689
timestamp 1677677812
transform 1 0 532 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2314
timestamp 1677677812
transform 1 0 580 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2331
timestamp 1677677812
transform 1 0 580 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2690
timestamp 1677677812
transform 1 0 580 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2691
timestamp 1677677812
transform 1 0 644 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2692
timestamp 1677677812
transform 1 0 652 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2789
timestamp 1677677812
transform 1 0 556 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2302
timestamp 1677677812
transform 1 0 684 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2344
timestamp 1677677812
transform 1 0 684 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2790
timestamp 1677677812
transform 1 0 684 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2791
timestamp 1677677812
transform 1 0 692 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2864
timestamp 1677677812
transform 1 0 676 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_2435
timestamp 1677677812
transform 1 0 668 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2315
timestamp 1677677812
transform 1 0 708 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2303
timestamp 1677677812
transform 1 0 732 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2332
timestamp 1677677812
transform 1 0 724 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2345
timestamp 1677677812
transform 1 0 716 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2693
timestamp 1677677812
transform 1 0 740 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2436
timestamp 1677677812
transform 1 0 732 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2316
timestamp 1677677812
transform 1 0 796 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2333
timestamp 1677677812
transform 1 0 772 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2694
timestamp 1677677812
transform 1 0 812 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2792
timestamp 1677677812
transform 1 0 780 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2394
timestamp 1677677812
transform 1 0 876 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2865
timestamp 1677677812
transform 1 0 876 0 1 3395
box -2 -2 2 2
use M2_M1  M2_M1_2695
timestamp 1677677812
transform 1 0 908 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2793
timestamp 1677677812
transform 1 0 980 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2304
timestamp 1677677812
transform 1 0 1028 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2696
timestamp 1677677812
transform 1 0 1028 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2395
timestamp 1677677812
transform 1 0 1028 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2794
timestamp 1677677812
transform 1 0 1036 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2334
timestamp 1677677812
transform 1 0 1060 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2697
timestamp 1677677812
transform 1 0 1060 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2396
timestamp 1677677812
transform 1 0 1068 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2296
timestamp 1677677812
transform 1 0 1084 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_2795
timestamp 1677677812
transform 1 0 1076 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2796
timestamp 1677677812
transform 1 0 1084 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2297
timestamp 1677677812
transform 1 0 1108 0 1 3465
box -3 -3 3 3
use M2_M1  M2_M1_2673
timestamp 1677677812
transform 1 0 1124 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2374
timestamp 1677677812
transform 1 0 1124 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2317
timestamp 1677677812
transform 1 0 1156 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2335
timestamp 1677677812
transform 1 0 1148 0 1 3435
box -3 -3 3 3
use M2_M1  M2_M1_2698
timestamp 1677677812
transform 1 0 1132 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2699
timestamp 1677677812
transform 1 0 1148 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2700
timestamp 1677677812
transform 1 0 1172 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2797
timestamp 1677677812
transform 1 0 1156 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2798
timestamp 1677677812
transform 1 0 1164 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2336
timestamp 1677677812
transform 1 0 1196 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2416
timestamp 1677677812
transform 1 0 1188 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2305
timestamp 1677677812
transform 1 0 1212 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2318
timestamp 1677677812
transform 1 0 1228 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2346
timestamp 1677677812
transform 1 0 1236 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2319
timestamp 1677677812
transform 1 0 1252 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2347
timestamp 1677677812
transform 1 0 1276 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2701
timestamp 1677677812
transform 1 0 1236 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2702
timestamp 1677677812
transform 1 0 1244 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2417
timestamp 1677677812
transform 1 0 1236 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2375
timestamp 1677677812
transform 1 0 1260 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2703
timestamp 1677677812
transform 1 0 1276 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2799
timestamp 1677677812
transform 1 0 1324 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2800
timestamp 1677677812
transform 1 0 1340 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2376
timestamp 1677677812
transform 1 0 1380 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2704
timestamp 1677677812
transform 1 0 1388 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2705
timestamp 1677677812
transform 1 0 1452 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2801
timestamp 1677677812
transform 1 0 1404 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2418
timestamp 1677677812
transform 1 0 1404 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2706
timestamp 1677677812
transform 1 0 1500 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2707
timestamp 1677677812
transform 1 0 1516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2708
timestamp 1677677812
transform 1 0 1564 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2802
timestamp 1677677812
transform 1 0 1596 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2419
timestamp 1677677812
transform 1 0 1596 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2298
timestamp 1677677812
transform 1 0 1620 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2348
timestamp 1677677812
transform 1 0 1636 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2420
timestamp 1677677812
transform 1 0 1628 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2397
timestamp 1677677812
transform 1 0 1644 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2320
timestamp 1677677812
transform 1 0 1708 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2709
timestamp 1677677812
transform 1 0 1684 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2803
timestamp 1677677812
transform 1 0 1660 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2398
timestamp 1677677812
transform 1 0 1684 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2399
timestamp 1677677812
transform 1 0 1700 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2400
timestamp 1677677812
transform 1 0 1724 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2421
timestamp 1677677812
transform 1 0 1660 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2349
timestamp 1677677812
transform 1 0 1756 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2710
timestamp 1677677812
transform 1 0 1748 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2711
timestamp 1677677812
transform 1 0 1756 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2321
timestamp 1677677812
transform 1 0 1772 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2712
timestamp 1677677812
transform 1 0 1772 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2804
timestamp 1677677812
transform 1 0 1764 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2322
timestamp 1677677812
transform 1 0 1788 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2713
timestamp 1677677812
transform 1 0 1796 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2805
timestamp 1677677812
transform 1 0 1788 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2714
timestamp 1677677812
transform 1 0 1844 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2806
timestamp 1677677812
transform 1 0 1892 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2422
timestamp 1677677812
transform 1 0 1892 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2306
timestamp 1677677812
transform 1 0 1948 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2307
timestamp 1677677812
transform 1 0 1964 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2350
timestamp 1677677812
transform 1 0 1972 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2377
timestamp 1677677812
transform 1 0 1948 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2351
timestamp 1677677812
transform 1 0 2012 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2715
timestamp 1677677812
transform 1 0 1972 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2716
timestamp 1677677812
transform 1 0 2004 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2717
timestamp 1677677812
transform 1 0 2012 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2807
timestamp 1677677812
transform 1 0 1924 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2423
timestamp 1677677812
transform 1 0 1924 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2424
timestamp 1677677812
transform 1 0 1972 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2808
timestamp 1677677812
transform 1 0 2052 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2425
timestamp 1677677812
transform 1 0 2052 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2352
timestamp 1677677812
transform 1 0 2116 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2353
timestamp 1677677812
transform 1 0 2156 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2718
timestamp 1677677812
transform 1 0 2116 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2719
timestamp 1677677812
transform 1 0 2148 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2720
timestamp 1677677812
transform 1 0 2156 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2809
timestamp 1677677812
transform 1 0 2068 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2426
timestamp 1677677812
transform 1 0 2100 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2810
timestamp 1677677812
transform 1 0 2172 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2427
timestamp 1677677812
transform 1 0 2180 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2354
timestamp 1677677812
transform 1 0 2196 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2721
timestamp 1677677812
transform 1 0 2204 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2722
timestamp 1677677812
transform 1 0 2260 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2811
timestamp 1677677812
transform 1 0 2284 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2428
timestamp 1677677812
transform 1 0 2212 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2723
timestamp 1677677812
transform 1 0 2308 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2724
timestamp 1677677812
transform 1 0 2324 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2725
timestamp 1677677812
transform 1 0 2356 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2812
timestamp 1677677812
transform 1 0 2332 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2813
timestamp 1677677812
transform 1 0 2348 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2814
timestamp 1677677812
transform 1 0 2364 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2429
timestamp 1677677812
transform 1 0 2348 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2726
timestamp 1677677812
transform 1 0 2380 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2323
timestamp 1677677812
transform 1 0 2404 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2727
timestamp 1677677812
transform 1 0 2404 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2437
timestamp 1677677812
transform 1 0 2404 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2815
timestamp 1677677812
transform 1 0 2420 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2866
timestamp 1677677812
transform 1 0 2428 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_2308
timestamp 1677677812
transform 1 0 2452 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2816
timestamp 1677677812
transform 1 0 2452 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2355
timestamp 1677677812
transform 1 0 2492 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2356
timestamp 1677677812
transform 1 0 2508 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2728
timestamp 1677677812
transform 1 0 2508 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2729
timestamp 1677677812
transform 1 0 2516 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2730
timestamp 1677677812
transform 1 0 2532 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2817
timestamp 1677677812
transform 1 0 2508 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2818
timestamp 1677677812
transform 1 0 2516 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2430
timestamp 1677677812
transform 1 0 2508 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2357
timestamp 1677677812
transform 1 0 2556 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2819
timestamp 1677677812
transform 1 0 2556 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2358
timestamp 1677677812
transform 1 0 2572 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2731
timestamp 1677677812
transform 1 0 2564 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2820
timestamp 1677677812
transform 1 0 2572 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2732
timestamp 1677677812
transform 1 0 2596 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2674
timestamp 1677677812
transform 1 0 2612 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2359
timestamp 1677677812
transform 1 0 2692 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2733
timestamp 1677677812
transform 1 0 2676 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2734
timestamp 1677677812
transform 1 0 2692 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2821
timestamp 1677677812
transform 1 0 2660 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2378
timestamp 1677677812
transform 1 0 2700 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2735
timestamp 1677677812
transform 1 0 2708 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2822
timestamp 1677677812
transform 1 0 2708 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2360
timestamp 1677677812
transform 1 0 2732 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2736
timestamp 1677677812
transform 1 0 2732 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2867
timestamp 1677677812
transform 1 0 2748 0 1 3395
box -2 -2 2 2
use M3_M2  M3_M2_2438
timestamp 1677677812
transform 1 0 2748 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2675
timestamp 1677677812
transform 1 0 2812 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2379
timestamp 1677677812
transform 1 0 2804 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2823
timestamp 1677677812
transform 1 0 2788 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2824
timestamp 1677677812
transform 1 0 2796 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2825
timestamp 1677677812
transform 1 0 2804 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2439
timestamp 1677677812
transform 1 0 2788 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2380
timestamp 1677677812
transform 1 0 2828 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2440
timestamp 1677677812
transform 1 0 2828 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2676
timestamp 1677677812
transform 1 0 2844 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2737
timestamp 1677677812
transform 1 0 2844 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2441
timestamp 1677677812
transform 1 0 2844 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2677
timestamp 1677677812
transform 1 0 2884 0 1 3425
box -2 -2 2 2
use M3_M2  M3_M2_2381
timestamp 1677677812
transform 1 0 2876 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2826
timestamp 1677677812
transform 1 0 2884 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2442
timestamp 1677677812
transform 1 0 2884 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2309
timestamp 1677677812
transform 1 0 2900 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2827
timestamp 1677677812
transform 1 0 2892 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2310
timestamp 1677677812
transform 1 0 2948 0 1 3455
box -3 -3 3 3
use M3_M2  M3_M2_2361
timestamp 1677677812
transform 1 0 2948 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2738
timestamp 1677677812
transform 1 0 2948 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2324
timestamp 1677677812
transform 1 0 2972 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2739
timestamp 1677677812
transform 1 0 2996 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2401
timestamp 1677677812
transform 1 0 2988 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2311
timestamp 1677677812
transform 1 0 3084 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2740
timestamp 1677677812
transform 1 0 3044 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2828
timestamp 1677677812
transform 1 0 3020 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2741
timestamp 1677677812
transform 1 0 3108 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2443
timestamp 1677677812
transform 1 0 3068 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2444
timestamp 1677677812
transform 1 0 3100 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2742
timestamp 1677677812
transform 1 0 3164 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2743
timestamp 1677677812
transform 1 0 3220 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2829
timestamp 1677677812
transform 1 0 3140 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2445
timestamp 1677677812
transform 1 0 3140 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2446
timestamp 1677677812
transform 1 0 3228 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2299
timestamp 1677677812
transform 1 0 3268 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2312
timestamp 1677677812
transform 1 0 3300 0 1 3455
box -3 -3 3 3
use M2_M1  M2_M1_2744
timestamp 1677677812
transform 1 0 3284 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2745
timestamp 1677677812
transform 1 0 3324 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2830
timestamp 1677677812
transform 1 0 3244 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2447
timestamp 1677677812
transform 1 0 3244 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2382
timestamp 1677677812
transform 1 0 3340 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2362
timestamp 1677677812
transform 1 0 3364 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2746
timestamp 1677677812
transform 1 0 3348 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2747
timestamp 1677677812
transform 1 0 3364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2831
timestamp 1677677812
transform 1 0 3340 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2448
timestamp 1677677812
transform 1 0 3340 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2300
timestamp 1677677812
transform 1 0 3404 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2301
timestamp 1677677812
transform 1 0 3436 0 1 3465
box -3 -3 3 3
use M3_M2  M3_M2_2337
timestamp 1677677812
transform 1 0 3476 0 1 3435
box -3 -3 3 3
use M3_M2  M3_M2_2363
timestamp 1677677812
transform 1 0 3492 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2748
timestamp 1677677812
transform 1 0 3460 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2832
timestamp 1677677812
transform 1 0 3412 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2402
timestamp 1677677812
transform 1 0 3460 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2749
timestamp 1677677812
transform 1 0 3500 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2383
timestamp 1677677812
transform 1 0 3516 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2833
timestamp 1677677812
transform 1 0 3516 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2364
timestamp 1677677812
transform 1 0 3540 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2750
timestamp 1677677812
transform 1 0 3540 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2751
timestamp 1677677812
transform 1 0 3556 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2384
timestamp 1677677812
transform 1 0 3564 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2403
timestamp 1677677812
transform 1 0 3540 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2834
timestamp 1677677812
transform 1 0 3548 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2835
timestamp 1677677812
transform 1 0 3564 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2836
timestamp 1677677812
transform 1 0 3580 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2752
timestamp 1677677812
transform 1 0 3660 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2385
timestamp 1677677812
transform 1 0 3684 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2837
timestamp 1677677812
transform 1 0 3668 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2838
timestamp 1677677812
transform 1 0 3684 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2839
timestamp 1677677812
transform 1 0 3692 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2449
timestamp 1677677812
transform 1 0 3684 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2753
timestamp 1677677812
transform 1 0 3708 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2325
timestamp 1677677812
transform 1 0 3724 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2754
timestamp 1677677812
transform 1 0 3724 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2365
timestamp 1677677812
transform 1 0 3780 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2386
timestamp 1677677812
transform 1 0 3772 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2755
timestamp 1677677812
transform 1 0 3780 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2840
timestamp 1677677812
transform 1 0 3772 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2756
timestamp 1677677812
transform 1 0 3828 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2366
timestamp 1677677812
transform 1 0 3852 0 1 3425
box -3 -3 3 3
use M3_M2  M3_M2_2367
timestamp 1677677812
transform 1 0 3868 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2678
timestamp 1677677812
transform 1 0 3876 0 1 3425
box -2 -2 2 2
use M2_M1  M2_M1_2757
timestamp 1677677812
transform 1 0 3860 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2841
timestamp 1677677812
transform 1 0 3852 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2404
timestamp 1677677812
transform 1 0 3860 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2368
timestamp 1677677812
transform 1 0 3884 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2842
timestamp 1677677812
transform 1 0 3892 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2450
timestamp 1677677812
transform 1 0 3892 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2326
timestamp 1677677812
transform 1 0 3940 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2327
timestamp 1677677812
transform 1 0 3972 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2758
timestamp 1677677812
transform 1 0 3932 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2759
timestamp 1677677812
transform 1 0 3988 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2387
timestamp 1677677812
transform 1 0 3996 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2843
timestamp 1677677812
transform 1 0 3908 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2405
timestamp 1677677812
transform 1 0 3932 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2406
timestamp 1677677812
transform 1 0 3948 0 1 3405
box -3 -3 3 3
use M3_M2  M3_M2_2407
timestamp 1677677812
transform 1 0 3988 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2844
timestamp 1677677812
transform 1 0 3996 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2369
timestamp 1677677812
transform 1 0 4044 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2760
timestamp 1677677812
transform 1 0 4028 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2761
timestamp 1677677812
transform 1 0 4044 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2845
timestamp 1677677812
transform 1 0 4036 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2408
timestamp 1677677812
transform 1 0 4044 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2846
timestamp 1677677812
transform 1 0 4052 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2370
timestamp 1677677812
transform 1 0 4180 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2762
timestamp 1677677812
transform 1 0 4124 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2847
timestamp 1677677812
transform 1 0 4100 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2409
timestamp 1677677812
transform 1 0 4124 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2763
timestamp 1677677812
transform 1 0 4188 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2848
timestamp 1677677812
transform 1 0 4196 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2328
timestamp 1677677812
transform 1 0 4220 0 1 3445
box -3 -3 3 3
use M3_M2  M3_M2_2329
timestamp 1677677812
transform 1 0 4236 0 1 3445
box -3 -3 3 3
use M2_M1  M2_M1_2764
timestamp 1677677812
transform 1 0 4220 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2765
timestamp 1677677812
transform 1 0 4236 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2388
timestamp 1677677812
transform 1 0 4244 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2849
timestamp 1677677812
transform 1 0 4228 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2850
timestamp 1677677812
transform 1 0 4244 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2451
timestamp 1677677812
transform 1 0 4244 0 1 3385
box -3 -3 3 3
use M3_M2  M3_M2_2389
timestamp 1677677812
transform 1 0 4284 0 1 3415
box -3 -3 3 3
use M2_M1  M2_M1_2851
timestamp 1677677812
transform 1 0 4300 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2766
timestamp 1677677812
transform 1 0 4316 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2390
timestamp 1677677812
transform 1 0 4324 0 1 3415
box -3 -3 3 3
use M3_M2  M3_M2_2410
timestamp 1677677812
transform 1 0 4316 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2852
timestamp 1677677812
transform 1 0 4324 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2431
timestamp 1677677812
transform 1 0 4332 0 1 3395
box -3 -3 3 3
use M2_M1  M2_M1_2767
timestamp 1677677812
transform 1 0 4348 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2768
timestamp 1677677812
transform 1 0 4364 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2769
timestamp 1677677812
transform 1 0 4380 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2853
timestamp 1677677812
transform 1 0 4372 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2411
timestamp 1677677812
transform 1 0 4380 0 1 3405
box -3 -3 3 3
use M2_M1  M2_M1_2770
timestamp 1677677812
transform 1 0 4452 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2771
timestamp 1677677812
transform 1 0 4476 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2772
timestamp 1677677812
transform 1 0 4492 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2854
timestamp 1677677812
transform 1 0 4460 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2855
timestamp 1677677812
transform 1 0 4468 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2432
timestamp 1677677812
transform 1 0 4468 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2371
timestamp 1677677812
transform 1 0 4508 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2773
timestamp 1677677812
transform 1 0 4508 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2372
timestamp 1677677812
transform 1 0 4644 0 1 3425
box -3 -3 3 3
use M2_M1  M2_M1_2774
timestamp 1677677812
transform 1 0 4580 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2775
timestamp 1677677812
transform 1 0 4636 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2776
timestamp 1677677812
transform 1 0 4644 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2856
timestamp 1677677812
transform 1 0 4556 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2452
timestamp 1677677812
transform 1 0 4556 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2777
timestamp 1677677812
transform 1 0 4660 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2857
timestamp 1677677812
transform 1 0 4652 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2858
timestamp 1677677812
transform 1 0 4660 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2778
timestamp 1677677812
transform 1 0 4692 0 1 3415
box -2 -2 2 2
use M2_M1  M2_M1_2859
timestamp 1677677812
transform 1 0 4684 0 1 3405
box -2 -2 2 2
use M3_M2  M3_M2_2433
timestamp 1677677812
transform 1 0 4692 0 1 3395
box -3 -3 3 3
use M3_M2  M3_M2_2453
timestamp 1677677812
transform 1 0 4676 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2779
timestamp 1677677812
transform 1 0 4708 0 1 3415
box -2 -2 2 2
use M3_M2  M3_M2_2454
timestamp 1677677812
transform 1 0 4708 0 1 3385
box -3 -3 3 3
use M2_M1  M2_M1_2860
timestamp 1677677812
transform 1 0 4740 0 1 3405
box -2 -2 2 2
use M2_M1  M2_M1_2861
timestamp 1677677812
transform 1 0 4780 0 1 3405
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_26
timestamp 1677677812
transform 1 0 48 0 1 3370
box -10 -3 10 3
use FILL  FILL_2739
timestamp 1677677812
transform 1 0 72 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_186
timestamp 1677677812
transform 1 0 80 0 1 3370
box -8 -3 104 105
use FILL  FILL_2741
timestamp 1677677812
transform 1 0 176 0 1 3370
box -8 -3 16 105
use FILL  FILL_2742
timestamp 1677677812
transform 1 0 184 0 1 3370
box -8 -3 16 105
use FILL  FILL_2743
timestamp 1677677812
transform 1 0 192 0 1 3370
box -8 -3 16 105
use FILL  FILL_2744
timestamp 1677677812
transform 1 0 200 0 1 3370
box -8 -3 16 105
use FILL  FILL_2745
timestamp 1677677812
transform 1 0 208 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_119
timestamp 1677677812
transform 1 0 216 0 1 3370
box -8 -3 46 105
use FILL  FILL_2749
timestamp 1677677812
transform 1 0 256 0 1 3370
box -8 -3 16 105
use FILL  FILL_2750
timestamp 1677677812
transform 1 0 264 0 1 3370
box -8 -3 16 105
use FILL  FILL_2753
timestamp 1677677812
transform 1 0 272 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_188
timestamp 1677677812
transform 1 0 280 0 1 3370
box -8 -3 104 105
use FILL  FILL_2755
timestamp 1677677812
transform 1 0 376 0 1 3370
box -8 -3 16 105
use FILL  FILL_2756
timestamp 1677677812
transform 1 0 384 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_217
timestamp 1677677812
transform 1 0 392 0 1 3370
box -9 -3 26 105
use FILL  FILL_2757
timestamp 1677677812
transform 1 0 408 0 1 3370
box -8 -3 16 105
use FILL  FILL_2758
timestamp 1677677812
transform 1 0 416 0 1 3370
box -8 -3 16 105
use FILL  FILL_2767
timestamp 1677677812
transform 1 0 424 0 1 3370
box -8 -3 16 105
use FILL  FILL_2769
timestamp 1677677812
transform 1 0 432 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_121
timestamp 1677677812
transform -1 0 480 0 1 3370
box -8 -3 46 105
use FILL  FILL_2770
timestamp 1677677812
transform 1 0 480 0 1 3370
box -8 -3 16 105
use FILL  FILL_2771
timestamp 1677677812
transform 1 0 488 0 1 3370
box -8 -3 16 105
use FILL  FILL_2772
timestamp 1677677812
transform 1 0 496 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_218
timestamp 1677677812
transform 1 0 504 0 1 3370
box -9 -3 26 105
use FILL  FILL_2773
timestamp 1677677812
transform 1 0 520 0 1 3370
box -8 -3 16 105
use FILL  FILL_2781
timestamp 1677677812
transform 1 0 528 0 1 3370
box -8 -3 16 105
use FILL  FILL_2783
timestamp 1677677812
transform 1 0 536 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2455
timestamp 1677677812
transform 1 0 588 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_189
timestamp 1677677812
transform 1 0 544 0 1 3370
box -8 -3 104 105
use FILL  FILL_2785
timestamp 1677677812
transform 1 0 640 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2456
timestamp 1677677812
transform 1 0 676 0 1 3375
box -3 -3 3 3
use BUFX2  BUFX2_16
timestamp 1677677812
transform 1 0 648 0 1 3370
box -5 -3 28 105
use FILL  FILL_2786
timestamp 1677677812
transform 1 0 672 0 1 3370
box -8 -3 16 105
use FILL  FILL_2792
timestamp 1677677812
transform 1 0 680 0 1 3370
box -8 -3 16 105
use FILL  FILL_2794
timestamp 1677677812
transform 1 0 688 0 1 3370
box -8 -3 16 105
use FILL  FILL_2796
timestamp 1677677812
transform 1 0 696 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_28
timestamp 1677677812
transform 1 0 704 0 1 3370
box -8 -3 32 105
use FILL  FILL_2797
timestamp 1677677812
transform 1 0 728 0 1 3370
box -8 -3 16 105
use FILL  FILL_2798
timestamp 1677677812
transform 1 0 736 0 1 3370
box -8 -3 16 105
use FILL  FILL_2800
timestamp 1677677812
transform 1 0 744 0 1 3370
box -8 -3 16 105
use FILL  FILL_2802
timestamp 1677677812
transform 1 0 752 0 1 3370
box -8 -3 16 105
use FILL  FILL_2804
timestamp 1677677812
transform 1 0 760 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_191
timestamp 1677677812
transform 1 0 768 0 1 3370
box -8 -3 104 105
use FILL  FILL_2806
timestamp 1677677812
transform 1 0 864 0 1 3370
box -8 -3 16 105
use FILL  FILL_2807
timestamp 1677677812
transform 1 0 872 0 1 3370
box -8 -3 16 105
use FILL  FILL_2808
timestamp 1677677812
transform 1 0 880 0 1 3370
box -8 -3 16 105
use FILL  FILL_2809
timestamp 1677677812
transform 1 0 888 0 1 3370
box -8 -3 16 105
use FILL  FILL_2810
timestamp 1677677812
transform 1 0 896 0 1 3370
box -8 -3 16 105
use FILL  FILL_2811
timestamp 1677677812
transform 1 0 904 0 1 3370
box -8 -3 16 105
use FILL  FILL_2812
timestamp 1677677812
transform 1 0 912 0 1 3370
box -8 -3 16 105
use FILL  FILL_2813
timestamp 1677677812
transform 1 0 920 0 1 3370
box -8 -3 16 105
use FILL  FILL_2814
timestamp 1677677812
transform 1 0 928 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2457
timestamp 1677677812
transform 1 0 948 0 1 3375
box -3 -3 3 3
use FILL  FILL_2815
timestamp 1677677812
transform 1 0 936 0 1 3370
box -8 -3 16 105
use FILL  FILL_2816
timestamp 1677677812
transform 1 0 944 0 1 3370
box -8 -3 16 105
use FILL  FILL_2817
timestamp 1677677812
transform 1 0 952 0 1 3370
box -8 -3 16 105
use FILL  FILL_2818
timestamp 1677677812
transform 1 0 960 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_29
timestamp 1677677812
transform 1 0 968 0 1 3370
box -8 -3 32 105
use FILL  FILL_2830
timestamp 1677677812
transform 1 0 992 0 1 3370
box -8 -3 16 105
use FILL  FILL_2831
timestamp 1677677812
transform 1 0 1000 0 1 3370
box -8 -3 16 105
use FILL  FILL_2835
timestamp 1677677812
transform 1 0 1008 0 1 3370
box -8 -3 16 105
use FILL  FILL_2837
timestamp 1677677812
transform 1 0 1016 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2458
timestamp 1677677812
transform 1 0 1036 0 1 3375
box -3 -3 3 3
use FILL  FILL_2839
timestamp 1677677812
transform 1 0 1024 0 1 3370
box -8 -3 16 105
use FILL  FILL_2841
timestamp 1677677812
transform 1 0 1032 0 1 3370
box -8 -3 16 105
use FILL  FILL_2843
timestamp 1677677812
transform 1 0 1040 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_62
timestamp 1677677812
transform 1 0 1048 0 1 3370
box -8 -3 34 105
use FILL  FILL_2845
timestamp 1677677812
transform 1 0 1080 0 1 3370
box -8 -3 16 105
use FILL  FILL_2846
timestamp 1677677812
transform 1 0 1088 0 1 3370
box -8 -3 16 105
use FILL  FILL_2848
timestamp 1677677812
transform 1 0 1096 0 1 3370
box -8 -3 16 105
use FILL  FILL_2850
timestamp 1677677812
transform 1 0 1104 0 1 3370
box -8 -3 16 105
use FILL  FILL_2852
timestamp 1677677812
transform 1 0 1112 0 1 3370
box -8 -3 16 105
use FILL  FILL_2854
timestamp 1677677812
transform 1 0 1120 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_128
timestamp 1677677812
transform 1 0 1128 0 1 3370
box -8 -3 46 105
use FILL  FILL_2856
timestamp 1677677812
transform 1 0 1168 0 1 3370
box -8 -3 16 105
use FILL  FILL_2857
timestamp 1677677812
transform 1 0 1176 0 1 3370
box -8 -3 16 105
use FILL  FILL_2861
timestamp 1677677812
transform 1 0 1184 0 1 3370
box -8 -3 16 105
use FILL  FILL_2863
timestamp 1677677812
transform 1 0 1192 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2459
timestamp 1677677812
transform 1 0 1212 0 1 3375
box -3 -3 3 3
use FILL  FILL_2865
timestamp 1677677812
transform 1 0 1200 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_221
timestamp 1677677812
transform 1 0 1208 0 1 3370
box -9 -3 26 105
use FILL  FILL_2867
timestamp 1677677812
transform 1 0 1224 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2460
timestamp 1677677812
transform 1 0 1244 0 1 3375
box -3 -3 3 3
use FILL  FILL_2868
timestamp 1677677812
transform 1 0 1232 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_193
timestamp 1677677812
transform -1 0 1336 0 1 3370
box -8 -3 104 105
use FILL  FILL_2869
timestamp 1677677812
transform 1 0 1336 0 1 3370
box -8 -3 16 105
use FILL  FILL_2880
timestamp 1677677812
transform 1 0 1344 0 1 3370
box -8 -3 16 105
use BUFX2  BUFX2_17
timestamp 1677677812
transform -1 0 1376 0 1 3370
box -5 -3 28 105
use FILL  FILL_2881
timestamp 1677677812
transform 1 0 1376 0 1 3370
box -8 -3 16 105
use FILL  FILL_2882
timestamp 1677677812
transform 1 0 1384 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2461
timestamp 1677677812
transform 1 0 1428 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_194
timestamp 1677677812
transform 1 0 1392 0 1 3370
box -8 -3 104 105
use INVX2  INVX2_222
timestamp 1677677812
transform 1 0 1488 0 1 3370
box -9 -3 26 105
use FILL  FILL_2885
timestamp 1677677812
transform 1 0 1504 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2462
timestamp 1677677812
transform 1 0 1596 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_195
timestamp 1677677812
transform -1 0 1608 0 1 3370
box -8 -3 104 105
use FILL  FILL_2886
timestamp 1677677812
transform 1 0 1608 0 1 3370
box -8 -3 16 105
use FILL  FILL_2908
timestamp 1677677812
transform 1 0 1616 0 1 3370
box -8 -3 16 105
use FILL  FILL_2909
timestamp 1677677812
transform 1 0 1624 0 1 3370
box -8 -3 16 105
use FILL  FILL_2910
timestamp 1677677812
transform 1 0 1632 0 1 3370
box -8 -3 16 105
use FILL  FILL_2911
timestamp 1677677812
transform 1 0 1640 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_196
timestamp 1677677812
transform 1 0 1648 0 1 3370
box -8 -3 104 105
use FILL  FILL_2912
timestamp 1677677812
transform 1 0 1744 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_224
timestamp 1677677812
transform -1 0 1768 0 1 3370
box -9 -3 26 105
use BUFX2  BUFX2_18
timestamp 1677677812
transform 1 0 1768 0 1 3370
box -5 -3 28 105
use FILL  FILL_2913
timestamp 1677677812
transform 1 0 1792 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2463
timestamp 1677677812
transform 1 0 1812 0 1 3375
box -3 -3 3 3
use FILL  FILL_2914
timestamp 1677677812
transform 1 0 1800 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_197
timestamp 1677677812
transform -1 0 1904 0 1 3370
box -8 -3 104 105
use FILL  FILL_2915
timestamp 1677677812
transform 1 0 1904 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_198
timestamp 1677677812
transform 1 0 1912 0 1 3370
box -8 -3 104 105
use FILL  FILL_2938
timestamp 1677677812
transform 1 0 2008 0 1 3370
box -8 -3 16 105
use FILL  FILL_2939
timestamp 1677677812
transform 1 0 2016 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_226
timestamp 1677677812
transform -1 0 2040 0 1 3370
box -9 -3 26 105
use FILL  FILL_2940
timestamp 1677677812
transform 1 0 2040 0 1 3370
box -8 -3 16 105
use FILL  FILL_2941
timestamp 1677677812
transform 1 0 2048 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_199
timestamp 1677677812
transform 1 0 2056 0 1 3370
box -8 -3 104 105
use M3_M2  M3_M2_2464
timestamp 1677677812
transform 1 0 2164 0 1 3375
box -3 -3 3 3
use FILL  FILL_2942
timestamp 1677677812
transform 1 0 2152 0 1 3370
box -8 -3 16 105
use FILL  FILL_2943
timestamp 1677677812
transform 1 0 2160 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_227
timestamp 1677677812
transform 1 0 2168 0 1 3370
box -9 -3 26 105
use FILL  FILL_2944
timestamp 1677677812
transform 1 0 2184 0 1 3370
box -8 -3 16 105
use FILL  FILL_2945
timestamp 1677677812
transform 1 0 2192 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_200
timestamp 1677677812
transform -1 0 2296 0 1 3370
box -8 -3 104 105
use FILL  FILL_2946
timestamp 1677677812
transform 1 0 2296 0 1 3370
box -8 -3 16 105
use FILL  FILL_2972
timestamp 1677677812
transform 1 0 2304 0 1 3370
box -8 -3 16 105
use FILL  FILL_2974
timestamp 1677677812
transform 1 0 2312 0 1 3370
box -8 -3 16 105
use FILL  FILL_2976
timestamp 1677677812
transform 1 0 2320 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_126
timestamp 1677677812
transform 1 0 2328 0 1 3370
box -8 -3 46 105
use FILL  FILL_2977
timestamp 1677677812
transform 1 0 2368 0 1 3370
box -8 -3 16 105
use FILL  FILL_2978
timestamp 1677677812
transform 1 0 2376 0 1 3370
box -8 -3 16 105
use AND2X2  AND2X2_5
timestamp 1677677812
transform -1 0 2416 0 1 3370
box -8 -3 40 105
use FILL  FILL_2979
timestamp 1677677812
transform 1 0 2416 0 1 3370
box -8 -3 16 105
use FILL  FILL_2981
timestamp 1677677812
transform 1 0 2424 0 1 3370
box -8 -3 16 105
use FILL  FILL_2983
timestamp 1677677812
transform 1 0 2432 0 1 3370
box -8 -3 16 105
use FILL  FILL_2985
timestamp 1677677812
transform 1 0 2440 0 1 3370
box -8 -3 16 105
use FILL  FILL_2987
timestamp 1677677812
transform 1 0 2448 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_31
timestamp 1677677812
transform 1 0 2456 0 1 3370
box -8 -3 32 105
use FILL  FILL_2989
timestamp 1677677812
transform 1 0 2480 0 1 3370
box -8 -3 16 105
use FILL  FILL_2994
timestamp 1677677812
transform 1 0 2488 0 1 3370
box -8 -3 16 105
use FILL  FILL_2996
timestamp 1677677812
transform 1 0 2496 0 1 3370
box -8 -3 16 105
use FILL  FILL_2998
timestamp 1677677812
transform 1 0 2504 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_131
timestamp 1677677812
transform 1 0 2512 0 1 3370
box -8 -3 46 105
use FILL  FILL_3000
timestamp 1677677812
transform 1 0 2552 0 1 3370
box -8 -3 16 105
use FILL  FILL_3001
timestamp 1677677812
transform 1 0 2560 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_229
timestamp 1677677812
transform 1 0 2568 0 1 3370
box -9 -3 26 105
use FILL  FILL_3002
timestamp 1677677812
transform 1 0 2584 0 1 3370
box -8 -3 16 105
use FILL  FILL_3003
timestamp 1677677812
transform 1 0 2592 0 1 3370
box -8 -3 16 105
use FILL  FILL_3004
timestamp 1677677812
transform 1 0 2600 0 1 3370
box -8 -3 16 105
use FILL  FILL_3005
timestamp 1677677812
transform 1 0 2608 0 1 3370
box -8 -3 16 105
use FILL  FILL_3006
timestamp 1677677812
transform 1 0 2616 0 1 3370
box -8 -3 16 105
use FILL  FILL_3007
timestamp 1677677812
transform 1 0 2624 0 1 3370
box -8 -3 16 105
use FILL  FILL_3008
timestamp 1677677812
transform 1 0 2632 0 1 3370
box -8 -3 16 105
use FILL  FILL_3009
timestamp 1677677812
transform 1 0 2640 0 1 3370
box -8 -3 16 105
use FILL  FILL_3010
timestamp 1677677812
transform 1 0 2648 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_132
timestamp 1677677812
transform 1 0 2656 0 1 3370
box -8 -3 46 105
use FILL  FILL_3015
timestamp 1677677812
transform 1 0 2696 0 1 3370
box -8 -3 16 105
use FILL  FILL_3016
timestamp 1677677812
transform 1 0 2704 0 1 3370
box -8 -3 16 105
use AND2X2  AND2X2_6
timestamp 1677677812
transform -1 0 2744 0 1 3370
box -8 -3 40 105
use FILL  FILL_3017
timestamp 1677677812
transform 1 0 2744 0 1 3370
box -8 -3 16 105
use FILL  FILL_3018
timestamp 1677677812
transform 1 0 2752 0 1 3370
box -8 -3 16 105
use FILL  FILL_3019
timestamp 1677677812
transform 1 0 2760 0 1 3370
box -8 -3 16 105
use FILL  FILL_3020
timestamp 1677677812
transform 1 0 2768 0 1 3370
box -8 -3 16 105
use FILL  FILL_3021
timestamp 1677677812
transform 1 0 2776 0 1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_32
timestamp 1677677812
transform 1 0 2784 0 1 3370
box -8 -3 32 105
use FILL  FILL_3022
timestamp 1677677812
transform 1 0 2808 0 1 3370
box -8 -3 16 105
use FILL  FILL_3023
timestamp 1677677812
transform 1 0 2816 0 1 3370
box -8 -3 16 105
use FILL  FILL_3024
timestamp 1677677812
transform 1 0 2824 0 1 3370
box -8 -3 16 105
use FILL  FILL_3025
timestamp 1677677812
transform 1 0 2832 0 1 3370
box -8 -3 16 105
use FILL  FILL_3026
timestamp 1677677812
transform 1 0 2840 0 1 3370
box -8 -3 16 105
use FILL  FILL_3027
timestamp 1677677812
transform 1 0 2848 0 1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_66
timestamp 1677677812
transform 1 0 2856 0 1 3370
box -8 -3 34 105
use FILL  FILL_3037
timestamp 1677677812
transform 1 0 2888 0 1 3370
box -8 -3 16 105
use FILL  FILL_3039
timestamp 1677677812
transform 1 0 2896 0 1 3370
box -8 -3 16 105
use FILL  FILL_3040
timestamp 1677677812
transform 1 0 2904 0 1 3370
box -8 -3 16 105
use FILL  FILL_3041
timestamp 1677677812
transform 1 0 2912 0 1 3370
box -8 -3 16 105
use FILL  FILL_3042
timestamp 1677677812
transform 1 0 2920 0 1 3370
box -8 -3 16 105
use FILL  FILL_3043
timestamp 1677677812
transform 1 0 2928 0 1 3370
box -8 -3 16 105
use AND2X2  AND2X2_7
timestamp 1677677812
transform 1 0 2936 0 1 3370
box -8 -3 40 105
use FILL  FILL_3045
timestamp 1677677812
transform 1 0 2968 0 1 3370
box -8 -3 16 105
use FILL  FILL_3046
timestamp 1677677812
transform 1 0 2976 0 1 3370
box -8 -3 16 105
use FILL  FILL_3047
timestamp 1677677812
transform 1 0 2984 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2465
timestamp 1677677812
transform 1 0 3004 0 1 3375
box -3 -3 3 3
use FILL  FILL_3048
timestamp 1677677812
transform 1 0 2992 0 1 3370
box -8 -3 16 105
use FILL  FILL_3049
timestamp 1677677812
transform 1 0 3000 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_205
timestamp 1677677812
transform 1 0 3008 0 1 3370
box -8 -3 104 105
use FILL  FILL_3055
timestamp 1677677812
transform 1 0 3104 0 1 3370
box -8 -3 16 105
use FILL  FILL_3065
timestamp 1677677812
transform 1 0 3112 0 1 3370
box -8 -3 16 105
use FILL  FILL_3067
timestamp 1677677812
transform 1 0 3120 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_206
timestamp 1677677812
transform 1 0 3128 0 1 3370
box -8 -3 104 105
use FILL  FILL_3069
timestamp 1677677812
transform 1 0 3224 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2466
timestamp 1677677812
transform 1 0 3252 0 1 3375
box -3 -3 3 3
use M3_M2  M3_M2_2467
timestamp 1677677812
transform 1 0 3316 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_207
timestamp 1677677812
transform 1 0 3232 0 1 3370
box -8 -3 104 105
use FILL  FILL_3076
timestamp 1677677812
transform 1 0 3328 0 1 3370
box -8 -3 16 105
use AND2X2  AND2X2_8
timestamp 1677677812
transform 1 0 3336 0 1 3370
box -8 -3 40 105
use M3_M2  M3_M2_2468
timestamp 1677677812
transform 1 0 3380 0 1 3375
box -3 -3 3 3
use FILL  FILL_3077
timestamp 1677677812
transform 1 0 3368 0 1 3370
box -8 -3 16 105
use FILL  FILL_3089
timestamp 1677677812
transform 1 0 3376 0 1 3370
box -8 -3 16 105
use FILL  FILL_3090
timestamp 1677677812
transform 1 0 3384 0 1 3370
box -8 -3 16 105
use FILL  FILL_3091
timestamp 1677677812
transform 1 0 3392 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2469
timestamp 1677677812
transform 1 0 3420 0 1 3375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_208
timestamp 1677677812
transform 1 0 3400 0 1 3370
box -8 -3 104 105
use FILL  FILL_3092
timestamp 1677677812
transform 1 0 3496 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2470
timestamp 1677677812
transform 1 0 3516 0 1 3375
box -3 -3 3 3
use FILL  FILL_3100
timestamp 1677677812
transform 1 0 3504 0 1 3370
box -8 -3 16 105
use FILL  FILL_3102
timestamp 1677677812
transform 1 0 3512 0 1 3370
box -8 -3 16 105
use FILL  FILL_3103
timestamp 1677677812
transform 1 0 3520 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2471
timestamp 1677677812
transform 1 0 3572 0 1 3375
box -3 -3 3 3
use OAI22X1  OAI22X1_129
timestamp 1677677812
transform -1 0 3568 0 1 3370
box -8 -3 46 105
use FILL  FILL_3104
timestamp 1677677812
transform 1 0 3568 0 1 3370
box -8 -3 16 105
use FILL  FILL_3105
timestamp 1677677812
transform 1 0 3576 0 1 3370
box -8 -3 16 105
use FILL  FILL_3106
timestamp 1677677812
transform 1 0 3584 0 1 3370
box -8 -3 16 105
use FILL  FILL_3107
timestamp 1677677812
transform 1 0 3592 0 1 3370
box -8 -3 16 105
use FILL  FILL_3108
timestamp 1677677812
transform 1 0 3600 0 1 3370
box -8 -3 16 105
use FILL  FILL_3109
timestamp 1677677812
transform 1 0 3608 0 1 3370
box -8 -3 16 105
use FILL  FILL_3110
timestamp 1677677812
transform 1 0 3616 0 1 3370
box -8 -3 16 105
use FILL  FILL_3111
timestamp 1677677812
transform 1 0 3624 0 1 3370
box -8 -3 16 105
use FILL  FILL_3112
timestamp 1677677812
transform 1 0 3632 0 1 3370
box -8 -3 16 105
use FILL  FILL_3113
timestamp 1677677812
transform 1 0 3640 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_130
timestamp 1677677812
transform -1 0 3688 0 1 3370
box -8 -3 46 105
use FILL  FILL_3114
timestamp 1677677812
transform 1 0 3688 0 1 3370
box -8 -3 16 105
use FILL  FILL_3115
timestamp 1677677812
transform 1 0 3696 0 1 3370
box -8 -3 16 105
use FILL  FILL_3116
timestamp 1677677812
transform 1 0 3704 0 1 3370
box -8 -3 16 105
use AND2X2  AND2X2_9
timestamp 1677677812
transform 1 0 3712 0 1 3370
box -8 -3 40 105
use FILL  FILL_3117
timestamp 1677677812
transform 1 0 3744 0 1 3370
box -8 -3 16 105
use FILL  FILL_3118
timestamp 1677677812
transform 1 0 3752 0 1 3370
box -8 -3 16 105
use FILL  FILL_3119
timestamp 1677677812
transform 1 0 3760 0 1 3370
box -8 -3 16 105
use FILL  FILL_3120
timestamp 1677677812
transform 1 0 3768 0 1 3370
box -8 -3 16 105
use FILL  FILL_3121
timestamp 1677677812
transform 1 0 3776 0 1 3370
box -8 -3 16 105
use FILL  FILL_3122
timestamp 1677677812
transform 1 0 3784 0 1 3370
box -8 -3 16 105
use FILL  FILL_3123
timestamp 1677677812
transform 1 0 3792 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2472
timestamp 1677677812
transform 1 0 3812 0 1 3375
box -3 -3 3 3
use FILL  FILL_3124
timestamp 1677677812
transform 1 0 3800 0 1 3370
box -8 -3 16 105
use FILL  FILL_3125
timestamp 1677677812
transform 1 0 3808 0 1 3370
box -8 -3 16 105
use FILL  FILL_3132
timestamp 1677677812
transform 1 0 3816 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2473
timestamp 1677677812
transform 1 0 3836 0 1 3375
box -3 -3 3 3
use FILL  FILL_3134
timestamp 1677677812
transform 1 0 3824 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_131
timestamp 1677677812
transform 1 0 3832 0 1 3370
box -8 -3 46 105
use FILL  FILL_3136
timestamp 1677677812
transform 1 0 3872 0 1 3370
box -8 -3 16 105
use FILL  FILL_3137
timestamp 1677677812
transform 1 0 3880 0 1 3370
box -8 -3 16 105
use FILL  FILL_3138
timestamp 1677677812
transform 1 0 3888 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_211
timestamp 1677677812
transform 1 0 3896 0 1 3370
box -8 -3 104 105
use FILL  FILL_3142
timestamp 1677677812
transform 1 0 3992 0 1 3370
box -8 -3 16 105
use FILL  FILL_3143
timestamp 1677677812
transform 1 0 4000 0 1 3370
box -8 -3 16 105
use FILL  FILL_3144
timestamp 1677677812
transform 1 0 4008 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_132
timestamp 1677677812
transform 1 0 4016 0 1 3370
box -8 -3 46 105
use FILL  FILL_3145
timestamp 1677677812
transform 1 0 4056 0 1 3370
box -8 -3 16 105
use FILL  FILL_3153
timestamp 1677677812
transform 1 0 4064 0 1 3370
box -8 -3 16 105
use FILL  FILL_3155
timestamp 1677677812
transform 1 0 4072 0 1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2474
timestamp 1677677812
transform 1 0 4092 0 1 3375
box -3 -3 3 3
use FILL  FILL_3157
timestamp 1677677812
transform 1 0 4080 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_213
timestamp 1677677812
transform 1 0 4088 0 1 3370
box -8 -3 104 105
use FILL  FILL_3158
timestamp 1677677812
transform 1 0 4184 0 1 3370
box -8 -3 16 105
use FILL  FILL_3161
timestamp 1677677812
transform 1 0 4192 0 1 3370
box -8 -3 16 105
use FILL  FILL_3163
timestamp 1677677812
transform 1 0 4200 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_133
timestamp 1677677812
transform 1 0 4208 0 1 3370
box -8 -3 46 105
use FILL  FILL_3165
timestamp 1677677812
transform 1 0 4248 0 1 3370
box -8 -3 16 105
use FILL  FILL_3166
timestamp 1677677812
transform 1 0 4256 0 1 3370
box -8 -3 16 105
use FILL  FILL_3167
timestamp 1677677812
transform 1 0 4264 0 1 3370
box -8 -3 16 105
use FILL  FILL_3168
timestamp 1677677812
transform 1 0 4272 0 1 3370
box -8 -3 16 105
use FILL  FILL_3169
timestamp 1677677812
transform 1 0 4280 0 1 3370
box -8 -3 16 105
use FILL  FILL_3170
timestamp 1677677812
transform 1 0 4288 0 1 3370
box -8 -3 16 105
use BUFX2  BUFX2_20
timestamp 1677677812
transform -1 0 4320 0 1 3370
box -5 -3 28 105
use FILL  FILL_3171
timestamp 1677677812
transform 1 0 4320 0 1 3370
box -8 -3 16 105
use FILL  FILL_3172
timestamp 1677677812
transform 1 0 4328 0 1 3370
box -8 -3 16 105
use FILL  FILL_3173
timestamp 1677677812
transform 1 0 4336 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_135
timestamp 1677677812
transform -1 0 4384 0 1 3370
box -8 -3 46 105
use FILL  FILL_3174
timestamp 1677677812
transform 1 0 4384 0 1 3370
box -8 -3 16 105
use FILL  FILL_3175
timestamp 1677677812
transform 1 0 4392 0 1 3370
box -8 -3 16 105
use FILL  FILL_3176
timestamp 1677677812
transform 1 0 4400 0 1 3370
box -8 -3 16 105
use FILL  FILL_3177
timestamp 1677677812
transform 1 0 4408 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_238
timestamp 1677677812
transform -1 0 4432 0 1 3370
box -9 -3 26 105
use FILL  FILL_3178
timestamp 1677677812
transform 1 0 4432 0 1 3370
box -8 -3 16 105
use FILL  FILL_3192
timestamp 1677677812
transform 1 0 4440 0 1 3370
box -8 -3 16 105
use FILL  FILL_3194
timestamp 1677677812
transform 1 0 4448 0 1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_137
timestamp 1677677812
transform 1 0 4456 0 1 3370
box -8 -3 46 105
use FILL  FILL_3196
timestamp 1677677812
transform 1 0 4496 0 1 3370
box -8 -3 16 105
use FILL  FILL_3197
timestamp 1677677812
transform 1 0 4504 0 1 3370
box -8 -3 16 105
use FILL  FILL_3198
timestamp 1677677812
transform 1 0 4512 0 1 3370
box -8 -3 16 105
use FILL  FILL_3199
timestamp 1677677812
transform 1 0 4520 0 1 3370
box -8 -3 16 105
use FILL  FILL_3204
timestamp 1677677812
transform 1 0 4528 0 1 3370
box -8 -3 16 105
use FILL  FILL_3206
timestamp 1677677812
transform 1 0 4536 0 1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_215
timestamp 1677677812
transform 1 0 4544 0 1 3370
box -8 -3 104 105
use INVX2  INVX2_241
timestamp 1677677812
transform -1 0 4656 0 1 3370
box -9 -3 26 105
use FILL  FILL_3208
timestamp 1677677812
transform 1 0 4656 0 1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_136
timestamp 1677677812
transform 1 0 4664 0 1 3370
box -8 -3 46 105
use FILL  FILL_3217
timestamp 1677677812
transform 1 0 4704 0 1 3370
box -8 -3 16 105
use FILL  FILL_3218
timestamp 1677677812
transform 1 0 4712 0 1 3370
box -8 -3 16 105
use FILL  FILL_3219
timestamp 1677677812
transform 1 0 4720 0 1 3370
box -8 -3 16 105
use FILL  FILL_3220
timestamp 1677677812
transform 1 0 4728 0 1 3370
box -8 -3 16 105
use FILL  FILL_3221
timestamp 1677677812
transform 1 0 4736 0 1 3370
box -8 -3 16 105
use INVX2  INVX2_243
timestamp 1677677812
transform -1 0 4760 0 1 3370
box -9 -3 26 105
use FILL  FILL_3222
timestamp 1677677812
transform 1 0 4760 0 1 3370
box -8 -3 16 105
use FILL  FILL_3223
timestamp 1677677812
transform 1 0 4768 0 1 3370
box -8 -3 16 105
use FILL  FILL_3224
timestamp 1677677812
transform 1 0 4776 0 1 3370
box -8 -3 16 105
use FILL  FILL_3225
timestamp 1677677812
transform 1 0 4784 0 1 3370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_27
timestamp 1677677812
transform 1 0 4819 0 1 3370
box -10 -3 10 3
use M3_M2  M3_M2_2535
timestamp 1677677812
transform 1 0 100 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2869
timestamp 1677677812
transform 1 0 180 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2956
timestamp 1677677812
transform 1 0 100 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2957
timestamp 1677677812
transform 1 0 148 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2958
timestamp 1677677812
transform 1 0 196 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2600
timestamp 1677677812
transform 1 0 148 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2601
timestamp 1677677812
transform 1 0 196 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2663
timestamp 1677677812
transform 1 0 180 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2536
timestamp 1677677812
transform 1 0 252 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2870
timestamp 1677677812
transform 1 0 228 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2871
timestamp 1677677812
transform 1 0 236 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2872
timestamp 1677677812
transform 1 0 252 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2873
timestamp 1677677812
transform 1 0 268 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2959
timestamp 1677677812
transform 1 0 228 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2960
timestamp 1677677812
transform 1 0 244 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2961
timestamp 1677677812
transform 1 0 260 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2602
timestamp 1677677812
transform 1 0 220 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2603
timestamp 1677677812
transform 1 0 244 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2604
timestamp 1677677812
transform 1 0 260 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2643
timestamp 1677677812
transform 1 0 236 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2537
timestamp 1677677812
transform 1 0 332 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2874
timestamp 1677677812
transform 1 0 316 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2875
timestamp 1677677812
transform 1 0 332 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2962
timestamp 1677677812
transform 1 0 308 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2573
timestamp 1677677812
transform 1 0 316 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2963
timestamp 1677677812
transform 1 0 324 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2475
timestamp 1677677812
transform 1 0 356 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2664
timestamp 1677677812
transform 1 0 356 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2510
timestamp 1677677812
transform 1 0 372 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2876
timestamp 1677677812
transform 1 0 372 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2964
timestamp 1677677812
transform 1 0 372 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2965
timestamp 1677677812
transform 1 0 396 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2877
timestamp 1677677812
transform 1 0 436 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2966
timestamp 1677677812
transform 1 0 444 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2538
timestamp 1677677812
transform 1 0 508 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2878
timestamp 1677677812
transform 1 0 484 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2879
timestamp 1677677812
transform 1 0 508 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2967
timestamp 1677677812
transform 1 0 492 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2968
timestamp 1677677812
transform 1 0 508 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2605
timestamp 1677677812
transform 1 0 508 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2644
timestamp 1677677812
transform 1 0 484 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2476
timestamp 1677677812
transform 1 0 556 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2477
timestamp 1677677812
transform 1 0 612 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2539
timestamp 1677677812
transform 1 0 644 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2880
timestamp 1677677812
transform 1 0 564 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2969
timestamp 1677677812
transform 1 0 604 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2970
timestamp 1677677812
transform 1 0 644 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2606
timestamp 1677677812
transform 1 0 564 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2645
timestamp 1677677812
transform 1 0 588 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2478
timestamp 1677677812
transform 1 0 660 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2540
timestamp 1677677812
transform 1 0 660 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2881
timestamp 1677677812
transform 1 0 660 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2479
timestamp 1677677812
transform 1 0 716 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2511
timestamp 1677677812
transform 1 0 732 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2882
timestamp 1677677812
transform 1 0 716 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2883
timestamp 1677677812
transform 1 0 732 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2971
timestamp 1677677812
transform 1 0 708 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2972
timestamp 1677677812
transform 1 0 724 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2646
timestamp 1677677812
transform 1 0 724 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2512
timestamp 1677677812
transform 1 0 780 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2884
timestamp 1677677812
transform 1 0 788 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2973
timestamp 1677677812
transform 1 0 812 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2574
timestamp 1677677812
transform 1 0 820 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2885
timestamp 1677677812
transform 1 0 876 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2974
timestamp 1677677812
transform 1 0 924 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2575
timestamp 1677677812
transform 1 0 948 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2975
timestamp 1677677812
transform 1 0 956 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2976
timestamp 1677677812
transform 1 0 964 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2607
timestamp 1677677812
transform 1 0 924 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2665
timestamp 1677677812
transform 1 0 900 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2666
timestamp 1677677812
transform 1 0 924 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2608
timestamp 1677677812
transform 1 0 964 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2977
timestamp 1677677812
transform 1 0 996 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2886
timestamp 1677677812
transform 1 0 1028 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2609
timestamp 1677677812
transform 1 0 1028 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2541
timestamp 1677677812
transform 1 0 1084 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2887
timestamp 1677677812
transform 1 0 1060 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2888
timestamp 1677677812
transform 1 0 1076 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2978
timestamp 1677677812
transform 1 0 1068 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2576
timestamp 1677677812
transform 1 0 1076 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2979
timestamp 1677677812
transform 1 0 1084 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2610
timestamp 1677677812
transform 1 0 1068 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2480
timestamp 1677677812
transform 1 0 1180 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2542
timestamp 1677677812
transform 1 0 1172 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2554
timestamp 1677677812
transform 1 0 1164 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2889
timestamp 1677677812
transform 1 0 1172 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2980
timestamp 1677677812
transform 1 0 1156 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2868
timestamp 1677677812
transform 1 0 1180 0 1 3345
box -2 -2 2 2
use M3_M2  M3_M2_2555
timestamp 1677677812
transform 1 0 1204 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2890
timestamp 1677677812
transform 1 0 1212 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2577
timestamp 1677677812
transform 1 0 1204 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3059
timestamp 1677677812
transform 1 0 1204 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2891
timestamp 1677677812
transform 1 0 1228 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2543
timestamp 1677677812
transform 1 0 1260 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2981
timestamp 1677677812
transform 1 0 1260 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2544
timestamp 1677677812
transform 1 0 1300 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2556
timestamp 1677677812
transform 1 0 1284 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2892
timestamp 1677677812
transform 1 0 1300 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2982
timestamp 1677677812
transform 1 0 1284 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2893
timestamp 1677677812
transform 1 0 1308 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2578
timestamp 1677677812
transform 1 0 1308 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3060
timestamp 1677677812
transform 1 0 1308 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2513
timestamp 1677677812
transform 1 0 1324 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2983
timestamp 1677677812
transform 1 0 1324 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2579
timestamp 1677677812
transform 1 0 1364 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2984
timestamp 1677677812
transform 1 0 1380 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2481
timestamp 1677677812
transform 1 0 1460 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2482
timestamp 1677677812
transform 1 0 1484 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2894
timestamp 1677677812
transform 1 0 1452 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2895
timestamp 1677677812
transform 1 0 1460 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2896
timestamp 1677677812
transform 1 0 1476 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2985
timestamp 1677677812
transform 1 0 1460 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2611
timestamp 1677677812
transform 1 0 1452 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2580
timestamp 1677677812
transform 1 0 1476 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2986
timestamp 1677677812
transform 1 0 1484 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2667
timestamp 1677677812
transform 1 0 1460 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2545
timestamp 1677677812
transform 1 0 1508 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2897
timestamp 1677677812
transform 1 0 1508 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2898
timestamp 1677677812
transform 1 0 1516 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2581
timestamp 1677677812
transform 1 0 1516 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_2987
timestamp 1677677812
transform 1 0 1556 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2546
timestamp 1677677812
transform 1 0 1580 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2899
timestamp 1677677812
transform 1 0 1580 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2582
timestamp 1677677812
transform 1 0 1572 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2647
timestamp 1677677812
transform 1 0 1588 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2668
timestamp 1677677812
transform 1 0 1580 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2483
timestamp 1677677812
transform 1 0 1612 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2900
timestamp 1677677812
transform 1 0 1644 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2988
timestamp 1677677812
transform 1 0 1636 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2989
timestamp 1677677812
transform 1 0 1652 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2612
timestamp 1677677812
transform 1 0 1636 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2669
timestamp 1677677812
transform 1 0 1652 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2484
timestamp 1677677812
transform 1 0 1668 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2485
timestamp 1677677812
transform 1 0 1692 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2547
timestamp 1677677812
transform 1 0 1716 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2901
timestamp 1677677812
transform 1 0 1716 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2990
timestamp 1677677812
transform 1 0 1724 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2902
timestamp 1677677812
transform 1 0 1780 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2903
timestamp 1677677812
transform 1 0 1788 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2904
timestamp 1677677812
transform 1 0 1804 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2613
timestamp 1677677812
transform 1 0 1780 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2991
timestamp 1677677812
transform 1 0 1796 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2992
timestamp 1677677812
transform 1 0 1812 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2614
timestamp 1677677812
transform 1 0 1812 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2648
timestamp 1677677812
transform 1 0 1804 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2548
timestamp 1677677812
transform 1 0 1828 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2905
timestamp 1677677812
transform 1 0 1836 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2993
timestamp 1677677812
transform 1 0 1844 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2994
timestamp 1677677812
transform 1 0 1924 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2514
timestamp 1677677812
transform 1 0 1940 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2486
timestamp 1677677812
transform 1 0 1972 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2515
timestamp 1677677812
transform 1 0 1964 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2906
timestamp 1677677812
transform 1 0 1972 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2487
timestamp 1677677812
transform 1 0 2068 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2995
timestamp 1677677812
transform 1 0 2004 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2996
timestamp 1677677812
transform 1 0 2052 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2997
timestamp 1677677812
transform 1 0 2060 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2516
timestamp 1677677812
transform 1 0 2124 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2907
timestamp 1677677812
transform 1 0 2148 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2908
timestamp 1677677812
transform 1 0 2180 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2557
timestamp 1677677812
transform 1 0 2196 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2998
timestamp 1677677812
transform 1 0 2156 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_2999
timestamp 1677677812
transform 1 0 2172 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3000
timestamp 1677677812
transform 1 0 2188 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2615
timestamp 1677677812
transform 1 0 2156 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2558
timestamp 1677677812
transform 1 0 2212 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2583
timestamp 1677677812
transform 1 0 2204 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2670
timestamp 1677677812
transform 1 0 2204 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2517
timestamp 1677677812
transform 1 0 2244 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2559
timestamp 1677677812
transform 1 0 2228 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2909
timestamp 1677677812
transform 1 0 2252 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2910
timestamp 1677677812
transform 1 0 2260 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3001
timestamp 1677677812
transform 1 0 2228 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3002
timestamp 1677677812
transform 1 0 2244 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2584
timestamp 1677677812
transform 1 0 2252 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3003
timestamp 1677677812
transform 1 0 2260 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3004
timestamp 1677677812
transform 1 0 2268 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2616
timestamp 1677677812
transform 1 0 2260 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2488
timestamp 1677677812
transform 1 0 2284 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2671
timestamp 1677677812
transform 1 0 2308 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2489
timestamp 1677677812
transform 1 0 2332 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2518
timestamp 1677677812
transform 1 0 2356 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2911
timestamp 1677677812
transform 1 0 2332 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2560
timestamp 1677677812
transform 1 0 2372 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3005
timestamp 1677677812
transform 1 0 2356 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2617
timestamp 1677677812
transform 1 0 2364 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2678
timestamp 1677677812
transform 1 0 2404 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_3006
timestamp 1677677812
transform 1 0 2420 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2490
timestamp 1677677812
transform 1 0 2436 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2679
timestamp 1677677812
transform 1 0 2460 0 1 3285
box -3 -3 3 3
use M2_M1  M2_M1_2912
timestamp 1677677812
transform 1 0 2532 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2491
timestamp 1677677812
transform 1 0 2596 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2519
timestamp 1677677812
transform 1 0 2572 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2520
timestamp 1677677812
transform 1 0 2620 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2913
timestamp 1677677812
transform 1 0 2636 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3007
timestamp 1677677812
transform 1 0 2548 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3008
timestamp 1677677812
transform 1 0 2556 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3009
timestamp 1677677812
transform 1 0 2596 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2618
timestamp 1677677812
transform 1 0 2548 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2619
timestamp 1677677812
transform 1 0 2596 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2649
timestamp 1677677812
transform 1 0 2564 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2561
timestamp 1677677812
transform 1 0 2652 0 1 3335
box -3 -3 3 3
use M3_M2  M3_M2_2521
timestamp 1677677812
transform 1 0 2676 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_3010
timestamp 1677677812
transform 1 0 2668 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2492
timestamp 1677677812
transform 1 0 2708 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2522
timestamp 1677677812
transform 1 0 2708 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2914
timestamp 1677677812
transform 1 0 2708 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2585
timestamp 1677677812
transform 1 0 2740 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2493
timestamp 1677677812
transform 1 0 2844 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2523
timestamp 1677677812
transform 1 0 2812 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2524
timestamp 1677677812
transform 1 0 2860 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2915
timestamp 1677677812
transform 1 0 2772 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2562
timestamp 1677677812
transform 1 0 2796 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2916
timestamp 1677677812
transform 1 0 2860 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3011
timestamp 1677677812
transform 1 0 2748 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3012
timestamp 1677677812
transform 1 0 2756 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2586
timestamp 1677677812
transform 1 0 2772 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2494
timestamp 1677677812
transform 1 0 2892 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2917
timestamp 1677677812
transform 1 0 2884 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3013
timestamp 1677677812
transform 1 0 2796 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3014
timestamp 1677677812
transform 1 0 2860 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3015
timestamp 1677677812
transform 1 0 2868 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2620
timestamp 1677677812
transform 1 0 2756 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2621
timestamp 1677677812
transform 1 0 2796 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2622
timestamp 1677677812
transform 1 0 2844 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2623
timestamp 1677677812
transform 1 0 2860 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2650
timestamp 1677677812
transform 1 0 2748 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2651
timestamp 1677677812
transform 1 0 2772 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2652
timestamp 1677677812
transform 1 0 2836 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2653
timestamp 1677677812
transform 1 0 2868 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2918
timestamp 1677677812
transform 1 0 2892 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2587
timestamp 1677677812
transform 1 0 2892 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3016
timestamp 1677677812
transform 1 0 2908 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3061
timestamp 1677677812
transform 1 0 2892 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2919
timestamp 1677677812
transform 1 0 2932 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2588
timestamp 1677677812
transform 1 0 2932 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3062
timestamp 1677677812
transform 1 0 2924 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2654
timestamp 1677677812
transform 1 0 2908 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2655
timestamp 1677677812
transform 1 0 2924 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_3063
timestamp 1677677812
transform 1 0 2932 0 1 3315
box -2 -2 2 2
use M2_M1  M2_M1_2920
timestamp 1677677812
transform 1 0 2996 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2921
timestamp 1677677812
transform 1 0 3004 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3017
timestamp 1677677812
transform 1 0 2988 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2589
timestamp 1677677812
transform 1 0 2996 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3064
timestamp 1677677812
transform 1 0 2972 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2624
timestamp 1677677812
transform 1 0 2988 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2672
timestamp 1677677812
transform 1 0 2972 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3065
timestamp 1677677812
transform 1 0 3012 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2656
timestamp 1677677812
transform 1 0 3004 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2673
timestamp 1677677812
transform 1 0 3012 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3018
timestamp 1677677812
transform 1 0 3076 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2625
timestamp 1677677812
transform 1 0 3076 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2549
timestamp 1677677812
transform 1 0 3132 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2922
timestamp 1677677812
transform 1 0 3124 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2923
timestamp 1677677812
transform 1 0 3132 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2924
timestamp 1677677812
transform 1 0 3148 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3019
timestamp 1677677812
transform 1 0 3132 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3020
timestamp 1677677812
transform 1 0 3156 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2626
timestamp 1677677812
transform 1 0 3124 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2627
timestamp 1677677812
transform 1 0 3156 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2525
timestamp 1677677812
transform 1 0 3172 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2925
timestamp 1677677812
transform 1 0 3172 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3021
timestamp 1677677812
transform 1 0 3172 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2628
timestamp 1677677812
transform 1 0 3172 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2926
timestamp 1677677812
transform 1 0 3220 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2526
timestamp 1677677812
transform 1 0 3244 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2495
timestamp 1677677812
transform 1 0 3276 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2527
timestamp 1677677812
transform 1 0 3300 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2927
timestamp 1677677812
transform 1 0 3284 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2928
timestamp 1677677812
transform 1 0 3300 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3022
timestamp 1677677812
transform 1 0 3268 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3023
timestamp 1677677812
transform 1 0 3276 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2590
timestamp 1677677812
transform 1 0 3284 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3024
timestamp 1677677812
transform 1 0 3292 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3025
timestamp 1677677812
transform 1 0 3308 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2496
timestamp 1677677812
transform 1 0 3316 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2929
timestamp 1677677812
transform 1 0 3324 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3066
timestamp 1677677812
transform 1 0 3380 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2563
timestamp 1677677812
transform 1 0 3412 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3026
timestamp 1677677812
transform 1 0 3404 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2629
timestamp 1677677812
transform 1 0 3404 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2674
timestamp 1677677812
transform 1 0 3388 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_3070
timestamp 1677677812
transform 1 0 3412 0 1 3305
box -2 -2 2 2
use M3_M2  M3_M2_2497
timestamp 1677677812
transform 1 0 3484 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2528
timestamp 1677677812
transform 1 0 3484 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2930
timestamp 1677677812
transform 1 0 3460 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2564
timestamp 1677677812
transform 1 0 3468 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2931
timestamp 1677677812
transform 1 0 3484 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2565
timestamp 1677677812
transform 1 0 3492 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2932
timestamp 1677677812
transform 1 0 3500 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3027
timestamp 1677677812
transform 1 0 3452 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3028
timestamp 1677677812
transform 1 0 3468 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3029
timestamp 1677677812
transform 1 0 3484 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3030
timestamp 1677677812
transform 1 0 3492 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3067
timestamp 1677677812
transform 1 0 3444 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2657
timestamp 1677677812
transform 1 0 3444 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2630
timestamp 1677677812
transform 1 0 3468 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2675
timestamp 1677677812
transform 1 0 3484 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2498
timestamp 1677677812
transform 1 0 3556 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2676
timestamp 1677677812
transform 1 0 3548 0 1 3295
box -3 -3 3 3
use M3_M2  M3_M2_2499
timestamp 1677677812
transform 1 0 3572 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2500
timestamp 1677677812
transform 1 0 3652 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2933
timestamp 1677677812
transform 1 0 3572 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2566
timestamp 1677677812
transform 1 0 3620 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3031
timestamp 1677677812
transform 1 0 3620 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2529
timestamp 1677677812
transform 1 0 3660 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2530
timestamp 1677677812
transform 1 0 3676 0 1 3355
box -3 -3 3 3
use M3_M2  M3_M2_2567
timestamp 1677677812
transform 1 0 3668 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2934
timestamp 1677677812
transform 1 0 3684 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2531
timestamp 1677677812
transform 1 0 3708 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2935
timestamp 1677677812
transform 1 0 3796 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3032
timestamp 1677677812
transform 1 0 3676 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3033
timestamp 1677677812
transform 1 0 3692 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3034
timestamp 1677677812
transform 1 0 3708 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3035
timestamp 1677677812
transform 1 0 3716 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3036
timestamp 1677677812
transform 1 0 3772 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2631
timestamp 1677677812
transform 1 0 3692 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2680
timestamp 1677677812
transform 1 0 3684 0 1 3285
box -3 -3 3 3
use M3_M2  M3_M2_2591
timestamp 1677677812
transform 1 0 3796 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2632
timestamp 1677677812
transform 1 0 3724 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2633
timestamp 1677677812
transform 1 0 3772 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3037
timestamp 1677677812
transform 1 0 3812 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2634
timestamp 1677677812
transform 1 0 3812 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2936
timestamp 1677677812
transform 1 0 3860 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2568
timestamp 1677677812
transform 1 0 3868 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2937
timestamp 1677677812
transform 1 0 3884 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3038
timestamp 1677677812
transform 1 0 3852 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3039
timestamp 1677677812
transform 1 0 3868 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3040
timestamp 1677677812
transform 1 0 3884 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2658
timestamp 1677677812
transform 1 0 3868 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2501
timestamp 1677677812
transform 1 0 3908 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2569
timestamp 1677677812
transform 1 0 3900 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3041
timestamp 1677677812
transform 1 0 3900 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2592
timestamp 1677677812
transform 1 0 3908 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2635
timestamp 1677677812
transform 1 0 3916 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_2938
timestamp 1677677812
transform 1 0 3948 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2502
timestamp 1677677812
transform 1 0 4036 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2939
timestamp 1677677812
transform 1 0 4036 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3042
timestamp 1677677812
transform 1 0 3956 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3043
timestamp 1677677812
transform 1 0 4012 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2593
timestamp 1677677812
transform 1 0 4036 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2503
timestamp 1677677812
transform 1 0 4060 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2532
timestamp 1677677812
transform 1 0 4052 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2940
timestamp 1677677812
transform 1 0 4092 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2504
timestamp 1677677812
transform 1 0 4196 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2941
timestamp 1677677812
transform 1 0 4188 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3044
timestamp 1677677812
transform 1 0 4116 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3045
timestamp 1677677812
transform 1 0 4172 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3046
timestamp 1677677812
transform 1 0 4180 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3047
timestamp 1677677812
transform 1 0 4244 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2505
timestamp 1677677812
transform 1 0 4276 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2533
timestamp 1677677812
transform 1 0 4260 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2942
timestamp 1677677812
transform 1 0 4260 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2943
timestamp 1677677812
transform 1 0 4284 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2570
timestamp 1677677812
transform 1 0 4292 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3048
timestamp 1677677812
transform 1 0 4276 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3049
timestamp 1677677812
transform 1 0 4292 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2677
timestamp 1677677812
transform 1 0 4276 0 1 3295
box -3 -3 3 3
use M2_M1  M2_M1_2944
timestamp 1677677812
transform 1 0 4316 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2550
timestamp 1677677812
transform 1 0 4340 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2945
timestamp 1677677812
transform 1 0 4340 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3068
timestamp 1677677812
transform 1 0 4324 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2636
timestamp 1677677812
transform 1 0 4348 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3071
timestamp 1677677812
transform 1 0 4332 0 1 3305
box -2 -2 2 2
use M3_M2  M3_M2_2506
timestamp 1677677812
transform 1 0 4372 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2946
timestamp 1677677812
transform 1 0 4372 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3069
timestamp 1677677812
transform 1 0 4364 0 1 3315
box -2 -2 2 2
use M3_M2  M3_M2_2659
timestamp 1677677812
transform 1 0 4372 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2947
timestamp 1677677812
transform 1 0 4404 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2571
timestamp 1677677812
transform 1 0 4412 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_2948
timestamp 1677677812
transform 1 0 4420 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3050
timestamp 1677677812
transform 1 0 4396 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2594
timestamp 1677677812
transform 1 0 4404 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3051
timestamp 1677677812
transform 1 0 4412 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3052
timestamp 1677677812
transform 1 0 4452 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2660
timestamp 1677677812
transform 1 0 4444 0 1 3305
box -3 -3 3 3
use M3_M2  M3_M2_2551
timestamp 1677677812
transform 1 0 4476 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2572
timestamp 1677677812
transform 1 0 4484 0 1 3335
box -3 -3 3 3
use M2_M1  M2_M1_3053
timestamp 1677677812
transform 1 0 4484 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2552
timestamp 1677677812
transform 1 0 4500 0 1 3345
box -3 -3 3 3
use M2_M1  M2_M1_2949
timestamp 1677677812
transform 1 0 4500 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2637
timestamp 1677677812
transform 1 0 4492 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2595
timestamp 1677677812
transform 1 0 4516 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2507
timestamp 1677677812
transform 1 0 4532 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2553
timestamp 1677677812
transform 1 0 4540 0 1 3345
box -3 -3 3 3
use M3_M2  M3_M2_2638
timestamp 1677677812
transform 1 0 4532 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2508
timestamp 1677677812
transform 1 0 4556 0 1 3365
box -3 -3 3 3
use M3_M2  M3_M2_2534
timestamp 1677677812
transform 1 0 4580 0 1 3355
box -3 -3 3 3
use M2_M1  M2_M1_2950
timestamp 1677677812
transform 1 0 4548 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2951
timestamp 1677677812
transform 1 0 4556 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_2952
timestamp 1677677812
transform 1 0 4572 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2596
timestamp 1677677812
transform 1 0 4548 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3054
timestamp 1677677812
transform 1 0 4564 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2597
timestamp 1677677812
transform 1 0 4572 0 1 3325
box -3 -3 3 3
use M2_M1  M2_M1_3055
timestamp 1677677812
transform 1 0 4580 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2639
timestamp 1677677812
transform 1 0 4564 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2640
timestamp 1677677812
transform 1 0 4580 0 1 3315
box -3 -3 3 3
use M2_M1  M2_M1_3056
timestamp 1677677812
transform 1 0 4596 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2661
timestamp 1677677812
transform 1 0 4588 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2953
timestamp 1677677812
transform 1 0 4612 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2598
timestamp 1677677812
transform 1 0 4612 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2662
timestamp 1677677812
transform 1 0 4620 0 1 3305
box -3 -3 3 3
use M2_M1  M2_M1_2954
timestamp 1677677812
transform 1 0 4636 0 1 3335
box -2 -2 2 2
use M3_M2  M3_M2_2599
timestamp 1677677812
transform 1 0 4636 0 1 3325
box -3 -3 3 3
use M3_M2  M3_M2_2509
timestamp 1677677812
transform 1 0 4660 0 1 3365
box -3 -3 3 3
use M2_M1  M2_M1_2955
timestamp 1677677812
transform 1 0 4708 0 1 3335
box -2 -2 2 2
use M2_M1  M2_M1_3057
timestamp 1677677812
transform 1 0 4740 0 1 3325
box -2 -2 2 2
use M2_M1  M2_M1_3058
timestamp 1677677812
transform 1 0 4788 0 1 3325
box -2 -2 2 2
use M3_M2  M3_M2_2641
timestamp 1677677812
transform 1 0 4748 0 1 3315
box -3 -3 3 3
use M3_M2  M3_M2_2642
timestamp 1677677812
transform 1 0 4788 0 1 3315
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_28
timestamp 1677677812
transform 1 0 24 0 1 3270
box -10 -3 10 3
use FILL  FILL_2740
timestamp 1677677812
transform 1 0 72 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2746
timestamp 1677677812
transform 1 0 80 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2747
timestamp 1677677812
transform 1 0 88 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_187
timestamp 1677677812
transform -1 0 192 0 -1 3370
box -8 -3 104 105
use INVX2  INVX2_216
timestamp 1677677812
transform -1 0 208 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2748
timestamp 1677677812
transform 1 0 208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2751
timestamp 1677677812
transform 1 0 216 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_124
timestamp 1677677812
transform 1 0 224 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2752
timestamp 1677677812
transform 1 0 264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2754
timestamp 1677677812
transform 1 0 272 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2759
timestamp 1677677812
transform 1 0 280 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2760
timestamp 1677677812
transform 1 0 288 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_120
timestamp 1677677812
transform -1 0 336 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2761
timestamp 1677677812
transform 1 0 336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2762
timestamp 1677677812
transform 1 0 344 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2763
timestamp 1677677812
transform 1 0 352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2764
timestamp 1677677812
transform 1 0 360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2765
timestamp 1677677812
transform 1 0 368 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_125
timestamp 1677677812
transform -1 0 416 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2766
timestamp 1677677812
transform 1 0 416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2768
timestamp 1677677812
transform 1 0 424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2774
timestamp 1677677812
transform 1 0 432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2775
timestamp 1677677812
transform 1 0 440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2776
timestamp 1677677812
transform 1 0 448 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2777
timestamp 1677677812
transform 1 0 456 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2778
timestamp 1677677812
transform 1 0 464 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_126
timestamp 1677677812
transform 1 0 472 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2779
timestamp 1677677812
transform 1 0 512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2780
timestamp 1677677812
transform 1 0 520 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2681
timestamp 1677677812
transform 1 0 540 0 1 3275
box -3 -3 3 3
use FILL  FILL_2782
timestamp 1677677812
transform 1 0 528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2784
timestamp 1677677812
transform 1 0 536 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2787
timestamp 1677677812
transform 1 0 544 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_190
timestamp 1677677812
transform 1 0 552 0 -1 3370
box -8 -3 104 105
use M3_M2  M3_M2_2682
timestamp 1677677812
transform 1 0 660 0 1 3275
box -3 -3 3 3
use FILL  FILL_2788
timestamp 1677677812
transform 1 0 648 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2789
timestamp 1677677812
transform 1 0 656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2790
timestamp 1677677812
transform 1 0 664 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2791
timestamp 1677677812
transform 1 0 672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2793
timestamp 1677677812
transform 1 0 680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2795
timestamp 1677677812
transform 1 0 688 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_122
timestamp 1677677812
transform 1 0 696 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2799
timestamp 1677677812
transform 1 0 736 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2801
timestamp 1677677812
transform 1 0 744 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2803
timestamp 1677677812
transform 1 0 752 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2805
timestamp 1677677812
transform 1 0 760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2819
timestamp 1677677812
transform 1 0 768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2820
timestamp 1677677812
transform 1 0 776 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2821
timestamp 1677677812
transform 1 0 784 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2822
timestamp 1677677812
transform 1 0 792 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_219
timestamp 1677677812
transform 1 0 800 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2823
timestamp 1677677812
transform 1 0 816 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2824
timestamp 1677677812
transform 1 0 824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2825
timestamp 1677677812
transform 1 0 832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2826
timestamp 1677677812
transform 1 0 840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2827
timestamp 1677677812
transform 1 0 848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2828
timestamp 1677677812
transform 1 0 856 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_192
timestamp 1677677812
transform 1 0 864 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2829
timestamp 1677677812
transform 1 0 960 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2832
timestamp 1677677812
transform 1 0 968 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2833
timestamp 1677677812
transform 1 0 976 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_220
timestamp 1677677812
transform -1 0 1000 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2834
timestamp 1677677812
transform 1 0 1000 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2836
timestamp 1677677812
transform 1 0 1008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2838
timestamp 1677677812
transform 1 0 1016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2840
timestamp 1677677812
transform 1 0 1024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2842
timestamp 1677677812
transform 1 0 1032 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2844
timestamp 1677677812
transform 1 0 1040 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_127
timestamp 1677677812
transform 1 0 1048 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2847
timestamp 1677677812
transform 1 0 1088 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2849
timestamp 1677677812
transform 1 0 1096 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2851
timestamp 1677677812
transform 1 0 1104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2853
timestamp 1677677812
transform 1 0 1112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2855
timestamp 1677677812
transform 1 0 1120 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2858
timestamp 1677677812
transform 1 0 1128 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2859
timestamp 1677677812
transform 1 0 1136 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_63
timestamp 1677677812
transform 1 0 1144 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2860
timestamp 1677677812
transform 1 0 1176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2862
timestamp 1677677812
transform 1 0 1184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2864
timestamp 1677677812
transform 1 0 1192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2866
timestamp 1677677812
transform 1 0 1200 0 -1 3370
box -8 -3 16 105
use NOR2X1  NOR2X1_30
timestamp 1677677812
transform 1 0 1208 0 -1 3370
box -8 -3 32 105
use FILL  FILL_2870
timestamp 1677677812
transform 1 0 1232 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2871
timestamp 1677677812
transform 1 0 1240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2872
timestamp 1677677812
transform 1 0 1248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2873
timestamp 1677677812
transform 1 0 1256 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2874
timestamp 1677677812
transform 1 0 1264 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_64
timestamp 1677677812
transform 1 0 1272 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2875
timestamp 1677677812
transform 1 0 1304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2876
timestamp 1677677812
transform 1 0 1312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2877
timestamp 1677677812
transform 1 0 1320 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2878
timestamp 1677677812
transform 1 0 1328 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2879
timestamp 1677677812
transform 1 0 1336 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2883
timestamp 1677677812
transform 1 0 1344 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_65
timestamp 1677677812
transform -1 0 1384 0 -1 3370
box -8 -3 34 105
use FILL  FILL_2884
timestamp 1677677812
transform 1 0 1384 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2887
timestamp 1677677812
transform 1 0 1392 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2888
timestamp 1677677812
transform 1 0 1400 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2889
timestamp 1677677812
transform 1 0 1408 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2890
timestamp 1677677812
transform 1 0 1416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2891
timestamp 1677677812
transform 1 0 1424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2892
timestamp 1677677812
transform 1 0 1432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2893
timestamp 1677677812
transform 1 0 1440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2894
timestamp 1677677812
transform 1 0 1448 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_123
timestamp 1677677812
transform 1 0 1456 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2895
timestamp 1677677812
transform 1 0 1496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2896
timestamp 1677677812
transform 1 0 1504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2897
timestamp 1677677812
transform 1 0 1512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2898
timestamp 1677677812
transform 1 0 1520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2899
timestamp 1677677812
transform 1 0 1528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2900
timestamp 1677677812
transform 1 0 1536 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_223
timestamp 1677677812
transform 1 0 1544 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2901
timestamp 1677677812
transform 1 0 1560 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2902
timestamp 1677677812
transform 1 0 1568 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2903
timestamp 1677677812
transform 1 0 1576 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2904
timestamp 1677677812
transform 1 0 1584 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2905
timestamp 1677677812
transform 1 0 1592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2906
timestamp 1677677812
transform 1 0 1600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2907
timestamp 1677677812
transform 1 0 1608 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2916
timestamp 1677677812
transform 1 0 1616 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_124
timestamp 1677677812
transform -1 0 1664 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2917
timestamp 1677677812
transform 1 0 1664 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2918
timestamp 1677677812
transform 1 0 1672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2919
timestamp 1677677812
transform 1 0 1680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2920
timestamp 1677677812
transform 1 0 1688 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2921
timestamp 1677677812
transform 1 0 1696 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2922
timestamp 1677677812
transform 1 0 1704 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2923
timestamp 1677677812
transform 1 0 1712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2924
timestamp 1677677812
transform 1 0 1720 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2683
timestamp 1677677812
transform 1 0 1748 0 1 3275
box -3 -3 3 3
use BUFX2  BUFX2_19
timestamp 1677677812
transform 1 0 1728 0 -1 3370
box -5 -3 28 105
use FILL  FILL_2925
timestamp 1677677812
transform 1 0 1752 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2926
timestamp 1677677812
transform 1 0 1760 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2927
timestamp 1677677812
transform 1 0 1768 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2928
timestamp 1677677812
transform 1 0 1776 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_125
timestamp 1677677812
transform -1 0 1824 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2929
timestamp 1677677812
transform 1 0 1824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2930
timestamp 1677677812
transform 1 0 1832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2931
timestamp 1677677812
transform 1 0 1840 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2932
timestamp 1677677812
transform 1 0 1848 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2933
timestamp 1677677812
transform 1 0 1856 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_225
timestamp 1677677812
transform -1 0 1880 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2934
timestamp 1677677812
transform 1 0 1880 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2935
timestamp 1677677812
transform 1 0 1888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2936
timestamp 1677677812
transform 1 0 1896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2937
timestamp 1677677812
transform 1 0 1904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2947
timestamp 1677677812
transform 1 0 1912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2948
timestamp 1677677812
transform 1 0 1920 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2949
timestamp 1677677812
transform 1 0 1928 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2950
timestamp 1677677812
transform 1 0 1936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2951
timestamp 1677677812
transform 1 0 1944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2952
timestamp 1677677812
transform 1 0 1952 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_201
timestamp 1677677812
transform 1 0 1960 0 -1 3370
box -8 -3 104 105
use FILL  FILL_2953
timestamp 1677677812
transform 1 0 2056 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2684
timestamp 1677677812
transform 1 0 2076 0 1 3275
box -3 -3 3 3
use FILL  FILL_2954
timestamp 1677677812
transform 1 0 2064 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2955
timestamp 1677677812
transform 1 0 2072 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2956
timestamp 1677677812
transform 1 0 2080 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2957
timestamp 1677677812
transform 1 0 2088 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2958
timestamp 1677677812
transform 1 0 2096 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2959
timestamp 1677677812
transform 1 0 2104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2960
timestamp 1677677812
transform 1 0 2112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2961
timestamp 1677677812
transform 1 0 2120 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2962
timestamp 1677677812
transform 1 0 2128 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2963
timestamp 1677677812
transform 1 0 2136 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2964
timestamp 1677677812
transform 1 0 2144 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_129
timestamp 1677677812
transform -1 0 2192 0 -1 3370
box -8 -3 46 105
use FILL  FILL_2965
timestamp 1677677812
transform 1 0 2192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2966
timestamp 1677677812
transform 1 0 2200 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2685
timestamp 1677677812
transform 1 0 2220 0 1 3275
box -3 -3 3 3
use FILL  FILL_2967
timestamp 1677677812
transform 1 0 2208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2968
timestamp 1677677812
transform 1 0 2216 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_130
timestamp 1677677812
transform 1 0 2224 0 -1 3370
box -8 -3 46 105
use M3_M2  M3_M2_2686
timestamp 1677677812
transform 1 0 2284 0 1 3275
box -3 -3 3 3
use FILL  FILL_2969
timestamp 1677677812
transform 1 0 2264 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2970
timestamp 1677677812
transform 1 0 2272 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_228
timestamp 1677677812
transform 1 0 2280 0 -1 3370
box -9 -3 26 105
use FILL  FILL_2971
timestamp 1677677812
transform 1 0 2296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2973
timestamp 1677677812
transform 1 0 2304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2975
timestamp 1677677812
transform 1 0 2312 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_202
timestamp 1677677812
transform 1 0 2320 0 -1 3370
box -8 -3 104 105
use M3_M2  M3_M2_2687
timestamp 1677677812
transform 1 0 2428 0 1 3275
box -3 -3 3 3
use FILL  FILL_2980
timestamp 1677677812
transform 1 0 2416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2982
timestamp 1677677812
transform 1 0 2424 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2688
timestamp 1677677812
transform 1 0 2444 0 1 3275
box -3 -3 3 3
use FILL  FILL_2984
timestamp 1677677812
transform 1 0 2432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2986
timestamp 1677677812
transform 1 0 2440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2988
timestamp 1677677812
transform 1 0 2448 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2990
timestamp 1677677812
transform 1 0 2456 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2991
timestamp 1677677812
transform 1 0 2464 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2992
timestamp 1677677812
transform 1 0 2472 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2993
timestamp 1677677812
transform 1 0 2480 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2995
timestamp 1677677812
transform 1 0 2488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2997
timestamp 1677677812
transform 1 0 2496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_2999
timestamp 1677677812
transform 1 0 2504 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3011
timestamp 1677677812
transform 1 0 2512 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3012
timestamp 1677677812
transform 1 0 2520 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_230
timestamp 1677677812
transform 1 0 2528 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3013
timestamp 1677677812
transform 1 0 2544 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_203
timestamp 1677677812
transform -1 0 2648 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3014
timestamp 1677677812
transform 1 0 2648 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3028
timestamp 1677677812
transform 1 0 2656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3029
timestamp 1677677812
transform 1 0 2664 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3030
timestamp 1677677812
transform 1 0 2672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3031
timestamp 1677677812
transform 1 0 2680 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_231
timestamp 1677677812
transform 1 0 2688 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3032
timestamp 1677677812
transform 1 0 2704 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3033
timestamp 1677677812
transform 1 0 2712 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3034
timestamp 1677677812
transform 1 0 2720 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3035
timestamp 1677677812
transform 1 0 2728 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3036
timestamp 1677677812
transform 1 0 2736 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_232
timestamp 1677677812
transform 1 0 2744 0 -1 3370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_204
timestamp 1677677812
transform 1 0 2760 0 -1 3370
box -8 -3 104 105
use OAI21X1  OAI21X1_67
timestamp 1677677812
transform 1 0 2856 0 -1 3370
box -8 -3 34 105
use FILL  FILL_3038
timestamp 1677677812
transform 1 0 2888 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_68
timestamp 1677677812
transform 1 0 2896 0 -1 3370
box -8 -3 34 105
use FILL  FILL_3044
timestamp 1677677812
transform 1 0 2928 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3050
timestamp 1677677812
transform 1 0 2936 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3051
timestamp 1677677812
transform 1 0 2944 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3052
timestamp 1677677812
transform 1 0 2952 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3053
timestamp 1677677812
transform 1 0 2960 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_69
timestamp 1677677812
transform -1 0 3000 0 -1 3370
box -8 -3 34 105
use FILL  FILL_3054
timestamp 1677677812
transform 1 0 3000 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2689
timestamp 1677677812
transform 1 0 3020 0 1 3275
box -3 -3 3 3
use FILL  FILL_3056
timestamp 1677677812
transform 1 0 3008 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3057
timestamp 1677677812
transform 1 0 3016 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3058
timestamp 1677677812
transform 1 0 3024 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3059
timestamp 1677677812
transform 1 0 3032 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3060
timestamp 1677677812
transform 1 0 3040 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3061
timestamp 1677677812
transform 1 0 3048 0 -1 3370
box -8 -3 16 105
use OAI21X1  OAI21X1_70
timestamp 1677677812
transform -1 0 3088 0 -1 3370
box -8 -3 34 105
use FILL  FILL_3062
timestamp 1677677812
transform 1 0 3088 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3063
timestamp 1677677812
transform 1 0 3096 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3064
timestamp 1677677812
transform 1 0 3104 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3066
timestamp 1677677812
transform 1 0 3112 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3068
timestamp 1677677812
transform 1 0 3120 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_127
timestamp 1677677812
transform 1 0 3128 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3070
timestamp 1677677812
transform 1 0 3168 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3071
timestamp 1677677812
transform 1 0 3176 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3072
timestamp 1677677812
transform 1 0 3184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3073
timestamp 1677677812
transform 1 0 3192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3074
timestamp 1677677812
transform 1 0 3200 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_233
timestamp 1677677812
transform -1 0 3224 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3075
timestamp 1677677812
transform 1 0 3224 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3078
timestamp 1677677812
transform 1 0 3232 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3079
timestamp 1677677812
transform 1 0 3240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3080
timestamp 1677677812
transform 1 0 3248 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3081
timestamp 1677677812
transform 1 0 3256 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_128
timestamp 1677677812
transform 1 0 3264 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3082
timestamp 1677677812
transform 1 0 3304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3083
timestamp 1677677812
transform 1 0 3312 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3084
timestamp 1677677812
transform 1 0 3320 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_234
timestamp 1677677812
transform 1 0 3328 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3085
timestamp 1677677812
transform 1 0 3344 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3086
timestamp 1677677812
transform 1 0 3352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3087
timestamp 1677677812
transform 1 0 3360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3088
timestamp 1677677812
transform 1 0 3368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3093
timestamp 1677677812
transform 1 0 3376 0 -1 3370
box -8 -3 16 105
use NAND3X1  NAND3X1_14
timestamp 1677677812
transform -1 0 3416 0 -1 3370
box -8 -3 40 105
use FILL  FILL_3094
timestamp 1677677812
transform 1 0 3416 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3095
timestamp 1677677812
transform 1 0 3424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3096
timestamp 1677677812
transform 1 0 3432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3097
timestamp 1677677812
transform 1 0 3440 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_133
timestamp 1677677812
transform 1 0 3448 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3098
timestamp 1677677812
transform 1 0 3488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3099
timestamp 1677677812
transform 1 0 3496 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3101
timestamp 1677677812
transform 1 0 3504 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_235
timestamp 1677677812
transform 1 0 3512 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3126
timestamp 1677677812
transform 1 0 3528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3127
timestamp 1677677812
transform 1 0 3536 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3128
timestamp 1677677812
transform 1 0 3544 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3129
timestamp 1677677812
transform 1 0 3552 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2690
timestamp 1677677812
transform 1 0 3572 0 1 3275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_209
timestamp 1677677812
transform 1 0 3560 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3130
timestamp 1677677812
transform 1 0 3656 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_236
timestamp 1677677812
transform 1 0 3664 0 -1 3370
box -9 -3 26 105
use AND2X2  AND2X2_10
timestamp 1677677812
transform 1 0 3680 0 -1 3370
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_210
timestamp 1677677812
transform -1 0 3808 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3131
timestamp 1677677812
transform 1 0 3808 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3133
timestamp 1677677812
transform 1 0 3816 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3135
timestamp 1677677812
transform 1 0 3824 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3139
timestamp 1677677812
transform 1 0 3832 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3140
timestamp 1677677812
transform 1 0 3840 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_134
timestamp 1677677812
transform -1 0 3888 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3141
timestamp 1677677812
transform 1 0 3888 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3146
timestamp 1677677812
transform 1 0 3896 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3147
timestamp 1677677812
transform 1 0 3904 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3148
timestamp 1677677812
transform 1 0 3912 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3149
timestamp 1677677812
transform 1 0 3920 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_237
timestamp 1677677812
transform -1 0 3944 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3150
timestamp 1677677812
transform 1 0 3944 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_212
timestamp 1677677812
transform -1 0 4048 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3151
timestamp 1677677812
transform 1 0 4048 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3152
timestamp 1677677812
transform 1 0 4056 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3154
timestamp 1677677812
transform 1 0 4064 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3156
timestamp 1677677812
transform 1 0 4072 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_214
timestamp 1677677812
transform 1 0 4080 0 -1 3370
box -8 -3 104 105
use FILL  FILL_3159
timestamp 1677677812
transform 1 0 4176 0 -1 3370
box -8 -3 16 105
use M3_M2  M3_M2_2691
timestamp 1677677812
transform 1 0 4196 0 1 3275
box -3 -3 3 3
use FILL  FILL_3160
timestamp 1677677812
transform 1 0 4184 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3162
timestamp 1677677812
transform 1 0 4192 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3164
timestamp 1677677812
transform 1 0 4200 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3179
timestamp 1677677812
transform 1 0 4208 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3180
timestamp 1677677812
transform 1 0 4216 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_239
timestamp 1677677812
transform 1 0 4224 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3181
timestamp 1677677812
transform 1 0 4240 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3182
timestamp 1677677812
transform 1 0 4248 0 -1 3370
box -8 -3 16 105
use AOI22X1  AOI22X1_136
timestamp 1677677812
transform -1 0 4296 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3183
timestamp 1677677812
transform 1 0 4296 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3184
timestamp 1677677812
transform 1 0 4304 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3185
timestamp 1677677812
transform 1 0 4312 0 -1 3370
box -8 -3 16 105
use NAND3X1  NAND3X1_15
timestamp 1677677812
transform -1 0 4352 0 -1 3370
box -8 -3 40 105
use FILL  FILL_3186
timestamp 1677677812
transform 1 0 4352 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3187
timestamp 1677677812
transform 1 0 4360 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3188
timestamp 1677677812
transform 1 0 4368 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3189
timestamp 1677677812
transform 1 0 4376 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_134
timestamp 1677677812
transform 1 0 4384 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3190
timestamp 1677677812
transform 1 0 4424 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3191
timestamp 1677677812
transform 1 0 4432 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3193
timestamp 1677677812
transform 1 0 4440 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3195
timestamp 1677677812
transform 1 0 4448 0 -1 3370
box -8 -3 16 105
use BUFX2  BUFX2_21
timestamp 1677677812
transform 1 0 4456 0 -1 3370
box -5 -3 28 105
use FILL  FILL_3200
timestamp 1677677812
transform 1 0 4480 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3201
timestamp 1677677812
transform 1 0 4488 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3202
timestamp 1677677812
transform 1 0 4496 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_240
timestamp 1677677812
transform -1 0 4520 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3203
timestamp 1677677812
transform 1 0 4520 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3205
timestamp 1677677812
transform 1 0 4528 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3207
timestamp 1677677812
transform 1 0 4536 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3209
timestamp 1677677812
transform 1 0 4544 0 -1 3370
box -8 -3 16 105
use OAI22X1  OAI22X1_135
timestamp 1677677812
transform 1 0 4552 0 -1 3370
box -8 -3 46 105
use FILL  FILL_3210
timestamp 1677677812
transform 1 0 4592 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3211
timestamp 1677677812
transform 1 0 4600 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3212
timestamp 1677677812
transform 1 0 4608 0 -1 3370
box -8 -3 16 105
use INVX2  INVX2_242
timestamp 1677677812
transform -1 0 4632 0 -1 3370
box -9 -3 26 105
use FILL  FILL_3213
timestamp 1677677812
transform 1 0 4632 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3214
timestamp 1677677812
transform 1 0 4640 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3215
timestamp 1677677812
transform 1 0 4648 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3216
timestamp 1677677812
transform 1 0 4656 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3226
timestamp 1677677812
transform 1 0 4664 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3227
timestamp 1677677812
transform 1 0 4672 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3228
timestamp 1677677812
transform 1 0 4680 0 -1 3370
box -8 -3 16 105
use FILL  FILL_3229
timestamp 1677677812
transform 1 0 4688 0 -1 3370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_216
timestamp 1677677812
transform 1 0 4696 0 -1 3370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_29
timestamp 1677677812
transform 1 0 4843 0 1 3270
box -10 -3 10 3
use M3_M2  M3_M2_2733
timestamp 1677677812
transform 1 0 148 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2775
timestamp 1677677812
transform 1 0 4 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2714
timestamp 1677677812
transform 1 0 212 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2734
timestamp 1677677812
transform 1 0 180 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2747
timestamp 1677677812
transform 1 0 164 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3089
timestamp 1677677812
transform 1 0 132 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3090
timestamp 1677677812
transform 1 0 164 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3091
timestamp 1677677812
transform 1 0 172 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3190
timestamp 1677677812
transform 1 0 84 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2802
timestamp 1677677812
transform 1 0 132 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2844
timestamp 1677677812
transform 1 0 148 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2748
timestamp 1677677812
transform 1 0 196 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3092
timestamp 1677677812
transform 1 0 180 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3093
timestamp 1677677812
transform 1 0 204 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2776
timestamp 1677677812
transform 1 0 212 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2701
timestamp 1677677812
transform 1 0 228 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2715
timestamp 1677677812
transform 1 0 228 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3094
timestamp 1677677812
transform 1 0 220 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2803
timestamp 1677677812
transform 1 0 180 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3191
timestamp 1677677812
transform 1 0 188 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3192
timestamp 1677677812
transform 1 0 196 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3193
timestamp 1677677812
transform 1 0 220 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2817
timestamp 1677677812
transform 1 0 188 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2818
timestamp 1677677812
transform 1 0 212 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2845
timestamp 1677677812
transform 1 0 188 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3194
timestamp 1677677812
transform 1 0 252 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2819
timestamp 1677677812
transform 1 0 252 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2735
timestamp 1677677812
transform 1 0 268 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2749
timestamp 1677677812
transform 1 0 268 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2702
timestamp 1677677812
transform 1 0 364 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2716
timestamp 1677677812
transform 1 0 308 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2750
timestamp 1677677812
transform 1 0 308 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3095
timestamp 1677677812
transform 1 0 268 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3096
timestamp 1677677812
transform 1 0 276 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3097
timestamp 1677677812
transform 1 0 308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3195
timestamp 1677677812
transform 1 0 356 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2820
timestamp 1677677812
transform 1 0 292 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2821
timestamp 1677677812
transform 1 0 324 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2717
timestamp 1677677812
transform 1 0 404 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3098
timestamp 1677677812
transform 1 0 420 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3099
timestamp 1677677812
transform 1 0 468 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3196
timestamp 1677677812
transform 1 0 388 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2751
timestamp 1677677812
transform 1 0 508 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3197
timestamp 1677677812
transform 1 0 508 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2718
timestamp 1677677812
transform 1 0 556 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2736
timestamp 1677677812
transform 1 0 548 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3100
timestamp 1677677812
transform 1 0 548 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3198
timestamp 1677677812
transform 1 0 548 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2737
timestamp 1677677812
transform 1 0 604 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2752
timestamp 1677677812
transform 1 0 580 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2753
timestamp 1677677812
transform 1 0 596 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3101
timestamp 1677677812
transform 1 0 564 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2777
timestamp 1677677812
transform 1 0 572 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3102
timestamp 1677677812
transform 1 0 580 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3103
timestamp 1677677812
transform 1 0 596 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3199
timestamp 1677677812
transform 1 0 572 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3200
timestamp 1677677812
transform 1 0 588 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3201
timestamp 1677677812
transform 1 0 612 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3297
timestamp 1677677812
transform 1 0 620 0 1 3185
box -2 -2 2 2
use M3_M2  M3_M2_2778
timestamp 1677677812
transform 1 0 644 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3202
timestamp 1677677812
transform 1 0 644 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3104
timestamp 1677677812
transform 1 0 660 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3105
timestamp 1677677812
transform 1 0 676 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3203
timestamp 1677677812
transform 1 0 668 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3204
timestamp 1677677812
transform 1 0 684 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2703
timestamp 1677677812
transform 1 0 708 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3106
timestamp 1677677812
transform 1 0 708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3107
timestamp 1677677812
transform 1 0 788 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3205
timestamp 1677677812
transform 1 0 772 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3108
timestamp 1677677812
transform 1 0 828 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3291
timestamp 1677677812
transform 1 0 820 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3109
timestamp 1677677812
transform 1 0 852 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3206
timestamp 1677677812
transform 1 0 868 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2779
timestamp 1677677812
transform 1 0 884 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3110
timestamp 1677677812
transform 1 0 892 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3207
timestamp 1677677812
transform 1 0 892 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3208
timestamp 1677677812
transform 1 0 908 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3111
timestamp 1677677812
transform 1 0 924 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2780
timestamp 1677677812
transform 1 0 964 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3209
timestamp 1677677812
transform 1 0 964 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2754
timestamp 1677677812
transform 1 0 996 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3076
timestamp 1677677812
transform 1 0 1004 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2781
timestamp 1677677812
transform 1 0 1004 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3292
timestamp 1677677812
transform 1 0 996 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2738
timestamp 1677677812
transform 1 0 1028 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2704
timestamp 1677677812
transform 1 0 1052 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2755
timestamp 1677677812
transform 1 0 1052 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3293
timestamp 1677677812
transform 1 0 1044 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2705
timestamp 1677677812
transform 1 0 1076 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2756
timestamp 1677677812
transform 1 0 1068 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3112
timestamp 1677677812
transform 1 0 1068 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3294
timestamp 1677677812
transform 1 0 1068 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2739
timestamp 1677677812
transform 1 0 1084 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2740
timestamp 1677677812
transform 1 0 1100 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3113
timestamp 1677677812
transform 1 0 1092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3114
timestamp 1677677812
transform 1 0 1108 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3210
timestamp 1677677812
transform 1 0 1084 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3211
timestamp 1677677812
transform 1 0 1116 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2757
timestamp 1677677812
transform 1 0 1172 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3115
timestamp 1677677812
transform 1 0 1164 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3212
timestamp 1677677812
transform 1 0 1164 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3116
timestamp 1677677812
transform 1 0 1188 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3117
timestamp 1677677812
transform 1 0 1212 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3213
timestamp 1677677812
transform 1 0 1204 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2782
timestamp 1677677812
transform 1 0 1228 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3214
timestamp 1677677812
transform 1 0 1228 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3077
timestamp 1677677812
transform 1 0 1252 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2783
timestamp 1677677812
transform 1 0 1260 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2719
timestamp 1677677812
transform 1 0 1284 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3118
timestamp 1677677812
transform 1 0 1276 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3215
timestamp 1677677812
transform 1 0 1284 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3078
timestamp 1677677812
transform 1 0 1308 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2784
timestamp 1677677812
transform 1 0 1308 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3216
timestamp 1677677812
transform 1 0 1324 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3119
timestamp 1677677812
transform 1 0 1364 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3120
timestamp 1677677812
transform 1 0 1380 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3121
timestamp 1677677812
transform 1 0 1436 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3122
timestamp 1677677812
transform 1 0 1460 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3217
timestamp 1677677812
transform 1 0 1420 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3218
timestamp 1677677812
transform 1 0 1428 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3219
timestamp 1677677812
transform 1 0 1444 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2846
timestamp 1677677812
transform 1 0 1420 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2822
timestamp 1677677812
transform 1 0 1468 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2720
timestamp 1677677812
transform 1 0 1484 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3123
timestamp 1677677812
transform 1 0 1556 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3124
timestamp 1677677812
transform 1 0 1580 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3220
timestamp 1677677812
transform 1 0 1540 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3221
timestamp 1677677812
transform 1 0 1548 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3222
timestamp 1677677812
transform 1 0 1564 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3223
timestamp 1677677812
transform 1 0 1580 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3224
timestamp 1677677812
transform 1 0 1588 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2847
timestamp 1677677812
transform 1 0 1556 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2848
timestamp 1677677812
transform 1 0 1580 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3125
timestamp 1677677812
transform 1 0 1604 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2849
timestamp 1677677812
transform 1 0 1620 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2706
timestamp 1677677812
transform 1 0 1692 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3225
timestamp 1677677812
transform 1 0 1692 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2850
timestamp 1677677812
transform 1 0 1692 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2721
timestamp 1677677812
transform 1 0 1724 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3126
timestamp 1677677812
transform 1 0 1716 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3127
timestamp 1677677812
transform 1 0 1724 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2851
timestamp 1677677812
transform 1 0 1708 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3226
timestamp 1677677812
transform 1 0 1748 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2722
timestamp 1677677812
transform 1 0 1772 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3128
timestamp 1677677812
transform 1 0 1772 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2707
timestamp 1677677812
transform 1 0 1796 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2723
timestamp 1677677812
transform 1 0 1788 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3129
timestamp 1677677812
transform 1 0 1796 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2785
timestamp 1677677812
transform 1 0 1812 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3227
timestamp 1677677812
transform 1 0 1812 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2852
timestamp 1677677812
transform 1 0 1820 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3130
timestamp 1677677812
transform 1 0 1844 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2708
timestamp 1677677812
transform 1 0 1868 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2786
timestamp 1677677812
transform 1 0 1860 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2724
timestamp 1677677812
transform 1 0 1884 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3228
timestamp 1677677812
transform 1 0 1876 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3229
timestamp 1677677812
transform 1 0 1884 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2709
timestamp 1677677812
transform 1 0 1892 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2787
timestamp 1677677812
transform 1 0 1892 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3131
timestamp 1677677812
transform 1 0 1900 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2804
timestamp 1677677812
transform 1 0 1900 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2788
timestamp 1677677812
transform 1 0 1916 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3132
timestamp 1677677812
transform 1 0 1924 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2789
timestamp 1677677812
transform 1 0 1932 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3133
timestamp 1677677812
transform 1 0 1940 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3230
timestamp 1677677812
transform 1 0 1932 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2805
timestamp 1677677812
transform 1 0 1940 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2853
timestamp 1677677812
transform 1 0 1916 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2854
timestamp 1677677812
transform 1 0 1932 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3134
timestamp 1677677812
transform 1 0 1980 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2806
timestamp 1677677812
transform 1 0 1980 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3231
timestamp 1677677812
transform 1 0 2012 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2855
timestamp 1677677812
transform 1 0 2012 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3135
timestamp 1677677812
transform 1 0 2044 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3136
timestamp 1677677812
transform 1 0 2060 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3232
timestamp 1677677812
transform 1 0 2060 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3137
timestamp 1677677812
transform 1 0 2100 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2790
timestamp 1677677812
transform 1 0 2108 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3138
timestamp 1677677812
transform 1 0 2116 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2807
timestamp 1677677812
transform 1 0 2092 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3233
timestamp 1677677812
transform 1 0 2108 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2856
timestamp 1677677812
transform 1 0 2108 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2791
timestamp 1677677812
transform 1 0 2140 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2710
timestamp 1677677812
transform 1 0 2180 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3234
timestamp 1677677812
transform 1 0 2180 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3235
timestamp 1677677812
transform 1 0 2196 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3139
timestamp 1677677812
transform 1 0 2220 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2692
timestamp 1677677812
transform 1 0 2276 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2725
timestamp 1677677812
transform 1 0 2268 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2792
timestamp 1677677812
transform 1 0 2260 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3140
timestamp 1677677812
transform 1 0 2268 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3141
timestamp 1677677812
transform 1 0 2284 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3236
timestamp 1677677812
transform 1 0 2252 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3237
timestamp 1677677812
transform 1 0 2276 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3238
timestamp 1677677812
transform 1 0 2308 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2758
timestamp 1677677812
transform 1 0 2340 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3239
timestamp 1677677812
transform 1 0 2340 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3142
timestamp 1677677812
transform 1 0 2356 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3143
timestamp 1677677812
transform 1 0 2364 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2711
timestamp 1677677812
transform 1 0 2396 0 1 3255
box -3 -3 3 3
use M3_M2  M3_M2_2759
timestamp 1677677812
transform 1 0 2396 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2760
timestamp 1677677812
transform 1 0 2412 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2793
timestamp 1677677812
transform 1 0 2388 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3144
timestamp 1677677812
transform 1 0 2396 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3240
timestamp 1677677812
transform 1 0 2388 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3241
timestamp 1677677812
transform 1 0 2404 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2823
timestamp 1677677812
transform 1 0 2380 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2794
timestamp 1677677812
transform 1 0 2420 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3079
timestamp 1677677812
transform 1 0 2436 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3145
timestamp 1677677812
transform 1 0 2428 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3242
timestamp 1677677812
transform 1 0 2420 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2824
timestamp 1677677812
transform 1 0 2436 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2726
timestamp 1677677812
transform 1 0 2476 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2761
timestamp 1677677812
transform 1 0 2484 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3146
timestamp 1677677812
transform 1 0 2476 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2795
timestamp 1677677812
transform 1 0 2484 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3147
timestamp 1677677812
transform 1 0 2492 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3243
timestamp 1677677812
transform 1 0 2468 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2808
timestamp 1677677812
transform 1 0 2476 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3244
timestamp 1677677812
transform 1 0 2484 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2825
timestamp 1677677812
transform 1 0 2500 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2727
timestamp 1677677812
transform 1 0 2532 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3245
timestamp 1677677812
transform 1 0 2532 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2728
timestamp 1677677812
transform 1 0 2556 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2826
timestamp 1677677812
transform 1 0 2556 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3295
timestamp 1677677812
transform 1 0 2564 0 1 3195
box -2 -2 2 2
use M2_M1  M2_M1_3080
timestamp 1677677812
transform 1 0 2580 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2827
timestamp 1677677812
transform 1 0 2580 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3246
timestamp 1677677812
transform 1 0 2596 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3148
timestamp 1677677812
transform 1 0 2612 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2796
timestamp 1677677812
transform 1 0 2644 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2762
timestamp 1677677812
transform 1 0 2676 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3149
timestamp 1677677812
transform 1 0 2652 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3150
timestamp 1677677812
transform 1 0 2668 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3247
timestamp 1677677812
transform 1 0 2644 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3151
timestamp 1677677812
transform 1 0 2692 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3248
timestamp 1677677812
transform 1 0 2660 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3249
timestamp 1677677812
transform 1 0 2676 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3250
timestamp 1677677812
transform 1 0 2684 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2763
timestamp 1677677812
transform 1 0 2812 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2764
timestamp 1677677812
transform 1 0 2828 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3152
timestamp 1677677812
transform 1 0 2732 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3153
timestamp 1677677812
transform 1 0 2772 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3154
timestamp 1677677812
transform 1 0 2828 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3251
timestamp 1677677812
transform 1 0 2748 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2857
timestamp 1677677812
transform 1 0 2812 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2809
timestamp 1677677812
transform 1 0 2836 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3296
timestamp 1677677812
transform 1 0 2836 0 1 3195
box -2 -2 2 2
use M3_M2  M3_M2_2693
timestamp 1677677812
transform 1 0 2868 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2858
timestamp 1677677812
transform 1 0 2860 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2712
timestamp 1677677812
transform 1 0 2916 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3155
timestamp 1677677812
transform 1 0 2932 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3252
timestamp 1677677812
transform 1 0 2916 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3253
timestamp 1677677812
transform 1 0 2924 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2828
timestamp 1677677812
transform 1 0 2924 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3081
timestamp 1677677812
transform 1 0 2972 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3156
timestamp 1677677812
transform 1 0 2996 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3157
timestamp 1677677812
transform 1 0 3036 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2694
timestamp 1677677812
transform 1 0 3060 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3254
timestamp 1677677812
transform 1 0 3044 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2810
timestamp 1677677812
transform 1 0 3052 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2859
timestamp 1677677812
transform 1 0 3076 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2729
timestamp 1677677812
transform 1 0 3092 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2765
timestamp 1677677812
transform 1 0 3100 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3158
timestamp 1677677812
transform 1 0 3092 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2695
timestamp 1677677812
transform 1 0 3116 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2766
timestamp 1677677812
transform 1 0 3140 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3159
timestamp 1677677812
transform 1 0 3116 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3160
timestamp 1677677812
transform 1 0 3132 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3161
timestamp 1677677812
transform 1 0 3140 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3162
timestamp 1677677812
transform 1 0 3204 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3255
timestamp 1677677812
transform 1 0 3100 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3256
timestamp 1677677812
transform 1 0 3108 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3257
timestamp 1677677812
transform 1 0 3124 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3258
timestamp 1677677812
transform 1 0 3140 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3259
timestamp 1677677812
transform 1 0 3228 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2829
timestamp 1677677812
transform 1 0 3124 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2860
timestamp 1677677812
transform 1 0 3132 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2830
timestamp 1677677812
transform 1 0 3204 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2696
timestamp 1677677812
transform 1 0 3268 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2730
timestamp 1677677812
transform 1 0 3268 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3260
timestamp 1677677812
transform 1 0 3260 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2831
timestamp 1677677812
transform 1 0 3260 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3163
timestamp 1677677812
transform 1 0 3276 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3164
timestamp 1677677812
transform 1 0 3292 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3261
timestamp 1677677812
transform 1 0 3284 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2811
timestamp 1677677812
transform 1 0 3292 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3165
timestamp 1677677812
transform 1 0 3308 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3262
timestamp 1677677812
transform 1 0 3300 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2861
timestamp 1677677812
transform 1 0 3276 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2697
timestamp 1677677812
transform 1 0 3324 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2812
timestamp 1677677812
transform 1 0 3324 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2698
timestamp 1677677812
transform 1 0 3356 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3082
timestamp 1677677812
transform 1 0 3356 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3263
timestamp 1677677812
transform 1 0 3364 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2731
timestamp 1677677812
transform 1 0 3404 0 1 3245
box -3 -3 3 3
use M3_M2  M3_M2_2741
timestamp 1677677812
transform 1 0 3388 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3072
timestamp 1677677812
transform 1 0 3396 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_3083
timestamp 1677677812
transform 1 0 3412 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3166
timestamp 1677677812
transform 1 0 3404 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2699
timestamp 1677677812
transform 1 0 3484 0 1 3265
box -3 -3 3 3
use M2_M1  M2_M1_3073
timestamp 1677677812
transform 1 0 3468 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_3084
timestamp 1677677812
transform 1 0 3460 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2767
timestamp 1677677812
transform 1 0 3468 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3085
timestamp 1677677812
transform 1 0 3484 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2768
timestamp 1677677812
transform 1 0 3508 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3074
timestamp 1677677812
transform 1 0 3540 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_3086
timestamp 1677677812
transform 1 0 3548 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2797
timestamp 1677677812
transform 1 0 3540 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3167
timestamp 1677677812
transform 1 0 3548 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2732
timestamp 1677677812
transform 1 0 3564 0 1 3245
box -3 -3 3 3
use M2_M1  M2_M1_3087
timestamp 1677677812
transform 1 0 3564 0 1 3225
box -2 -2 2 2
use M3_M2  M3_M2_2832
timestamp 1677677812
transform 1 0 3572 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2713
timestamp 1677677812
transform 1 0 3604 0 1 3255
box -3 -3 3 3
use M2_M1  M2_M1_3075
timestamp 1677677812
transform 1 0 3604 0 1 3235
box -2 -2 2 2
use M2_M1  M2_M1_3264
timestamp 1677677812
transform 1 0 3612 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2813
timestamp 1677677812
transform 1 0 3620 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2742
timestamp 1677677812
transform 1 0 3708 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3088
timestamp 1677677812
transform 1 0 3708 0 1 3225
box -2 -2 2 2
use M2_M1  M2_M1_3265
timestamp 1677677812
transform 1 0 3716 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2798
timestamp 1677677812
transform 1 0 3780 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3266
timestamp 1677677812
transform 1 0 3780 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3168
timestamp 1677677812
transform 1 0 3788 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2769
timestamp 1677677812
transform 1 0 3820 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3169
timestamp 1677677812
transform 1 0 3804 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3170
timestamp 1677677812
transform 1 0 3820 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3171
timestamp 1677677812
transform 1 0 3836 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3267
timestamp 1677677812
transform 1 0 3812 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3268
timestamp 1677677812
transform 1 0 3828 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2833
timestamp 1677677812
transform 1 0 3828 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2743
timestamp 1677677812
transform 1 0 3900 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3172
timestamp 1677677812
transform 1 0 3900 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3173
timestamp 1677677812
transform 1 0 3916 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3269
timestamp 1677677812
transform 1 0 3892 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2834
timestamp 1677677812
transform 1 0 3892 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3174
timestamp 1677677812
transform 1 0 3932 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2770
timestamp 1677677812
transform 1 0 3940 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3270
timestamp 1677677812
transform 1 0 3940 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2835
timestamp 1677677812
transform 1 0 3932 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3271
timestamp 1677677812
transform 1 0 3956 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2862
timestamp 1677677812
transform 1 0 3948 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2799
timestamp 1677677812
transform 1 0 3988 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3272
timestamp 1677677812
transform 1 0 3988 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2863
timestamp 1677677812
transform 1 0 3988 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2744
timestamp 1677677812
transform 1 0 4028 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3175
timestamp 1677677812
transform 1 0 4012 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3176
timestamp 1677677812
transform 1 0 4028 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3273
timestamp 1677677812
transform 1 0 4020 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3274
timestamp 1677677812
transform 1 0 4036 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3275
timestamp 1677677812
transform 1 0 4044 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3276
timestamp 1677677812
transform 1 0 4052 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2836
timestamp 1677677812
transform 1 0 4012 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2837
timestamp 1677677812
transform 1 0 4044 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2864
timestamp 1677677812
transform 1 0 4044 0 1 3185
box -3 -3 3 3
use M3_M2  M3_M2_2745
timestamp 1677677812
transform 1 0 4108 0 1 3235
box -3 -3 3 3
use M3_M2  M3_M2_2771
timestamp 1677677812
transform 1 0 4092 0 1 3225
box -3 -3 3 3
use M3_M2  M3_M2_2772
timestamp 1677677812
transform 1 0 4116 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3177
timestamp 1677677812
transform 1 0 4092 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3178
timestamp 1677677812
transform 1 0 4108 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3179
timestamp 1677677812
transform 1 0 4116 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2814
timestamp 1677677812
transform 1 0 4092 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3277
timestamp 1677677812
transform 1 0 4100 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3278
timestamp 1677677812
transform 1 0 4116 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2838
timestamp 1677677812
transform 1 0 4116 0 1 3195
box -3 -3 3 3
use M2_M1  M2_M1_3279
timestamp 1677677812
transform 1 0 4172 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3280
timestamp 1677677812
transform 1 0 4196 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3180
timestamp 1677677812
transform 1 0 4228 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2815
timestamp 1677677812
transform 1 0 4220 0 1 3205
box -3 -3 3 3
use M3_M2  M3_M2_2800
timestamp 1677677812
transform 1 0 4236 0 1 3215
box -3 -3 3 3
use M2_M1  M2_M1_3181
timestamp 1677677812
transform 1 0 4244 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3182
timestamp 1677677812
transform 1 0 4260 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2839
timestamp 1677677812
transform 1 0 4228 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2865
timestamp 1677677812
transform 1 0 4228 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3281
timestamp 1677677812
transform 1 0 4244 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2816
timestamp 1677677812
transform 1 0 4268 0 1 3205
box -3 -3 3 3
use M2_M1  M2_M1_3282
timestamp 1677677812
transform 1 0 4276 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2840
timestamp 1677677812
transform 1 0 4252 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2841
timestamp 1677677812
transform 1 0 4276 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2866
timestamp 1677677812
transform 1 0 4276 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3183
timestamp 1677677812
transform 1 0 4308 0 1 3215
box -2 -2 2 2
use M3_M2  M3_M2_2700
timestamp 1677677812
transform 1 0 4324 0 1 3265
box -3 -3 3 3
use M3_M2  M3_M2_2801
timestamp 1677677812
transform 1 0 4420 0 1 3215
box -3 -3 3 3
use M3_M2  M3_M2_2746
timestamp 1677677812
transform 1 0 4580 0 1 3235
box -3 -3 3 3
use M2_M1  M2_M1_3184
timestamp 1677677812
transform 1 0 4516 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3185
timestamp 1677677812
transform 1 0 4572 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3186
timestamp 1677677812
transform 1 0 4580 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3283
timestamp 1677677812
transform 1 0 4492 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3284
timestamp 1677677812
transform 1 0 4596 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2867
timestamp 1677677812
transform 1 0 4596 0 1 3185
box -3 -3 3 3
use M2_M1  M2_M1_3285
timestamp 1677677812
transform 1 0 4628 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3286
timestamp 1677677812
transform 1 0 4644 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2842
timestamp 1677677812
transform 1 0 4636 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2773
timestamp 1677677812
transform 1 0 4684 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3187
timestamp 1677677812
transform 1 0 4692 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3188
timestamp 1677677812
transform 1 0 4708 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3287
timestamp 1677677812
transform 1 0 4684 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3288
timestamp 1677677812
transform 1 0 4700 0 1 3205
box -2 -2 2 2
use M3_M2  M3_M2_2843
timestamp 1677677812
transform 1 0 4700 0 1 3195
box -3 -3 3 3
use M3_M2  M3_M2_2774
timestamp 1677677812
transform 1 0 4740 0 1 3225
box -3 -3 3 3
use M2_M1  M2_M1_3189
timestamp 1677677812
transform 1 0 4756 0 1 3215
box -2 -2 2 2
use M2_M1  M2_M1_3289
timestamp 1677677812
transform 1 0 4748 0 1 3205
box -2 -2 2 2
use M2_M1  M2_M1_3290
timestamp 1677677812
transform 1 0 4764 0 1 3205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_30
timestamp 1677677812
transform 1 0 48 0 1 3170
box -10 -3 10 3
use M3_M2  M3_M2_2868
timestamp 1677677812
transform 1 0 116 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2869
timestamp 1677677812
transform 1 0 148 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_217
timestamp 1677677812
transform 1 0 72 0 1 3170
box -8 -3 104 105
use INVX2  INVX2_244
timestamp 1677677812
transform -1 0 184 0 1 3170
box -9 -3 26 105
use AOI22X1  AOI22X1_138
timestamp 1677677812
transform -1 0 224 0 1 3170
box -8 -3 46 105
use M3_M2  M3_M2_2870
timestamp 1677677812
transform 1 0 236 0 1 3175
box -3 -3 3 3
use FILL  FILL_3230
timestamp 1677677812
transform 1 0 224 0 1 3170
box -8 -3 16 105
use FILL  FILL_3231
timestamp 1677677812
transform 1 0 232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3234
timestamp 1677677812
transform 1 0 240 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_246
timestamp 1677677812
transform 1 0 248 0 1 3170
box -9 -3 26 105
use FILL  FILL_3236
timestamp 1677677812
transform 1 0 264 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2871
timestamp 1677677812
transform 1 0 300 0 1 3175
box -3 -3 3 3
use M3_M2  M3_M2_2872
timestamp 1677677812
transform 1 0 372 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_219
timestamp 1677677812
transform -1 0 368 0 1 3170
box -8 -3 104 105
use FILL  FILL_3237
timestamp 1677677812
transform 1 0 368 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2873
timestamp 1677677812
transform 1 0 404 0 1 3175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_220
timestamp 1677677812
transform 1 0 376 0 1 3170
box -8 -3 104 105
use FILL  FILL_3238
timestamp 1677677812
transform 1 0 472 0 1 3170
box -8 -3 16 105
use FILL  FILL_3239
timestamp 1677677812
transform 1 0 480 0 1 3170
box -8 -3 16 105
use FILL  FILL_3240
timestamp 1677677812
transform 1 0 488 0 1 3170
box -8 -3 16 105
use FILL  FILL_3241
timestamp 1677677812
transform 1 0 496 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_248
timestamp 1677677812
transform 1 0 504 0 1 3170
box -9 -3 26 105
use FILL  FILL_3257
timestamp 1677677812
transform 1 0 520 0 1 3170
box -8 -3 16 105
use FILL  FILL_3261
timestamp 1677677812
transform 1 0 528 0 1 3170
box -8 -3 16 105
use FILL  FILL_3262
timestamp 1677677812
transform 1 0 536 0 1 3170
box -8 -3 16 105
use FILL  FILL_3263
timestamp 1677677812
transform 1 0 544 0 1 3170
box -8 -3 16 105
use FILL  FILL_3264
timestamp 1677677812
transform 1 0 552 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_143
timestamp 1677677812
transform -1 0 600 0 1 3170
box -8 -3 46 105
use FILL  FILL_3265
timestamp 1677677812
transform 1 0 600 0 1 3170
box -8 -3 16 105
use FILL  FILL_3266
timestamp 1677677812
transform 1 0 608 0 1 3170
box -8 -3 16 105
use FILL  FILL_3267
timestamp 1677677812
transform 1 0 616 0 1 3170
box -8 -3 16 105
use FILL  FILL_3273
timestamp 1677677812
transform 1 0 624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3275
timestamp 1677677812
transform 1 0 632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3277
timestamp 1677677812
transform 1 0 640 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2874
timestamp 1677677812
transform 1 0 668 0 1 3175
box -3 -3 3 3
use OAI22X1  OAI22X1_137
timestamp 1677677812
transform 1 0 648 0 1 3170
box -8 -3 46 105
use FILL  FILL_3279
timestamp 1677677812
transform 1 0 688 0 1 3170
box -8 -3 16 105
use FILL  FILL_3280
timestamp 1677677812
transform 1 0 696 0 1 3170
box -8 -3 16 105
use FILL  FILL_3281
timestamp 1677677812
transform 1 0 704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3282
timestamp 1677677812
transform 1 0 712 0 1 3170
box -8 -3 16 105
use FILL  FILL_3283
timestamp 1677677812
transform 1 0 720 0 1 3170
box -8 -3 16 105
use FILL  FILL_3284
timestamp 1677677812
transform 1 0 728 0 1 3170
box -8 -3 16 105
use FILL  FILL_3285
timestamp 1677677812
transform 1 0 736 0 1 3170
box -8 -3 16 105
use FILL  FILL_3286
timestamp 1677677812
transform 1 0 744 0 1 3170
box -8 -3 16 105
use FILL  FILL_3288
timestamp 1677677812
transform 1 0 752 0 1 3170
box -8 -3 16 105
use FILL  FILL_3290
timestamp 1677677812
transform 1 0 760 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_145
timestamp 1677677812
transform 1 0 768 0 1 3170
box -8 -3 46 105
use FILL  FILL_3292
timestamp 1677677812
transform 1 0 808 0 1 3170
box -8 -3 16 105
use FILL  FILL_3293
timestamp 1677677812
transform 1 0 816 0 1 3170
box -8 -3 16 105
use FILL  FILL_3294
timestamp 1677677812
transform 1 0 824 0 1 3170
box -8 -3 16 105
use FILL  FILL_3298
timestamp 1677677812
transform 1 0 832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3300
timestamp 1677677812
transform 1 0 840 0 1 3170
box -8 -3 16 105
use FILL  FILL_3302
timestamp 1677677812
transform 1 0 848 0 1 3170
box -8 -3 16 105
use FILL  FILL_3304
timestamp 1677677812
transform 1 0 856 0 1 3170
box -8 -3 16 105
use FILL  FILL_3306
timestamp 1677677812
transform 1 0 864 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_33
timestamp 1677677812
transform 1 0 872 0 1 3170
box -8 -3 32 105
use FILL  FILL_3308
timestamp 1677677812
transform 1 0 896 0 1 3170
box -8 -3 16 105
use FILL  FILL_3309
timestamp 1677677812
transform 1 0 904 0 1 3170
box -8 -3 16 105
use FILL  FILL_3310
timestamp 1677677812
transform 1 0 912 0 1 3170
box -8 -3 16 105
use FILL  FILL_3311
timestamp 1677677812
transform 1 0 920 0 1 3170
box -8 -3 16 105
use FILL  FILL_3315
timestamp 1677677812
transform 1 0 928 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_72
timestamp 1677677812
transform 1 0 936 0 1 3170
box -8 -3 34 105
use FILL  FILL_3317
timestamp 1677677812
transform 1 0 968 0 1 3170
box -8 -3 16 105
use FILL  FILL_3323
timestamp 1677677812
transform 1 0 976 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2875
timestamp 1677677812
transform 1 0 996 0 1 3175
box -3 -3 3 3
use FILL  FILL_3325
timestamp 1677677812
transform 1 0 984 0 1 3170
box -8 -3 16 105
use FILL  FILL_3326
timestamp 1677677812
transform 1 0 992 0 1 3170
box -8 -3 16 105
use FILL  FILL_3327
timestamp 1677677812
transform 1 0 1000 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_34
timestamp 1677677812
transform 1 0 1008 0 1 3170
box -8 -3 32 105
use FILL  FILL_3328
timestamp 1677677812
transform 1 0 1032 0 1 3170
box -8 -3 16 105
use FILL  FILL_3331
timestamp 1677677812
transform 1 0 1040 0 1 3170
box -8 -3 16 105
use FILL  FILL_3333
timestamp 1677677812
transform 1 0 1048 0 1 3170
box -8 -3 16 105
use FILL  FILL_3335
timestamp 1677677812
transform 1 0 1056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3337
timestamp 1677677812
transform 1 0 1064 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_148
timestamp 1677677812
transform 1 0 1072 0 1 3170
box -8 -3 46 105
use FILL  FILL_3339
timestamp 1677677812
transform 1 0 1112 0 1 3170
box -8 -3 16 105
use FILL  FILL_3340
timestamp 1677677812
transform 1 0 1120 0 1 3170
box -8 -3 16 105
use FILL  FILL_3341
timestamp 1677677812
transform 1 0 1128 0 1 3170
box -8 -3 16 105
use FILL  FILL_3346
timestamp 1677677812
transform 1 0 1136 0 1 3170
box -8 -3 16 105
use FILL  FILL_3348
timestamp 1677677812
transform 1 0 1144 0 1 3170
box -8 -3 16 105
use FILL  FILL_3350
timestamp 1677677812
transform 1 0 1152 0 1 3170
box -8 -3 16 105
use FILL  FILL_3352
timestamp 1677677812
transform 1 0 1160 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_149
timestamp 1677677812
transform -1 0 1208 0 1 3170
box -8 -3 46 105
use FILL  FILL_3353
timestamp 1677677812
transform 1 0 1208 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2876
timestamp 1677677812
transform 1 0 1228 0 1 3175
box -3 -3 3 3
use FILL  FILL_3361
timestamp 1677677812
transform 1 0 1216 0 1 3170
box -8 -3 16 105
use FILL  FILL_3363
timestamp 1677677812
transform 1 0 1224 0 1 3170
box -8 -3 16 105
use FILL  FILL_3365
timestamp 1677677812
transform 1 0 1232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3367
timestamp 1677677812
transform 1 0 1240 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_74
timestamp 1677677812
transform -1 0 1280 0 1 3170
box -8 -3 34 105
use FILL  FILL_3368
timestamp 1677677812
transform 1 0 1280 0 1 3170
box -8 -3 16 105
use FILL  FILL_3369
timestamp 1677677812
transform 1 0 1288 0 1 3170
box -8 -3 16 105
use FILL  FILL_3370
timestamp 1677677812
transform 1 0 1296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3375
timestamp 1677677812
transform 1 0 1304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3377
timestamp 1677677812
transform 1 0 1312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3379
timestamp 1677677812
transform 1 0 1320 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_76
timestamp 1677677812
transform -1 0 1360 0 1 3170
box -8 -3 34 105
use FILL  FILL_3380
timestamp 1677677812
transform 1 0 1360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3381
timestamp 1677677812
transform 1 0 1368 0 1 3170
box -8 -3 16 105
use FILL  FILL_3382
timestamp 1677677812
transform 1 0 1376 0 1 3170
box -8 -3 16 105
use FILL  FILL_3387
timestamp 1677677812
transform 1 0 1384 0 1 3170
box -8 -3 16 105
use FILL  FILL_3389
timestamp 1677677812
transform 1 0 1392 0 1 3170
box -8 -3 16 105
use FILL  FILL_3391
timestamp 1677677812
transform 1 0 1400 0 1 3170
box -8 -3 16 105
use FILL  FILL_3393
timestamp 1677677812
transform 1 0 1408 0 1 3170
box -8 -3 16 105
use FILL  FILL_3395
timestamp 1677677812
transform 1 0 1416 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_138
timestamp 1677677812
transform -1 0 1464 0 1 3170
box -8 -3 46 105
use FILL  FILL_3396
timestamp 1677677812
transform 1 0 1464 0 1 3170
box -8 -3 16 105
use FILL  FILL_3402
timestamp 1677677812
transform 1 0 1472 0 1 3170
box -8 -3 16 105
use FILL  FILL_3404
timestamp 1677677812
transform 1 0 1480 0 1 3170
box -8 -3 16 105
use FILL  FILL_3406
timestamp 1677677812
transform 1 0 1488 0 1 3170
box -8 -3 16 105
use FILL  FILL_3407
timestamp 1677677812
transform 1 0 1496 0 1 3170
box -8 -3 16 105
use FILL  FILL_3408
timestamp 1677677812
transform 1 0 1504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3409
timestamp 1677677812
transform 1 0 1512 0 1 3170
box -8 -3 16 105
use FILL  FILL_3412
timestamp 1677677812
transform 1 0 1520 0 1 3170
box -8 -3 16 105
use FILL  FILL_3414
timestamp 1677677812
transform 1 0 1528 0 1 3170
box -8 -3 16 105
use FILL  FILL_3416
timestamp 1677677812
transform 1 0 1536 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_139
timestamp 1677677812
transform -1 0 1584 0 1 3170
box -8 -3 46 105
use FILL  FILL_3417
timestamp 1677677812
transform 1 0 1584 0 1 3170
box -8 -3 16 105
use FILL  FILL_3418
timestamp 1677677812
transform 1 0 1592 0 1 3170
box -8 -3 16 105
use FILL  FILL_3422
timestamp 1677677812
transform 1 0 1600 0 1 3170
box -8 -3 16 105
use FILL  FILL_3424
timestamp 1677677812
transform 1 0 1608 0 1 3170
box -8 -3 16 105
use FILL  FILL_3426
timestamp 1677677812
transform 1 0 1616 0 1 3170
box -8 -3 16 105
use FILL  FILL_3427
timestamp 1677677812
transform 1 0 1624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3428
timestamp 1677677812
transform 1 0 1632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3429
timestamp 1677677812
transform 1 0 1640 0 1 3170
box -8 -3 16 105
use FILL  FILL_3430
timestamp 1677677812
transform 1 0 1648 0 1 3170
box -8 -3 16 105
use FILL  FILL_3431
timestamp 1677677812
transform 1 0 1656 0 1 3170
box -8 -3 16 105
use FILL  FILL_3432
timestamp 1677677812
transform 1 0 1664 0 1 3170
box -8 -3 16 105
use FILL  FILL_3433
timestamp 1677677812
transform 1 0 1672 0 1 3170
box -8 -3 16 105
use FILL  FILL_3434
timestamp 1677677812
transform 1 0 1680 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_22
timestamp 1677677812
transform -1 0 1712 0 1 3170
box -5 -3 28 105
use FILL  FILL_3435
timestamp 1677677812
transform 1 0 1712 0 1 3170
box -8 -3 16 105
use FILL  FILL_3437
timestamp 1677677812
transform 1 0 1720 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_23
timestamp 1677677812
transform 1 0 1728 0 1 3170
box -5 -3 28 105
use FILL  FILL_3439
timestamp 1677677812
transform 1 0 1752 0 1 3170
box -8 -3 16 105
use FILL  FILL_3444
timestamp 1677677812
transform 1 0 1760 0 1 3170
box -8 -3 16 105
use FILL  FILL_3446
timestamp 1677677812
transform 1 0 1768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3448
timestamp 1677677812
transform 1 0 1776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3449
timestamp 1677677812
transform 1 0 1784 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_24
timestamp 1677677812
transform 1 0 1792 0 1 3170
box -5 -3 28 105
use FILL  FILL_3450
timestamp 1677677812
transform 1 0 1816 0 1 3170
box -8 -3 16 105
use FILL  FILL_3451
timestamp 1677677812
transform 1 0 1824 0 1 3170
box -8 -3 16 105
use FILL  FILL_3452
timestamp 1677677812
transform 1 0 1832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3453
timestamp 1677677812
transform 1 0 1840 0 1 3170
box -8 -3 16 105
use FILL  FILL_3454
timestamp 1677677812
transform 1 0 1848 0 1 3170
box -8 -3 16 105
use FILL  FILL_3455
timestamp 1677677812
transform 1 0 1856 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_252
timestamp 1677677812
transform -1 0 1880 0 1 3170
box -9 -3 26 105
use FILL  FILL_3456
timestamp 1677677812
transform 1 0 1880 0 1 3170
box -8 -3 16 105
use FILL  FILL_3459
timestamp 1677677812
transform 1 0 1888 0 1 3170
box -8 -3 16 105
use FILL  FILL_3461
timestamp 1677677812
transform 1 0 1896 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_150
timestamp 1677677812
transform -1 0 1944 0 1 3170
box -8 -3 46 105
use FILL  FILL_3462
timestamp 1677677812
transform 1 0 1944 0 1 3170
box -8 -3 16 105
use FILL  FILL_3465
timestamp 1677677812
transform 1 0 1952 0 1 3170
box -8 -3 16 105
use FILL  FILL_3467
timestamp 1677677812
transform 1 0 1960 0 1 3170
box -8 -3 16 105
use FILL  FILL_3469
timestamp 1677677812
transform 1 0 1968 0 1 3170
box -8 -3 16 105
use FILL  FILL_3471
timestamp 1677677812
transform 1 0 1976 0 1 3170
box -8 -3 16 105
use FILL  FILL_3472
timestamp 1677677812
transform 1 0 1984 0 1 3170
box -8 -3 16 105
use FILL  FILL_3473
timestamp 1677677812
transform 1 0 1992 0 1 3170
box -8 -3 16 105
use FILL  FILL_3475
timestamp 1677677812
transform 1 0 2000 0 1 3170
box -8 -3 16 105
use FILL  FILL_3477
timestamp 1677677812
transform 1 0 2008 0 1 3170
box -8 -3 16 105
use FILL  FILL_3478
timestamp 1677677812
transform 1 0 2016 0 1 3170
box -8 -3 16 105
use FILL  FILL_3479
timestamp 1677677812
transform 1 0 2024 0 1 3170
box -8 -3 16 105
use FILL  FILL_3480
timestamp 1677677812
transform 1 0 2032 0 1 3170
box -8 -3 16 105
use FILL  FILL_3481
timestamp 1677677812
transform 1 0 2040 0 1 3170
box -8 -3 16 105
use FILL  FILL_3482
timestamp 1677677812
transform 1 0 2048 0 1 3170
box -8 -3 16 105
use FILL  FILL_3484
timestamp 1677677812
transform 1 0 2056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3486
timestamp 1677677812
transform 1 0 2064 0 1 3170
box -8 -3 16 105
use FILL  FILL_3488
timestamp 1677677812
transform 1 0 2072 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_153
timestamp 1677677812
transform -1 0 2120 0 1 3170
box -8 -3 46 105
use FILL  FILL_3489
timestamp 1677677812
transform 1 0 2120 0 1 3170
box -8 -3 16 105
use FILL  FILL_3490
timestamp 1677677812
transform 1 0 2128 0 1 3170
box -8 -3 16 105
use FILL  FILL_3491
timestamp 1677677812
transform 1 0 2136 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2877
timestamp 1677677812
transform 1 0 2156 0 1 3175
box -3 -3 3 3
use FILL  FILL_3492
timestamp 1677677812
transform 1 0 2144 0 1 3170
box -8 -3 16 105
use FILL  FILL_3493
timestamp 1677677812
transform 1 0 2152 0 1 3170
box -8 -3 16 105
use FILL  FILL_3500
timestamp 1677677812
transform 1 0 2160 0 1 3170
box -8 -3 16 105
use FILL  FILL_3502
timestamp 1677677812
transform 1 0 2168 0 1 3170
box -8 -3 16 105
use FILL  FILL_3504
timestamp 1677677812
transform 1 0 2176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3506
timestamp 1677677812
transform 1 0 2184 0 1 3170
box -8 -3 16 105
use FILL  FILL_3507
timestamp 1677677812
transform 1 0 2192 0 1 3170
box -8 -3 16 105
use BUFX2  BUFX2_25
timestamp 1677677812
transform -1 0 2224 0 1 3170
box -5 -3 28 105
use FILL  FILL_3508
timestamp 1677677812
transform 1 0 2224 0 1 3170
box -8 -3 16 105
use FILL  FILL_3509
timestamp 1677677812
transform 1 0 2232 0 1 3170
box -8 -3 16 105
use FILL  FILL_3510
timestamp 1677677812
transform 1 0 2240 0 1 3170
box -8 -3 16 105
use FILL  FILL_3511
timestamp 1677677812
transform 1 0 2248 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_142
timestamp 1677677812
transform -1 0 2296 0 1 3170
box -8 -3 46 105
use FILL  FILL_3512
timestamp 1677677812
transform 1 0 2296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3513
timestamp 1677677812
transform 1 0 2304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3514
timestamp 1677677812
transform 1 0 2312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3515
timestamp 1677677812
transform 1 0 2320 0 1 3170
box -8 -3 16 105
use FILL  FILL_3519
timestamp 1677677812
transform 1 0 2328 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_254
timestamp 1677677812
transform 1 0 2336 0 1 3170
box -9 -3 26 105
use FILL  FILL_3520
timestamp 1677677812
transform 1 0 2352 0 1 3170
box -8 -3 16 105
use FILL  FILL_3521
timestamp 1677677812
transform 1 0 2360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3522
timestamp 1677677812
transform 1 0 2368 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_154
timestamp 1677677812
transform -1 0 2416 0 1 3170
box -8 -3 46 105
use FILL  FILL_3523
timestamp 1677677812
transform 1 0 2416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3524
timestamp 1677677812
transform 1 0 2424 0 1 3170
box -8 -3 16 105
use FILL  FILL_3526
timestamp 1677677812
transform 1 0 2432 0 1 3170
box -8 -3 16 105
use FILL  FILL_3528
timestamp 1677677812
transform 1 0 2440 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_143
timestamp 1677677812
transform 1 0 2448 0 1 3170
box -8 -3 46 105
use FILL  FILL_3530
timestamp 1677677812
transform 1 0 2488 0 1 3170
box -8 -3 16 105
use FILL  FILL_3535
timestamp 1677677812
transform 1 0 2496 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2878
timestamp 1677677812
transform 1 0 2516 0 1 3175
box -3 -3 3 3
use FILL  FILL_3537
timestamp 1677677812
transform 1 0 2504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3538
timestamp 1677677812
transform 1 0 2512 0 1 3170
box -8 -3 16 105
use FILL  FILL_3539
timestamp 1677677812
transform 1 0 2520 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_78
timestamp 1677677812
transform 1 0 2528 0 1 3170
box -8 -3 34 105
use FILL  FILL_3540
timestamp 1677677812
transform 1 0 2560 0 1 3170
box -8 -3 16 105
use FILL  FILL_3541
timestamp 1677677812
transform 1 0 2568 0 1 3170
box -8 -3 16 105
use FILL  FILL_3542
timestamp 1677677812
transform 1 0 2576 0 1 3170
box -8 -3 16 105
use FILL  FILL_3543
timestamp 1677677812
transform 1 0 2584 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_35
timestamp 1677677812
transform 1 0 2592 0 1 3170
box -8 -3 32 105
use FILL  FILL_3544
timestamp 1677677812
transform 1 0 2616 0 1 3170
box -8 -3 16 105
use FILL  FILL_3545
timestamp 1677677812
transform 1 0 2624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3546
timestamp 1677677812
transform 1 0 2632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3547
timestamp 1677677812
transform 1 0 2640 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2879
timestamp 1677677812
transform 1 0 2660 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_156
timestamp 1677677812
transform 1 0 2648 0 1 3170
box -8 -3 46 105
use FILL  FILL_3549
timestamp 1677677812
transform 1 0 2688 0 1 3170
box -8 -3 16 105
use FILL  FILL_3550
timestamp 1677677812
transform 1 0 2696 0 1 3170
box -8 -3 16 105
use FILL  FILL_3553
timestamp 1677677812
transform 1 0 2704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3554
timestamp 1677677812
transform 1 0 2712 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_256
timestamp 1677677812
transform 1 0 2720 0 1 3170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_227
timestamp 1677677812
transform 1 0 2736 0 1 3170
box -8 -3 104 105
use FILL  FILL_3555
timestamp 1677677812
transform 1 0 2832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3557
timestamp 1677677812
transform 1 0 2840 0 1 3170
box -8 -3 16 105
use FILL  FILL_3559
timestamp 1677677812
transform 1 0 2848 0 1 3170
box -8 -3 16 105
use FILL  FILL_3560
timestamp 1677677812
transform 1 0 2856 0 1 3170
box -8 -3 16 105
use FILL  FILL_3561
timestamp 1677677812
transform 1 0 2864 0 1 3170
box -8 -3 16 105
use FILL  FILL_3562
timestamp 1677677812
transform 1 0 2872 0 1 3170
box -8 -3 16 105
use FILL  FILL_3563
timestamp 1677677812
transform 1 0 2880 0 1 3170
box -8 -3 16 105
use FILL  FILL_3564
timestamp 1677677812
transform 1 0 2888 0 1 3170
box -8 -3 16 105
use FILL  FILL_3565
timestamp 1677677812
transform 1 0 2896 0 1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_38
timestamp 1677677812
transform 1 0 2904 0 1 3170
box -8 -3 32 105
use FILL  FILL_3567
timestamp 1677677812
transform 1 0 2928 0 1 3170
box -8 -3 16 105
use FILL  FILL_3568
timestamp 1677677812
transform 1 0 2936 0 1 3170
box -8 -3 16 105
use FILL  FILL_3569
timestamp 1677677812
transform 1 0 2944 0 1 3170
box -8 -3 16 105
use FILL  FILL_3570
timestamp 1677677812
transform 1 0 2952 0 1 3170
box -8 -3 16 105
use FILL  FILL_3571
timestamp 1677677812
transform 1 0 2960 0 1 3170
box -8 -3 16 105
use FILL  FILL_3576
timestamp 1677677812
transform 1 0 2968 0 1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_81
timestamp 1677677812
transform -1 0 3008 0 1 3170
box -8 -3 34 105
use FILL  FILL_3577
timestamp 1677677812
transform 1 0 3008 0 1 3170
box -8 -3 16 105
use FILL  FILL_3578
timestamp 1677677812
transform 1 0 3016 0 1 3170
box -8 -3 16 105
use FILL  FILL_3579
timestamp 1677677812
transform 1 0 3024 0 1 3170
box -8 -3 16 105
use FILL  FILL_3580
timestamp 1677677812
transform 1 0 3032 0 1 3170
box -8 -3 16 105
use FILL  FILL_3586
timestamp 1677677812
transform 1 0 3040 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_257
timestamp 1677677812
transform -1 0 3064 0 1 3170
box -9 -3 26 105
use FILL  FILL_3587
timestamp 1677677812
transform 1 0 3064 0 1 3170
box -8 -3 16 105
use FILL  FILL_3588
timestamp 1677677812
transform 1 0 3072 0 1 3170
box -8 -3 16 105
use FILL  FILL_3589
timestamp 1677677812
transform 1 0 3080 0 1 3170
box -8 -3 16 105
use FILL  FILL_3590
timestamp 1677677812
transform 1 0 3088 0 1 3170
box -8 -3 16 105
use FILL  FILL_3591
timestamp 1677677812
transform 1 0 3096 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_144
timestamp 1677677812
transform -1 0 3144 0 1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_229
timestamp 1677677812
transform -1 0 3240 0 1 3170
box -8 -3 104 105
use FILL  FILL_3592
timestamp 1677677812
transform 1 0 3240 0 1 3170
box -8 -3 16 105
use FILL  FILL_3602
timestamp 1677677812
transform 1 0 3248 0 1 3170
box -8 -3 16 105
use FILL  FILL_3603
timestamp 1677677812
transform 1 0 3256 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_146
timestamp 1677677812
transform 1 0 3264 0 1 3170
box -8 -3 46 105
use FILL  FILL_3604
timestamp 1677677812
transform 1 0 3304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3605
timestamp 1677677812
transform 1 0 3312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3606
timestamp 1677677812
transform 1 0 3320 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_258
timestamp 1677677812
transform -1 0 3344 0 1 3170
box -9 -3 26 105
use FILL  FILL_3607
timestamp 1677677812
transform 1 0 3344 0 1 3170
box -8 -3 16 105
use FILL  FILL_3608
timestamp 1677677812
transform 1 0 3352 0 1 3170
box -8 -3 16 105
use FILL  FILL_3609
timestamp 1677677812
transform 1 0 3360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3610
timestamp 1677677812
transform 1 0 3368 0 1 3170
box -8 -3 16 105
use FILL  FILL_3613
timestamp 1677677812
transform 1 0 3376 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_16
timestamp 1677677812
transform -1 0 3416 0 1 3170
box -8 -3 40 105
use FILL  FILL_3614
timestamp 1677677812
transform 1 0 3416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3615
timestamp 1677677812
transform 1 0 3424 0 1 3170
box -8 -3 16 105
use FILL  FILL_3619
timestamp 1677677812
transform 1 0 3432 0 1 3170
box -8 -3 16 105
use FILL  FILL_3621
timestamp 1677677812
transform 1 0 3440 0 1 3170
box -8 -3 16 105
use FILL  FILL_3623
timestamp 1677677812
transform 1 0 3448 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_18
timestamp 1677677812
transform -1 0 3488 0 1 3170
box -8 -3 40 105
use FILL  FILL_3624
timestamp 1677677812
transform 1 0 3488 0 1 3170
box -8 -3 16 105
use FILL  FILL_3631
timestamp 1677677812
transform 1 0 3496 0 1 3170
box -8 -3 16 105
use FILL  FILL_3632
timestamp 1677677812
transform 1 0 3504 0 1 3170
box -8 -3 16 105
use FILL  FILL_3633
timestamp 1677677812
transform 1 0 3512 0 1 3170
box -8 -3 16 105
use FILL  FILL_3634
timestamp 1677677812
transform 1 0 3520 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_19
timestamp 1677677812
transform -1 0 3560 0 1 3170
box -8 -3 40 105
use FILL  FILL_3635
timestamp 1677677812
transform 1 0 3560 0 1 3170
box -8 -3 16 105
use FILL  FILL_3640
timestamp 1677677812
transform 1 0 3568 0 1 3170
box -8 -3 16 105
use FILL  FILL_3642
timestamp 1677677812
transform 1 0 3576 0 1 3170
box -8 -3 16 105
use FILL  FILL_3644
timestamp 1677677812
transform 1 0 3584 0 1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_20
timestamp 1677677812
transform -1 0 3624 0 1 3170
box -8 -3 40 105
use FILL  FILL_3645
timestamp 1677677812
transform 1 0 3624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3646
timestamp 1677677812
transform 1 0 3632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3652
timestamp 1677677812
transform 1 0 3640 0 1 3170
box -8 -3 16 105
use FILL  FILL_3654
timestamp 1677677812
transform 1 0 3648 0 1 3170
box -8 -3 16 105
use FILL  FILL_3656
timestamp 1677677812
transform 1 0 3656 0 1 3170
box -8 -3 16 105
use FILL  FILL_3658
timestamp 1677677812
transform 1 0 3664 0 1 3170
box -8 -3 16 105
use FILL  FILL_3659
timestamp 1677677812
transform 1 0 3672 0 1 3170
box -8 -3 16 105
use FILL  FILL_3660
timestamp 1677677812
transform 1 0 3680 0 1 3170
box -8 -3 16 105
use FILL  FILL_3661
timestamp 1677677812
transform 1 0 3688 0 1 3170
box -8 -3 16 105
use FILL  FILL_3662
timestamp 1677677812
transform 1 0 3696 0 1 3170
box -8 -3 16 105
use FILL  FILL_3663
timestamp 1677677812
transform 1 0 3704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3666
timestamp 1677677812
transform 1 0 3712 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_261
timestamp 1677677812
transform 1 0 3720 0 1 3170
box -9 -3 26 105
use FILL  FILL_3668
timestamp 1677677812
transform 1 0 3736 0 1 3170
box -8 -3 16 105
use FILL  FILL_3672
timestamp 1677677812
transform 1 0 3744 0 1 3170
box -8 -3 16 105
use FILL  FILL_3674
timestamp 1677677812
transform 1 0 3752 0 1 3170
box -8 -3 16 105
use FILL  FILL_3676
timestamp 1677677812
transform 1 0 3760 0 1 3170
box -8 -3 16 105
use FILL  FILL_3678
timestamp 1677677812
transform 1 0 3768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3679
timestamp 1677677812
transform 1 0 3776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3680
timestamp 1677677812
transform 1 0 3784 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_147
timestamp 1677677812
transform -1 0 3832 0 1 3170
box -8 -3 46 105
use FILL  FILL_3681
timestamp 1677677812
transform 1 0 3832 0 1 3170
box -8 -3 16 105
use FILL  FILL_3682
timestamp 1677677812
transform 1 0 3840 0 1 3170
box -8 -3 16 105
use FILL  FILL_3683
timestamp 1677677812
transform 1 0 3848 0 1 3170
box -8 -3 16 105
use FILL  FILL_3684
timestamp 1677677812
transform 1 0 3856 0 1 3170
box -8 -3 16 105
use FILL  FILL_3685
timestamp 1677677812
transform 1 0 3864 0 1 3170
box -8 -3 16 105
use FILL  FILL_3686
timestamp 1677677812
transform 1 0 3872 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2880
timestamp 1677677812
transform 1 0 3924 0 1 3175
box -3 -3 3 3
use AOI22X1  AOI22X1_159
timestamp 1677677812
transform 1 0 3880 0 1 3170
box -8 -3 46 105
use FILL  FILL_3687
timestamp 1677677812
transform 1 0 3920 0 1 3170
box -8 -3 16 105
use FILL  FILL_3688
timestamp 1677677812
transform 1 0 3928 0 1 3170
box -8 -3 16 105
use FILL  FILL_3689
timestamp 1677677812
transform 1 0 3936 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_262
timestamp 1677677812
transform -1 0 3960 0 1 3170
box -9 -3 26 105
use FILL  FILL_3690
timestamp 1677677812
transform 1 0 3960 0 1 3170
box -8 -3 16 105
use FILL  FILL_3700
timestamp 1677677812
transform 1 0 3968 0 1 3170
box -8 -3 16 105
use FILL  FILL_3702
timestamp 1677677812
transform 1 0 3976 0 1 3170
box -8 -3 16 105
use FILL  FILL_3704
timestamp 1677677812
transform 1 0 3984 0 1 3170
box -8 -3 16 105
use FILL  FILL_3705
timestamp 1677677812
transform 1 0 3992 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_149
timestamp 1677677812
transform -1 0 4040 0 1 3170
box -8 -3 46 105
use M3_M2  M3_M2_2881
timestamp 1677677812
transform 1 0 4052 0 1 3175
box -3 -3 3 3
use FILL  FILL_3706
timestamp 1677677812
transform 1 0 4040 0 1 3170
box -8 -3 16 105
use FILL  FILL_3707
timestamp 1677677812
transform 1 0 4048 0 1 3170
box -8 -3 16 105
use FILL  FILL_3708
timestamp 1677677812
transform 1 0 4056 0 1 3170
box -8 -3 16 105
use FILL  FILL_3709
timestamp 1677677812
transform 1 0 4064 0 1 3170
box -8 -3 16 105
use FILL  FILL_3710
timestamp 1677677812
transform 1 0 4072 0 1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_150
timestamp 1677677812
transform -1 0 4120 0 1 3170
box -8 -3 46 105
use M3_M2  M3_M2_2882
timestamp 1677677812
transform 1 0 4132 0 1 3175
box -3 -3 3 3
use FILL  FILL_3711
timestamp 1677677812
transform 1 0 4120 0 1 3170
box -8 -3 16 105
use FILL  FILL_3712
timestamp 1677677812
transform 1 0 4128 0 1 3170
box -8 -3 16 105
use FILL  FILL_3713
timestamp 1677677812
transform 1 0 4136 0 1 3170
box -8 -3 16 105
use FILL  FILL_3714
timestamp 1677677812
transform 1 0 4144 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_264
timestamp 1677677812
transform -1 0 4168 0 1 3170
box -9 -3 26 105
use FILL  FILL_3715
timestamp 1677677812
transform 1 0 4168 0 1 3170
box -8 -3 16 105
use FILL  FILL_3716
timestamp 1677677812
transform 1 0 4176 0 1 3170
box -8 -3 16 105
use FILL  FILL_3717
timestamp 1677677812
transform 1 0 4184 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2883
timestamp 1677677812
transform 1 0 4204 0 1 3175
box -3 -3 3 3
use INVX2  INVX2_265
timestamp 1677677812
transform 1 0 4192 0 1 3170
box -9 -3 26 105
use FILL  FILL_3718
timestamp 1677677812
transform 1 0 4208 0 1 3170
box -8 -3 16 105
use FILL  FILL_3724
timestamp 1677677812
transform 1 0 4216 0 1 3170
box -8 -3 16 105
use FILL  FILL_3726
timestamp 1677677812
transform 1 0 4224 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2884
timestamp 1677677812
transform 1 0 4244 0 1 3175
box -3 -3 3 3
use FILL  FILL_3728
timestamp 1677677812
transform 1 0 4232 0 1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_161
timestamp 1677677812
transform -1 0 4280 0 1 3170
box -8 -3 46 105
use FILL  FILL_3730
timestamp 1677677812
transform 1 0 4280 0 1 3170
box -8 -3 16 105
use FILL  FILL_3732
timestamp 1677677812
transform 1 0 4288 0 1 3170
box -8 -3 16 105
use FILL  FILL_3734
timestamp 1677677812
transform 1 0 4296 0 1 3170
box -8 -3 16 105
use FILL  FILL_3736
timestamp 1677677812
transform 1 0 4304 0 1 3170
box -8 -3 16 105
use FILL  FILL_3738
timestamp 1677677812
transform 1 0 4312 0 1 3170
box -8 -3 16 105
use FILL  FILL_3739
timestamp 1677677812
transform 1 0 4320 0 1 3170
box -8 -3 16 105
use FILL  FILL_3740
timestamp 1677677812
transform 1 0 4328 0 1 3170
box -8 -3 16 105
use FILL  FILL_3741
timestamp 1677677812
transform 1 0 4336 0 1 3170
box -8 -3 16 105
use FILL  FILL_3742
timestamp 1677677812
transform 1 0 4344 0 1 3170
box -8 -3 16 105
use FILL  FILL_3743
timestamp 1677677812
transform 1 0 4352 0 1 3170
box -8 -3 16 105
use FILL  FILL_3745
timestamp 1677677812
transform 1 0 4360 0 1 3170
box -8 -3 16 105
use FILL  FILL_3747
timestamp 1677677812
transform 1 0 4368 0 1 3170
box -8 -3 16 105
use FILL  FILL_3749
timestamp 1677677812
transform 1 0 4376 0 1 3170
box -8 -3 16 105
use FILL  FILL_3751
timestamp 1677677812
transform 1 0 4384 0 1 3170
box -8 -3 16 105
use FILL  FILL_3752
timestamp 1677677812
transform 1 0 4392 0 1 3170
box -8 -3 16 105
use FILL  FILL_3753
timestamp 1677677812
transform 1 0 4400 0 1 3170
box -8 -3 16 105
use FILL  FILL_3754
timestamp 1677677812
transform 1 0 4408 0 1 3170
box -8 -3 16 105
use FILL  FILL_3755
timestamp 1677677812
transform 1 0 4416 0 1 3170
box -8 -3 16 105
use FILL  FILL_3756
timestamp 1677677812
transform 1 0 4424 0 1 3170
box -8 -3 16 105
use FILL  FILL_3758
timestamp 1677677812
transform 1 0 4432 0 1 3170
box -8 -3 16 105
use FILL  FILL_3760
timestamp 1677677812
transform 1 0 4440 0 1 3170
box -8 -3 16 105
use FILL  FILL_3762
timestamp 1677677812
transform 1 0 4448 0 1 3170
box -8 -3 16 105
use FILL  FILL_3764
timestamp 1677677812
transform 1 0 4456 0 1 3170
box -8 -3 16 105
use FILL  FILL_3765
timestamp 1677677812
transform 1 0 4464 0 1 3170
box -8 -3 16 105
use FILL  FILL_3766
timestamp 1677677812
transform 1 0 4472 0 1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_234
timestamp 1677677812
transform 1 0 4480 0 1 3170
box -8 -3 104 105
use FILL  FILL_3767
timestamp 1677677812
transform 1 0 4576 0 1 3170
box -8 -3 16 105
use FILL  FILL_3770
timestamp 1677677812
transform 1 0 4584 0 1 3170
box -8 -3 16 105
use FILL  FILL_3772
timestamp 1677677812
transform 1 0 4592 0 1 3170
box -8 -3 16 105
use FILL  FILL_3774
timestamp 1677677812
transform 1 0 4600 0 1 3170
box -8 -3 16 105
use FILL  FILL_3775
timestamp 1677677812
transform 1 0 4608 0 1 3170
box -8 -3 16 105
use FILL  FILL_3776
timestamp 1677677812
transform 1 0 4616 0 1 3170
box -8 -3 16 105
use FILL  FILL_3777
timestamp 1677677812
transform 1 0 4624 0 1 3170
box -8 -3 16 105
use FILL  FILL_3778
timestamp 1677677812
transform 1 0 4632 0 1 3170
box -8 -3 16 105
use FILL  FILL_3779
timestamp 1677677812
transform 1 0 4640 0 1 3170
box -8 -3 16 105
use FILL  FILL_3781
timestamp 1677677812
transform 1 0 4648 0 1 3170
box -8 -3 16 105
use FILL  FILL_3783
timestamp 1677677812
transform 1 0 4656 0 1 3170
box -8 -3 16 105
use M3_M2  M3_M2_2885
timestamp 1677677812
transform 1 0 4692 0 1 3175
box -3 -3 3 3
use OAI22X1  OAI22X1_154
timestamp 1677677812
transform 1 0 4664 0 1 3170
box -8 -3 46 105
use FILL  FILL_3785
timestamp 1677677812
transform 1 0 4704 0 1 3170
box -8 -3 16 105
use FILL  FILL_3786
timestamp 1677677812
transform 1 0 4712 0 1 3170
box -8 -3 16 105
use FILL  FILL_3787
timestamp 1677677812
transform 1 0 4720 0 1 3170
box -8 -3 16 105
use FILL  FILL_3788
timestamp 1677677812
transform 1 0 4728 0 1 3170
box -8 -3 16 105
use INVX2  INVX2_267
timestamp 1677677812
transform -1 0 4752 0 1 3170
box -9 -3 26 105
use INVX2  INVX2_268
timestamp 1677677812
transform -1 0 4768 0 1 3170
box -9 -3 26 105
use FILL  FILL_3789
timestamp 1677677812
transform 1 0 4768 0 1 3170
box -8 -3 16 105
use FILL  FILL_3792
timestamp 1677677812
transform 1 0 4776 0 1 3170
box -8 -3 16 105
use FILL  FILL_3794
timestamp 1677677812
transform 1 0 4784 0 1 3170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_31
timestamp 1677677812
transform 1 0 4819 0 1 3170
box -10 -3 10 3
use M3_M2  M3_M2_2951
timestamp 1677677812
transform 1 0 164 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3300
timestamp 1677677812
transform 1 0 84 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2984
timestamp 1677677812
transform 1 0 132 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2985
timestamp 1677677812
transform 1 0 172 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2952
timestamp 1677677812
transform 1 0 204 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3301
timestamp 1677677812
transform 1 0 196 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3302
timestamp 1677677812
transform 1 0 204 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3303
timestamp 1677677812
transform 1 0 220 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3391
timestamp 1677677812
transform 1 0 132 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3392
timestamp 1677677812
transform 1 0 164 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3393
timestamp 1677677812
transform 1 0 180 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3394
timestamp 1677677812
transform 1 0 188 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3395
timestamp 1677677812
transform 1 0 212 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2996
timestamp 1677677812
transform 1 0 220 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_3043
timestamp 1677677812
transform 1 0 212 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2953
timestamp 1677677812
transform 1 0 260 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3396
timestamp 1677677812
transform 1 0 252 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3009
timestamp 1677677812
transform 1 0 252 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3044
timestamp 1677677812
transform 1 0 244 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2910
timestamp 1677677812
transform 1 0 284 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3304
timestamp 1677677812
transform 1 0 276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3305
timestamp 1677677812
transform 1 0 284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3306
timestamp 1677677812
transform 1 0 300 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3397
timestamp 1677677812
transform 1 0 268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3398
timestamp 1677677812
transform 1 0 292 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3399
timestamp 1677677812
transform 1 0 308 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3010
timestamp 1677677812
transform 1 0 308 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3065
timestamp 1677677812
transform 1 0 308 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2911
timestamp 1677677812
transform 1 0 332 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2912
timestamp 1677677812
transform 1 0 348 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2954
timestamp 1677677812
transform 1 0 340 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3307
timestamp 1677677812
transform 1 0 340 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2997
timestamp 1677677812
transform 1 0 340 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3308
timestamp 1677677812
transform 1 0 372 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3309
timestamp 1677677812
transform 1 0 380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3400
timestamp 1677677812
transform 1 0 348 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3401
timestamp 1677677812
transform 1 0 364 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2998
timestamp 1677677812
transform 1 0 372 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3402
timestamp 1677677812
transform 1 0 404 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3011
timestamp 1677677812
transform 1 0 404 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3403
timestamp 1677677812
transform 1 0 420 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2955
timestamp 1677677812
transform 1 0 436 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3310
timestamp 1677677812
transform 1 0 436 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2956
timestamp 1677677812
transform 1 0 468 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3311
timestamp 1677677812
transform 1 0 484 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3404
timestamp 1677677812
transform 1 0 460 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3405
timestamp 1677677812
transform 1 0 476 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3406
timestamp 1677677812
transform 1 0 492 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3407
timestamp 1677677812
transform 1 0 500 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3045
timestamp 1677677812
transform 1 0 460 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3012
timestamp 1677677812
transform 1 0 492 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3013
timestamp 1677677812
transform 1 0 508 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3408
timestamp 1677677812
transform 1 0 548 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2913
timestamp 1677677812
transform 1 0 596 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3312
timestamp 1677677812
transform 1 0 572 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3313
timestamp 1677677812
transform 1 0 580 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3314
timestamp 1677677812
transform 1 0 612 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3409
timestamp 1677677812
transform 1 0 580 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3410
timestamp 1677677812
transform 1 0 596 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3411
timestamp 1677677812
transform 1 0 612 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3014
timestamp 1677677812
transform 1 0 572 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3015
timestamp 1677677812
transform 1 0 596 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3016
timestamp 1677677812
transform 1 0 612 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3046
timestamp 1677677812
transform 1 0 612 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3017
timestamp 1677677812
transform 1 0 628 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2914
timestamp 1677677812
transform 1 0 644 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2886
timestamp 1677677812
transform 1 0 724 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2915
timestamp 1677677812
transform 1 0 676 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2957
timestamp 1677677812
transform 1 0 684 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3315
timestamp 1677677812
transform 1 0 660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3412
timestamp 1677677812
transform 1 0 708 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3047
timestamp 1677677812
transform 1 0 660 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3048
timestamp 1677677812
transform 1 0 724 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2887
timestamp 1677677812
transform 1 0 780 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2916
timestamp 1677677812
transform 1 0 772 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2958
timestamp 1677677812
transform 1 0 780 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3316
timestamp 1677677812
transform 1 0 772 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2959
timestamp 1677677812
transform 1 0 812 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3317
timestamp 1677677812
transform 1 0 812 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3413
timestamp 1677677812
transform 1 0 780 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3414
timestamp 1677677812
transform 1 0 788 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3415
timestamp 1677677812
transform 1 0 804 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3066
timestamp 1677677812
transform 1 0 788 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3416
timestamp 1677677812
transform 1 0 828 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3067
timestamp 1677677812
transform 1 0 828 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2888
timestamp 1677677812
transform 1 0 884 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3417
timestamp 1677677812
transform 1 0 884 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2889
timestamp 1677677812
transform 1 0 924 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3418
timestamp 1677677812
transform 1 0 924 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3018
timestamp 1677677812
transform 1 0 924 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3504
timestamp 1677677812
transform 1 0 948 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3049
timestamp 1677677812
transform 1 0 948 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3318
timestamp 1677677812
transform 1 0 964 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2917
timestamp 1677677812
transform 1 0 996 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3319
timestamp 1677677812
transform 1 0 996 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2986
timestamp 1677677812
transform 1 0 1020 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3419
timestamp 1677677812
transform 1 0 988 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3420
timestamp 1677677812
transform 1 0 1004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3421
timestamp 1677677812
transform 1 0 1020 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3068
timestamp 1677677812
transform 1 0 1020 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2987
timestamp 1677677812
transform 1 0 1036 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2918
timestamp 1677677812
transform 1 0 1060 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3320
timestamp 1677677812
transform 1 0 1060 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2919
timestamp 1677677812
transform 1 0 1092 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2988
timestamp 1677677812
transform 1 0 1108 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3422
timestamp 1677677812
transform 1 0 1108 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2989
timestamp 1677677812
transform 1 0 1156 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3423
timestamp 1677677812
transform 1 0 1196 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3321
timestamp 1677677812
transform 1 0 1212 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3050
timestamp 1677677812
transform 1 0 1212 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2890
timestamp 1677677812
transform 1 0 1236 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2960
timestamp 1677677812
transform 1 0 1236 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2990
timestamp 1677677812
transform 1 0 1228 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3505
timestamp 1677677812
transform 1 0 1236 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3506
timestamp 1677677812
transform 1 0 1260 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3082
timestamp 1677677812
transform 1 0 1260 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2891
timestamp 1677677812
transform 1 0 1276 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2991
timestamp 1677677812
transform 1 0 1284 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3424
timestamp 1677677812
transform 1 0 1284 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2920
timestamp 1677677812
transform 1 0 1316 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2961
timestamp 1677677812
transform 1 0 1324 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3322
timestamp 1677677812
transform 1 0 1316 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3323
timestamp 1677677812
transform 1 0 1324 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3507
timestamp 1677677812
transform 1 0 1308 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3508
timestamp 1677677812
transform 1 0 1340 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_2892
timestamp 1677677812
transform 1 0 1348 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2992
timestamp 1677677812
transform 1 0 1364 0 1 3135
box -3 -3 3 3
use M2_M1  M2_M1_3425
timestamp 1677677812
transform 1 0 1364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3426
timestamp 1677677812
transform 1 0 1412 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2893
timestamp 1677677812
transform 1 0 1436 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2962
timestamp 1677677812
transform 1 0 1428 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3324
timestamp 1677677812
transform 1 0 1420 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2921
timestamp 1677677812
transform 1 0 1452 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3427
timestamp 1677677812
transform 1 0 1452 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2963
timestamp 1677677812
transform 1 0 1508 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_3069
timestamp 1677677812
transform 1 0 1508 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2894
timestamp 1677677812
transform 1 0 1532 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2922
timestamp 1677677812
transform 1 0 1548 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2993
timestamp 1677677812
transform 1 0 1540 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2895
timestamp 1677677812
transform 1 0 1588 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2964
timestamp 1677677812
transform 1 0 1556 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2965
timestamp 1677677812
transform 1 0 1580 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3325
timestamp 1677677812
transform 1 0 1548 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3326
timestamp 1677677812
transform 1 0 1556 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3327
timestamp 1677677812
transform 1 0 1572 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3328
timestamp 1677677812
transform 1 0 1588 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3428
timestamp 1677677812
transform 1 0 1548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3429
timestamp 1677677812
transform 1 0 1564 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3430
timestamp 1677677812
transform 1 0 1580 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3431
timestamp 1677677812
transform 1 0 1604 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3051
timestamp 1677677812
transform 1 0 1612 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3070
timestamp 1677677812
transform 1 0 1604 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2923
timestamp 1677677812
transform 1 0 1708 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2966
timestamp 1677677812
transform 1 0 1652 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3329
timestamp 1677677812
transform 1 0 1628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3432
timestamp 1677677812
transform 1 0 1652 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3433
timestamp 1677677812
transform 1 0 1708 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2967
timestamp 1677677812
transform 1 0 1788 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2999
timestamp 1677677812
transform 1 0 1780 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2924
timestamp 1677677812
transform 1 0 1876 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3330
timestamp 1677677812
transform 1 0 1868 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3434
timestamp 1677677812
transform 1 0 1788 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3435
timestamp 1677677812
transform 1 0 1844 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3071
timestamp 1677677812
transform 1 0 1828 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3072
timestamp 1677677812
transform 1 0 1852 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2925
timestamp 1677677812
transform 1 0 1924 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2968
timestamp 1677677812
transform 1 0 1932 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3331
timestamp 1677677812
transform 1 0 1916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3332
timestamp 1677677812
transform 1 0 1932 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3436
timestamp 1677677812
transform 1 0 1908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3437
timestamp 1677677812
transform 1 0 1924 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3438
timestamp 1677677812
transform 1 0 1940 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3073
timestamp 1677677812
transform 1 0 1908 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3333
timestamp 1677677812
transform 1 0 1980 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3019
timestamp 1677677812
transform 1 0 1980 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3334
timestamp 1677677812
transform 1 0 2012 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3335
timestamp 1677677812
transform 1 0 2020 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3336
timestamp 1677677812
transform 1 0 2036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3337
timestamp 1677677812
transform 1 0 2052 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3439
timestamp 1677677812
transform 1 0 2004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3440
timestamp 1677677812
transform 1 0 2012 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3441
timestamp 1677677812
transform 1 0 2028 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3442
timestamp 1677677812
transform 1 0 2044 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3020
timestamp 1677677812
transform 1 0 2028 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3443
timestamp 1677677812
transform 1 0 2076 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3338
timestamp 1677677812
transform 1 0 2108 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2969
timestamp 1677677812
transform 1 0 2132 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3339
timestamp 1677677812
transform 1 0 2132 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3340
timestamp 1677677812
transform 1 0 2148 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3341
timestamp 1677677812
transform 1 0 2156 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3000
timestamp 1677677812
transform 1 0 2132 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3444
timestamp 1677677812
transform 1 0 2140 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3021
timestamp 1677677812
transform 1 0 2116 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3022
timestamp 1677677812
transform 1 0 2140 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3023
timestamp 1677677812
transform 1 0 2188 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2926
timestamp 1677677812
transform 1 0 2212 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2927
timestamp 1677677812
transform 1 0 2236 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3342
timestamp 1677677812
transform 1 0 2236 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3445
timestamp 1677677812
transform 1 0 2220 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3001
timestamp 1677677812
transform 1 0 2236 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3446
timestamp 1677677812
transform 1 0 2268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3447
timestamp 1677677812
transform 1 0 2316 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3024
timestamp 1677677812
transform 1 0 2260 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3343
timestamp 1677677812
transform 1 0 2340 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3002
timestamp 1677677812
transform 1 0 2340 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2928
timestamp 1677677812
transform 1 0 2428 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3448
timestamp 1677677812
transform 1 0 2364 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3449
timestamp 1677677812
transform 1 0 2420 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2929
timestamp 1677677812
transform 1 0 2460 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3344
timestamp 1677677812
transform 1 0 2460 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3025
timestamp 1677677812
transform 1 0 2460 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3345
timestamp 1677677812
transform 1 0 2476 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3074
timestamp 1677677812
transform 1 0 2476 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3450
timestamp 1677677812
transform 1 0 2500 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3075
timestamp 1677677812
transform 1 0 2500 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3346
timestamp 1677677812
transform 1 0 2516 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3347
timestamp 1677677812
transform 1 0 2540 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3348
timestamp 1677677812
transform 1 0 2628 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3451
timestamp 1677677812
transform 1 0 2524 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3452
timestamp 1677677812
transform 1 0 2540 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3453
timestamp 1677677812
transform 1 0 2548 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3454
timestamp 1677677812
transform 1 0 2580 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3026
timestamp 1677677812
transform 1 0 2524 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3076
timestamp 1677677812
transform 1 0 2580 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3455
timestamp 1677677812
transform 1 0 2644 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3027
timestamp 1677677812
transform 1 0 2644 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3349
timestamp 1677677812
transform 1 0 2660 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3350
timestamp 1677677812
transform 1 0 2700 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2930
timestamp 1677677812
transform 1 0 2716 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2931
timestamp 1677677812
transform 1 0 2748 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3351
timestamp 1677677812
transform 1 0 2716 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3456
timestamp 1677677812
transform 1 0 2676 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3457
timestamp 1677677812
transform 1 0 2692 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3003
timestamp 1677677812
transform 1 0 2700 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3458
timestamp 1677677812
transform 1 0 2740 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3004
timestamp 1677677812
transform 1 0 2788 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2932
timestamp 1677677812
transform 1 0 2836 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2970
timestamp 1677677812
transform 1 0 2828 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3459
timestamp 1677677812
transform 1 0 2796 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3460
timestamp 1677677812
transform 1 0 2812 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3298
timestamp 1677677812
transform 1 0 2844 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3352
timestamp 1677677812
transform 1 0 2844 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3509
timestamp 1677677812
transform 1 0 2836 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3028
timestamp 1677677812
transform 1 0 2844 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3299
timestamp 1677677812
transform 1 0 2868 0 1 3145
box -2 -2 2 2
use M2_M1  M2_M1_3353
timestamp 1677677812
transform 1 0 2860 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3005
timestamp 1677677812
transform 1 0 2860 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2971
timestamp 1677677812
transform 1 0 2884 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3354
timestamp 1677677812
transform 1 0 2884 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3461
timestamp 1677677812
transform 1 0 2868 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3029
timestamp 1677677812
transform 1 0 2868 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3462
timestamp 1677677812
transform 1 0 2892 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3355
timestamp 1677677812
transform 1 0 2908 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3510
timestamp 1677677812
transform 1 0 2932 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_2933
timestamp 1677677812
transform 1 0 2964 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3356
timestamp 1677677812
transform 1 0 2956 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3357
timestamp 1677677812
transform 1 0 2964 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3077
timestamp 1677677812
transform 1 0 2956 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3511
timestamp 1677677812
transform 1 0 2972 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_2896
timestamp 1677677812
transform 1 0 2996 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3358
timestamp 1677677812
transform 1 0 3036 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3359
timestamp 1677677812
transform 1 0 3044 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3463
timestamp 1677677812
transform 1 0 3004 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3464
timestamp 1677677812
transform 1 0 3020 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3465
timestamp 1677677812
transform 1 0 3028 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2897
timestamp 1677677812
transform 1 0 3084 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3360
timestamp 1677677812
transform 1 0 3068 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3361
timestamp 1677677812
transform 1 0 3084 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3362
timestamp 1677677812
transform 1 0 3100 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3466
timestamp 1677677812
transform 1 0 3076 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3467
timestamp 1677677812
transform 1 0 3092 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3030
timestamp 1677677812
transform 1 0 3084 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3078
timestamp 1677677812
transform 1 0 3092 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2994
timestamp 1677677812
transform 1 0 3124 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_2934
timestamp 1677677812
transform 1 0 3140 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3363
timestamp 1677677812
transform 1 0 3140 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3468
timestamp 1677677812
transform 1 0 3164 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3031
timestamp 1677677812
transform 1 0 3164 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3052
timestamp 1677677812
transform 1 0 3188 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3053
timestamp 1677677812
transform 1 0 3212 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2935
timestamp 1677677812
transform 1 0 3228 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_3032
timestamp 1677677812
transform 1 0 3228 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2898
timestamp 1677677812
transform 1 0 3244 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3469
timestamp 1677677812
transform 1 0 3260 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3079
timestamp 1677677812
transform 1 0 3260 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_2899
timestamp 1677677812
transform 1 0 3300 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2936
timestamp 1677677812
transform 1 0 3284 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2937
timestamp 1677677812
transform 1 0 3308 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3364
timestamp 1677677812
transform 1 0 3284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3470
timestamp 1677677812
transform 1 0 3308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3471
timestamp 1677677812
transform 1 0 3364 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3033
timestamp 1677677812
transform 1 0 3284 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3512
timestamp 1677677812
transform 1 0 3372 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_2938
timestamp 1677677812
transform 1 0 3412 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3472
timestamp 1677677812
transform 1 0 3412 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3513
timestamp 1677677812
transform 1 0 3420 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3518
timestamp 1677677812
transform 1 0 3404 0 1 3105
box -2 -2 2 2
use M3_M2  M3_M2_3083
timestamp 1677677812
transform 1 0 3404 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3054
timestamp 1677677812
transform 1 0 3444 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3080
timestamp 1677677812
transform 1 0 3460 0 1 3095
box -3 -3 3 3
use M2_M1  M2_M1_3473
timestamp 1677677812
transform 1 0 3492 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2900
timestamp 1677677812
transform 1 0 3524 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3365
timestamp 1677677812
transform 1 0 3516 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3474
timestamp 1677677812
transform 1 0 3524 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3034
timestamp 1677677812
transform 1 0 3516 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3366
timestamp 1677677812
transform 1 0 3548 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2901
timestamp 1677677812
transform 1 0 3564 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3367
timestamp 1677677812
transform 1 0 3580 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2995
timestamp 1677677812
transform 1 0 3596 0 1 3135
box -3 -3 3 3
use M3_M2  M3_M2_3035
timestamp 1677677812
transform 1 0 3604 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3475
timestamp 1677677812
transform 1 0 3620 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3476
timestamp 1677677812
transform 1 0 3628 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3036
timestamp 1677677812
transform 1 0 3628 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3514
timestamp 1677677812
transform 1 0 3636 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3055
timestamp 1677677812
transform 1 0 3636 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2972
timestamp 1677677812
transform 1 0 3684 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3519
timestamp 1677677812
transform 1 0 3684 0 1 3105
box -2 -2 2 2
use M2_M1  M2_M1_3520
timestamp 1677677812
transform 1 0 3740 0 1 3105
box -2 -2 2 2
use M3_M2  M3_M2_3006
timestamp 1677677812
transform 1 0 3764 0 1 3125
box -3 -3 3 3
use M3_M2  M3_M2_2939
timestamp 1677677812
transform 1 0 3780 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2940
timestamp 1677677812
transform 1 0 3820 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3368
timestamp 1677677812
transform 1 0 3812 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3477
timestamp 1677677812
transform 1 0 3796 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3007
timestamp 1677677812
transform 1 0 3804 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3515
timestamp 1677677812
transform 1 0 3772 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3516
timestamp 1677677812
transform 1 0 3780 0 1 3115
box -2 -2 2 2
use M3_M2  M3_M2_3056
timestamp 1677677812
transform 1 0 3772 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3037
timestamp 1677677812
transform 1 0 3788 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3517
timestamp 1677677812
transform 1 0 3796 0 1 3115
box -2 -2 2 2
use M2_M1  M2_M1_3521
timestamp 1677677812
transform 1 0 3788 0 1 3105
box -2 -2 2 2
use M3_M2  M3_M2_2902
timestamp 1677677812
transform 1 0 3852 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3369
timestamp 1677677812
transform 1 0 3860 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3370
timestamp 1677677812
transform 1 0 3868 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3478
timestamp 1677677812
transform 1 0 3836 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3479
timestamp 1677677812
transform 1 0 3852 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3480
timestamp 1677677812
transform 1 0 3868 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3057
timestamp 1677677812
transform 1 0 3844 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3058
timestamp 1677677812
transform 1 0 3860 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2941
timestamp 1677677812
transform 1 0 3884 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3481
timestamp 1677677812
transform 1 0 3884 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3059
timestamp 1677677812
transform 1 0 3884 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2903
timestamp 1677677812
transform 1 0 3900 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2942
timestamp 1677677812
transform 1 0 3908 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2904
timestamp 1677677812
transform 1 0 3940 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2973
timestamp 1677677812
transform 1 0 3932 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2943
timestamp 1677677812
transform 1 0 3956 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3371
timestamp 1677677812
transform 1 0 3908 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3372
timestamp 1677677812
transform 1 0 3916 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3373
timestamp 1677677812
transform 1 0 3932 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3374
timestamp 1677677812
transform 1 0 3948 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3482
timestamp 1677677812
transform 1 0 3908 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3483
timestamp 1677677812
transform 1 0 3924 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3484
timestamp 1677677812
transform 1 0 3940 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3485
timestamp 1677677812
transform 1 0 3956 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2974
timestamp 1677677812
transform 1 0 4036 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2975
timestamp 1677677812
transform 1 0 4060 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3375
timestamp 1677677812
transform 1 0 4076 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3486
timestamp 1677677812
transform 1 0 4036 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3060
timestamp 1677677812
transform 1 0 4012 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2905
timestamp 1677677812
transform 1 0 4108 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2944
timestamp 1677677812
transform 1 0 4116 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2976
timestamp 1677677812
transform 1 0 4116 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2977
timestamp 1677677812
transform 1 0 4156 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3376
timestamp 1677677812
transform 1 0 4116 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3487
timestamp 1677677812
transform 1 0 4156 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3488
timestamp 1677677812
transform 1 0 4196 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_2906
timestamp 1677677812
transform 1 0 4212 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2945
timestamp 1677677812
transform 1 0 4212 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3377
timestamp 1677677812
transform 1 0 4228 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2946
timestamp 1677677812
transform 1 0 4260 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2978
timestamp 1677677812
transform 1 0 4260 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2947
timestamp 1677677812
transform 1 0 4284 0 1 3155
box -3 -3 3 3
use M2_M1  M2_M1_3378
timestamp 1677677812
transform 1 0 4260 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3379
timestamp 1677677812
transform 1 0 4276 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3380
timestamp 1677677812
transform 1 0 4284 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3489
timestamp 1677677812
transform 1 0 4252 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3490
timestamp 1677677812
transform 1 0 4268 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3491
timestamp 1677677812
transform 1 0 4276 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3061
timestamp 1677677812
transform 1 0 4268 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3084
timestamp 1677677812
transform 1 0 4268 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2907
timestamp 1677677812
transform 1 0 4308 0 1 3165
box -3 -3 3 3
use M2_M1  M2_M1_3492
timestamp 1677677812
transform 1 0 4308 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3381
timestamp 1677677812
transform 1 0 4324 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3493
timestamp 1677677812
transform 1 0 4332 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3494
timestamp 1677677812
transform 1 0 4348 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3495
timestamp 1677677812
transform 1 0 4356 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3038
timestamp 1677677812
transform 1 0 4340 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3062
timestamp 1677677812
transform 1 0 4324 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_3085
timestamp 1677677812
transform 1 0 4356 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_2948
timestamp 1677677812
transform 1 0 4380 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2979
timestamp 1677677812
transform 1 0 4388 0 1 3145
box -3 -3 3 3
use M3_M2  M3_M2_2980
timestamp 1677677812
transform 1 0 4404 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3382
timestamp 1677677812
transform 1 0 4380 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3383
timestamp 1677677812
transform 1 0 4388 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3384
timestamp 1677677812
transform 1 0 4404 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3385
timestamp 1677677812
transform 1 0 4420 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3496
timestamp 1677677812
transform 1 0 4396 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3497
timestamp 1677677812
transform 1 0 4412 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3039
timestamp 1677677812
transform 1 0 4388 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3063
timestamp 1677677812
transform 1 0 4412 0 1 3105
box -3 -3 3 3
use M3_M2  M3_M2_2908
timestamp 1677677812
transform 1 0 4468 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2909
timestamp 1677677812
transform 1 0 4492 0 1 3165
box -3 -3 3 3
use M3_M2  M3_M2_2981
timestamp 1677677812
transform 1 0 4492 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3386
timestamp 1677677812
transform 1 0 4468 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3498
timestamp 1677677812
transform 1 0 4492 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3040
timestamp 1677677812
transform 1 0 4500 0 1 3115
box -3 -3 3 3
use M2_M1  M2_M1_3499
timestamp 1677677812
transform 1 0 4572 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3500
timestamp 1677677812
transform 1 0 4580 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3064
timestamp 1677677812
transform 1 0 4572 0 1 3105
box -3 -3 3 3
use M2_M1  M2_M1_3387
timestamp 1677677812
transform 1 0 4596 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_2949
timestamp 1677677812
transform 1 0 4628 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2982
timestamp 1677677812
transform 1 0 4620 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3388
timestamp 1677677812
transform 1 0 4620 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3389
timestamp 1677677812
transform 1 0 4636 0 1 3135
box -2 -2 2 2
use M3_M2  M3_M2_3008
timestamp 1677677812
transform 1 0 4604 0 1 3125
box -3 -3 3 3
use M2_M1  M2_M1_3501
timestamp 1677677812
transform 1 0 4628 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3041
timestamp 1677677812
transform 1 0 4596 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_3042
timestamp 1677677812
transform 1 0 4668 0 1 3115
box -3 -3 3 3
use M3_M2  M3_M2_2950
timestamp 1677677812
transform 1 0 4756 0 1 3155
box -3 -3 3 3
use M3_M2  M3_M2_2983
timestamp 1677677812
transform 1 0 4708 0 1 3145
box -3 -3 3 3
use M2_M1  M2_M1_3390
timestamp 1677677812
transform 1 0 4684 0 1 3135
box -2 -2 2 2
use M2_M1  M2_M1_3502
timestamp 1677677812
transform 1 0 4708 0 1 3125
box -2 -2 2 2
use M2_M1  M2_M1_3503
timestamp 1677677812
transform 1 0 4764 0 1 3125
box -2 -2 2 2
use M3_M2  M3_M2_3081
timestamp 1677677812
transform 1 0 4764 0 1 3095
box -3 -3 3 3
use M3_M2  M3_M2_3086
timestamp 1677677812
transform 1 0 4740 0 1 3085
box -3 -3 3 3
use M3_M2  M3_M2_3087
timestamp 1677677812
transform 1 0 4772 0 1 3085
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_32
timestamp 1677677812
transform 1 0 24 0 1 3070
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_218
timestamp 1677677812
transform 1 0 72 0 -1 3170
box -8 -3 104 105
use INVX2  INVX2_245
timestamp 1677677812
transform -1 0 184 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3232
timestamp 1677677812
transform 1 0 184 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_139
timestamp 1677677812
transform -1 0 232 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3233
timestamp 1677677812
transform 1 0 232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3235
timestamp 1677677812
transform 1 0 240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3242
timestamp 1677677812
transform 1 0 248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3243
timestamp 1677677812
transform 1 0 256 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3244
timestamp 1677677812
transform 1 0 264 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_140
timestamp 1677677812
transform -1 0 312 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3245
timestamp 1677677812
transform 1 0 312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3246
timestamp 1677677812
transform 1 0 320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3247
timestamp 1677677812
transform 1 0 328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3248
timestamp 1677677812
transform 1 0 336 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_141
timestamp 1677677812
transform 1 0 344 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3249
timestamp 1677677812
transform 1 0 384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3250
timestamp 1677677812
transform 1 0 392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3251
timestamp 1677677812
transform 1 0 400 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_247
timestamp 1677677812
transform 1 0 408 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3252
timestamp 1677677812
transform 1 0 424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3253
timestamp 1677677812
transform 1 0 432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3254
timestamp 1677677812
transform 1 0 440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3255
timestamp 1677677812
transform 1 0 448 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_142
timestamp 1677677812
transform 1 0 456 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3256
timestamp 1677677812
transform 1 0 496 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3258
timestamp 1677677812
transform 1 0 504 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3259
timestamp 1677677812
transform 1 0 512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3260
timestamp 1677677812
transform 1 0 520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3268
timestamp 1677677812
transform 1 0 528 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_249
timestamp 1677677812
transform -1 0 552 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3269
timestamp 1677677812
transform 1 0 552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3270
timestamp 1677677812
transform 1 0 560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3271
timestamp 1677677812
transform 1 0 568 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_144
timestamp 1677677812
transform -1 0 616 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3272
timestamp 1677677812
transform 1 0 616 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3274
timestamp 1677677812
transform 1 0 624 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3276
timestamp 1677677812
transform 1 0 632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3278
timestamp 1677677812
transform 1 0 640 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_221
timestamp 1677677812
transform 1 0 648 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3287
timestamp 1677677812
transform 1 0 744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3289
timestamp 1677677812
transform 1 0 752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3291
timestamp 1677677812
transform 1 0 760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3295
timestamp 1677677812
transform 1 0 768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3296
timestamp 1677677812
transform 1 0 776 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_146
timestamp 1677677812
transform 1 0 784 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3297
timestamp 1677677812
transform 1 0 824 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3299
timestamp 1677677812
transform 1 0 832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3301
timestamp 1677677812
transform 1 0 840 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3303
timestamp 1677677812
transform 1 0 848 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3305
timestamp 1677677812
transform 1 0 856 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3307
timestamp 1677677812
transform 1 0 864 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3312
timestamp 1677677812
transform 1 0 872 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3313
timestamp 1677677812
transform 1 0 880 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_71
timestamp 1677677812
transform 1 0 888 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3314
timestamp 1677677812
transform 1 0 920 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3316
timestamp 1677677812
transform 1 0 928 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3318
timestamp 1677677812
transform 1 0 936 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3319
timestamp 1677677812
transform 1 0 944 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3320
timestamp 1677677812
transform 1 0 952 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3321
timestamp 1677677812
transform 1 0 960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3322
timestamp 1677677812
transform 1 0 968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3324
timestamp 1677677812
transform 1 0 976 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_147
timestamp 1677677812
transform 1 0 984 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3329
timestamp 1677677812
transform 1 0 1024 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3330
timestamp 1677677812
transform 1 0 1032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3332
timestamp 1677677812
transform 1 0 1040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3334
timestamp 1677677812
transform 1 0 1048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3336
timestamp 1677677812
transform 1 0 1056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3338
timestamp 1677677812
transform 1 0 1064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3342
timestamp 1677677812
transform 1 0 1072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3343
timestamp 1677677812
transform 1 0 1080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3344
timestamp 1677677812
transform 1 0 1088 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_73
timestamp 1677677812
transform 1 0 1096 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3345
timestamp 1677677812
transform 1 0 1128 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3347
timestamp 1677677812
transform 1 0 1136 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3349
timestamp 1677677812
transform 1 0 1144 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3351
timestamp 1677677812
transform 1 0 1152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3354
timestamp 1677677812
transform 1 0 1160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3355
timestamp 1677677812
transform 1 0 1168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3356
timestamp 1677677812
transform 1 0 1176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3357
timestamp 1677677812
transform 1 0 1184 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3358
timestamp 1677677812
transform 1 0 1192 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3359
timestamp 1677677812
transform 1 0 1200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3360
timestamp 1677677812
transform 1 0 1208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3362
timestamp 1677677812
transform 1 0 1216 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3364
timestamp 1677677812
transform 1 0 1224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3366
timestamp 1677677812
transform 1 0 1232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3371
timestamp 1677677812
transform 1 0 1240 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3372
timestamp 1677677812
transform 1 0 1248 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3373
timestamp 1677677812
transform 1 0 1256 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_75
timestamp 1677677812
transform -1 0 1296 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3374
timestamp 1677677812
transform 1 0 1296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3376
timestamp 1677677812
transform 1 0 1304 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3378
timestamp 1677677812
transform 1 0 1312 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3383
timestamp 1677677812
transform 1 0 1320 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3384
timestamp 1677677812
transform 1 0 1328 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3385
timestamp 1677677812
transform 1 0 1336 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_77
timestamp 1677677812
transform -1 0 1376 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3386
timestamp 1677677812
transform 1 0 1376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3388
timestamp 1677677812
transform 1 0 1384 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3390
timestamp 1677677812
transform 1 0 1392 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3392
timestamp 1677677812
transform 1 0 1400 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3394
timestamp 1677677812
transform 1 0 1408 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3397
timestamp 1677677812
transform 1 0 1416 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_250
timestamp 1677677812
transform 1 0 1424 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3398
timestamp 1677677812
transform 1 0 1440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3399
timestamp 1677677812
transform 1 0 1448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3400
timestamp 1677677812
transform 1 0 1456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3401
timestamp 1677677812
transform 1 0 1464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3403
timestamp 1677677812
transform 1 0 1472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3405
timestamp 1677677812
transform 1 0 1480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3410
timestamp 1677677812
transform 1 0 1488 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_251
timestamp 1677677812
transform -1 0 1512 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3411
timestamp 1677677812
transform 1 0 1512 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3413
timestamp 1677677812
transform 1 0 1520 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3415
timestamp 1677677812
transform 1 0 1528 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3419
timestamp 1677677812
transform 1 0 1536 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3420
timestamp 1677677812
transform 1 0 1544 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_140
timestamp 1677677812
transform -1 0 1592 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3421
timestamp 1677677812
transform 1 0 1592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3423
timestamp 1677677812
transform 1 0 1600 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3425
timestamp 1677677812
transform 1 0 1608 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_222
timestamp 1677677812
transform 1 0 1616 0 -1 3170
box -8 -3 104 105
use M3_M2  M3_M2_3088
timestamp 1677677812
transform 1 0 1724 0 1 3075
box -3 -3 3 3
use FILL  FILL_3436
timestamp 1677677812
transform 1 0 1712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3438
timestamp 1677677812
transform 1 0 1720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3440
timestamp 1677677812
transform 1 0 1728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3441
timestamp 1677677812
transform 1 0 1736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3442
timestamp 1677677812
transform 1 0 1744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3443
timestamp 1677677812
transform 1 0 1752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3445
timestamp 1677677812
transform 1 0 1760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3447
timestamp 1677677812
transform 1 0 1768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3457
timestamp 1677677812
transform 1 0 1776 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_223
timestamp 1677677812
transform -1 0 1880 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3458
timestamp 1677677812
transform 1 0 1880 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3460
timestamp 1677677812
transform 1 0 1888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3463
timestamp 1677677812
transform 1 0 1896 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_151
timestamp 1677677812
transform 1 0 1904 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3464
timestamp 1677677812
transform 1 0 1944 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3466
timestamp 1677677812
transform 1 0 1952 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3468
timestamp 1677677812
transform 1 0 1960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3470
timestamp 1677677812
transform 1 0 1968 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_253
timestamp 1677677812
transform 1 0 1976 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3474
timestamp 1677677812
transform 1 0 1992 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3476
timestamp 1677677812
transform 1 0 2000 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_152
timestamp 1677677812
transform 1 0 2008 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3483
timestamp 1677677812
transform 1 0 2048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3485
timestamp 1677677812
transform 1 0 2056 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3487
timestamp 1677677812
transform 1 0 2064 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3494
timestamp 1677677812
transform 1 0 2072 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3495
timestamp 1677677812
transform 1 0 2080 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3496
timestamp 1677677812
transform 1 0 2088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3497
timestamp 1677677812
transform 1 0 2096 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3498
timestamp 1677677812
transform 1 0 2104 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_141
timestamp 1677677812
transform 1 0 2112 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3499
timestamp 1677677812
transform 1 0 2152 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3501
timestamp 1677677812
transform 1 0 2160 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3503
timestamp 1677677812
transform 1 0 2168 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3505
timestamp 1677677812
transform 1 0 2176 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3516
timestamp 1677677812
transform 1 0 2184 0 -1 3170
box -8 -3 16 105
use BUFX2  BUFX2_26
timestamp 1677677812
transform -1 0 2216 0 -1 3170
box -5 -3 28 105
use FILL  FILL_3517
timestamp 1677677812
transform 1 0 2216 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_224
timestamp 1677677812
transform 1 0 2224 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3518
timestamp 1677677812
transform 1 0 2320 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_225
timestamp 1677677812
transform 1 0 2328 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3525
timestamp 1677677812
transform 1 0 2424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3527
timestamp 1677677812
transform 1 0 2432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3529
timestamp 1677677812
transform 1 0 2440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3531
timestamp 1677677812
transform 1 0 2448 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_255
timestamp 1677677812
transform 1 0 2456 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3532
timestamp 1677677812
transform 1 0 2472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3533
timestamp 1677677812
transform 1 0 2480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3534
timestamp 1677677812
transform 1 0 2488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3536
timestamp 1677677812
transform 1 0 2496 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_155
timestamp 1677677812
transform 1 0 2504 0 -1 3170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_226
timestamp 1677677812
transform -1 0 2640 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3548
timestamp 1677677812
transform 1 0 2640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3551
timestamp 1677677812
transform 1 0 2648 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_157
timestamp 1677677812
transform 1 0 2656 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3552
timestamp 1677677812
transform 1 0 2696 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_228
timestamp 1677677812
transform 1 0 2704 0 -1 3170
box -8 -3 104 105
use OAI21X1  OAI21X1_79
timestamp 1677677812
transform 1 0 2800 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3556
timestamp 1677677812
transform 1 0 2832 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3558
timestamp 1677677812
transform 1 0 2840 0 -1 3170
box -8 -3 16 105
use NOR2X1  NOR2X1_36
timestamp 1677677812
transform 1 0 2848 0 -1 3170
box -8 -3 32 105
use NOR2X1  NOR2X1_37
timestamp 1677677812
transform 1 0 2872 0 -1 3170
box -8 -3 32 105
use FILL  FILL_3566
timestamp 1677677812
transform 1 0 2896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3572
timestamp 1677677812
transform 1 0 2904 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3573
timestamp 1677677812
transform 1 0 2912 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3574
timestamp 1677677812
transform 1 0 2920 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_80
timestamp 1677677812
transform -1 0 2960 0 -1 3170
box -8 -3 34 105
use FILL  FILL_3575
timestamp 1677677812
transform 1 0 2960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3581
timestamp 1677677812
transform 1 0 2968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3582
timestamp 1677677812
transform 1 0 2976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3583
timestamp 1677677812
transform 1 0 2984 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3584
timestamp 1677677812
transform 1 0 2992 0 -1 3170
box -8 -3 16 105
use OAI21X1  OAI21X1_82
timestamp 1677677812
transform -1 0 3032 0 -1 3170
box -8 -3 34 105
use M3_M2  M3_M2_3089
timestamp 1677677812
transform 1 0 3044 0 1 3075
box -3 -3 3 3
use FILL  FILL_3585
timestamp 1677677812
transform 1 0 3032 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3593
timestamp 1677677812
transform 1 0 3040 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3594
timestamp 1677677812
transform 1 0 3048 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3595
timestamp 1677677812
transform 1 0 3056 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_145
timestamp 1677677812
transform 1 0 3064 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3596
timestamp 1677677812
transform 1 0 3104 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3597
timestamp 1677677812
transform 1 0 3112 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3598
timestamp 1677677812
transform 1 0 3120 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_230
timestamp 1677677812
transform 1 0 3128 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3599
timestamp 1677677812
transform 1 0 3224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3600
timestamp 1677677812
transform 1 0 3232 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3601
timestamp 1677677812
transform 1 0 3240 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_259
timestamp 1677677812
transform 1 0 3248 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3611
timestamp 1677677812
transform 1 0 3264 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_231
timestamp 1677677812
transform 1 0 3272 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3612
timestamp 1677677812
transform 1 0 3368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3616
timestamp 1677677812
transform 1 0 3376 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3617
timestamp 1677677812
transform 1 0 3384 0 -1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_17
timestamp 1677677812
transform -1 0 3424 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3618
timestamp 1677677812
transform 1 0 3424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3620
timestamp 1677677812
transform 1 0 3432 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3622
timestamp 1677677812
transform 1 0 3440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3625
timestamp 1677677812
transform 1 0 3448 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3626
timestamp 1677677812
transform 1 0 3456 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3627
timestamp 1677677812
transform 1 0 3464 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3628
timestamp 1677677812
transform 1 0 3472 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3629
timestamp 1677677812
transform 1 0 3480 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3630
timestamp 1677677812
transform 1 0 3488 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3636
timestamp 1677677812
transform 1 0 3496 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_158
timestamp 1677677812
transform -1 0 3544 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3637
timestamp 1677677812
transform 1 0 3544 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3638
timestamp 1677677812
transform 1 0 3552 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3639
timestamp 1677677812
transform 1 0 3560 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3641
timestamp 1677677812
transform 1 0 3568 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3643
timestamp 1677677812
transform 1 0 3576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3647
timestamp 1677677812
transform 1 0 3584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3648
timestamp 1677677812
transform 1 0 3592 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3649
timestamp 1677677812
transform 1 0 3600 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3090
timestamp 1677677812
transform 1 0 3620 0 1 3075
box -3 -3 3 3
use FILL  FILL_3650
timestamp 1677677812
transform 1 0 3608 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_260
timestamp 1677677812
transform 1 0 3616 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3651
timestamp 1677677812
transform 1 0 3632 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3653
timestamp 1677677812
transform 1 0 3640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3655
timestamp 1677677812
transform 1 0 3648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3657
timestamp 1677677812
transform 1 0 3656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3664
timestamp 1677677812
transform 1 0 3664 0 -1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_21
timestamp 1677677812
transform -1 0 3704 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3665
timestamp 1677677812
transform 1 0 3704 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3667
timestamp 1677677812
transform 1 0 3712 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3669
timestamp 1677677812
transform 1 0 3720 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3670
timestamp 1677677812
transform 1 0 3728 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3671
timestamp 1677677812
transform 1 0 3736 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3673
timestamp 1677677812
transform 1 0 3744 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3675
timestamp 1677677812
transform 1 0 3752 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3677
timestamp 1677677812
transform 1 0 3760 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3691
timestamp 1677677812
transform 1 0 3768 0 -1 3170
box -8 -3 16 105
use NAND3X1  NAND3X1_22
timestamp 1677677812
transform -1 0 3808 0 -1 3170
box -8 -3 40 105
use FILL  FILL_3692
timestamp 1677677812
transform 1 0 3808 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3693
timestamp 1677677812
transform 1 0 3816 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3694
timestamp 1677677812
transform 1 0 3824 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_160
timestamp 1677677812
transform 1 0 3832 0 -1 3170
box -8 -3 46 105
use INVX2  INVX2_263
timestamp 1677677812
transform -1 0 3888 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3695
timestamp 1677677812
transform 1 0 3888 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3696
timestamp 1677677812
transform 1 0 3896 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3697
timestamp 1677677812
transform 1 0 3904 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_148
timestamp 1677677812
transform -1 0 3952 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3698
timestamp 1677677812
transform 1 0 3952 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3699
timestamp 1677677812
transform 1 0 3960 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3701
timestamp 1677677812
transform 1 0 3968 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3703
timestamp 1677677812
transform 1 0 3976 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3719
timestamp 1677677812
transform 1 0 3984 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3091
timestamp 1677677812
transform 1 0 4076 0 1 3075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_232
timestamp 1677677812
transform -1 0 4088 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3720
timestamp 1677677812
transform 1 0 4088 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3721
timestamp 1677677812
transform 1 0 4096 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_233
timestamp 1677677812
transform 1 0 4104 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3722
timestamp 1677677812
transform 1 0 4200 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3723
timestamp 1677677812
transform 1 0 4208 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3725
timestamp 1677677812
transform 1 0 4216 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3727
timestamp 1677677812
transform 1 0 4224 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3729
timestamp 1677677812
transform 1 0 4232 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_151
timestamp 1677677812
transform -1 0 4280 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3731
timestamp 1677677812
transform 1 0 4280 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3733
timestamp 1677677812
transform 1 0 4288 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3735
timestamp 1677677812
transform 1 0 4296 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3737
timestamp 1677677812
transform 1 0 4304 0 -1 3170
box -8 -3 16 105
use AOI22X1  AOI22X1_162
timestamp 1677677812
transform 1 0 4312 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3744
timestamp 1677677812
transform 1 0 4352 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3746
timestamp 1677677812
transform 1 0 4360 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3748
timestamp 1677677812
transform 1 0 4368 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3750
timestamp 1677677812
transform 1 0 4376 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_152
timestamp 1677677812
transform 1 0 4384 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3757
timestamp 1677677812
transform 1 0 4424 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3759
timestamp 1677677812
transform 1 0 4432 0 -1 3170
box -8 -3 16 105
use M3_M2  M3_M2_3092
timestamp 1677677812
transform 1 0 4452 0 1 3075
box -3 -3 3 3
use FILL  FILL_3761
timestamp 1677677812
transform 1 0 4440 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3763
timestamp 1677677812
transform 1 0 4448 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_235
timestamp 1677677812
transform 1 0 4456 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3768
timestamp 1677677812
transform 1 0 4552 0 -1 3170
box -8 -3 16 105
use INVX2  INVX2_266
timestamp 1677677812
transform 1 0 4560 0 -1 3170
box -9 -3 26 105
use FILL  FILL_3769
timestamp 1677677812
transform 1 0 4576 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3771
timestamp 1677677812
transform 1 0 4584 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3773
timestamp 1677677812
transform 1 0 4592 0 -1 3170
box -8 -3 16 105
use OAI22X1  OAI22X1_153
timestamp 1677677812
transform 1 0 4600 0 -1 3170
box -8 -3 46 105
use FILL  FILL_3780
timestamp 1677677812
transform 1 0 4640 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3782
timestamp 1677677812
transform 1 0 4648 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3784
timestamp 1677677812
transform 1 0 4656 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3790
timestamp 1677677812
transform 1 0 4664 0 -1 3170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_236
timestamp 1677677812
transform 1 0 4672 0 -1 3170
box -8 -3 104 105
use FILL  FILL_3791
timestamp 1677677812
transform 1 0 4768 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3793
timestamp 1677677812
transform 1 0 4776 0 -1 3170
box -8 -3 16 105
use FILL  FILL_3795
timestamp 1677677812
transform 1 0 4784 0 -1 3170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_33
timestamp 1677677812
transform 1 0 4843 0 1 3070
box -10 -3 10 3
use M3_M2  M3_M2_3153
timestamp 1677677812
transform 1 0 100 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3645
timestamp 1677677812
transform 1 0 100 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3131
timestamp 1677677812
transform 1 0 116 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3154
timestamp 1677677812
transform 1 0 132 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3530
timestamp 1677677812
transform 1 0 108 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3531
timestamp 1677677812
transform 1 0 116 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3532
timestamp 1677677812
transform 1 0 132 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3190
timestamp 1677677812
transform 1 0 140 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3533
timestamp 1677677812
transform 1 0 148 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3646
timestamp 1677677812
transform 1 0 124 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3647
timestamp 1677677812
transform 1 0 140 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3648
timestamp 1677677812
transform 1 0 148 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3232
timestamp 1677677812
transform 1 0 124 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3233
timestamp 1677677812
transform 1 0 148 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3649
timestamp 1677677812
transform 1 0 164 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3534
timestamp 1677677812
transform 1 0 172 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3132
timestamp 1677677812
transform 1 0 188 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3535
timestamp 1677677812
transform 1 0 188 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3213
timestamp 1677677812
transform 1 0 188 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3650
timestamp 1677677812
transform 1 0 196 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3191
timestamp 1677677812
transform 1 0 220 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3214
timestamp 1677677812
transform 1 0 228 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3155
timestamp 1677677812
transform 1 0 244 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3536
timestamp 1677677812
transform 1 0 244 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3265
timestamp 1677677812
transform 1 0 236 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3101
timestamp 1677677812
transform 1 0 268 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3156
timestamp 1677677812
transform 1 0 284 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3537
timestamp 1677677812
transform 1 0 268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3538
timestamp 1677677812
transform 1 0 284 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3651
timestamp 1677677812
transform 1 0 252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3652
timestamp 1677677812
transform 1 0 260 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3215
timestamp 1677677812
transform 1 0 268 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3102
timestamp 1677677812
transform 1 0 300 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3653
timestamp 1677677812
transform 1 0 276 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3654
timestamp 1677677812
transform 1 0 292 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3234
timestamp 1677677812
transform 1 0 276 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3266
timestamp 1677677812
transform 1 0 300 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3103
timestamp 1677677812
transform 1 0 396 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3157
timestamp 1677677812
transform 1 0 316 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3158
timestamp 1677677812
transform 1 0 364 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3159
timestamp 1677677812
transform 1 0 404 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3192
timestamp 1677677812
transform 1 0 316 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3539
timestamp 1677677812
transform 1 0 364 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3193
timestamp 1677677812
transform 1 0 388 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3540
timestamp 1677677812
transform 1 0 396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3541
timestamp 1677677812
transform 1 0 404 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3655
timestamp 1677677812
transform 1 0 316 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3216
timestamp 1677677812
transform 1 0 340 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3656
timestamp 1677677812
transform 1 0 460 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3104
timestamp 1677677812
transform 1 0 484 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3542
timestamp 1677677812
transform 1 0 500 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3657
timestamp 1677677812
transform 1 0 476 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3543
timestamp 1677677812
transform 1 0 564 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3544
timestamp 1677677812
transform 1 0 620 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3105
timestamp 1677677812
transform 1 0 676 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3133
timestamp 1677677812
transform 1 0 668 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3545
timestamp 1677677812
transform 1 0 644 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3546
timestamp 1677677812
transform 1 0 668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3658
timestamp 1677677812
transform 1 0 660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3659
timestamp 1677677812
transform 1 0 676 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3267
timestamp 1677677812
transform 1 0 660 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3547
timestamp 1677677812
transform 1 0 708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3747
timestamp 1677677812
transform 1 0 772 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3120
timestamp 1677677812
transform 1 0 788 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3160
timestamp 1677677812
transform 1 0 796 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3548
timestamp 1677677812
transform 1 0 804 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3161
timestamp 1677677812
transform 1 0 828 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3660
timestamp 1677677812
transform 1 0 812 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3661
timestamp 1677677812
transform 1 0 820 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3162
timestamp 1677677812
transform 1 0 876 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3549
timestamp 1677677812
transform 1 0 876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3550
timestamp 1677677812
transform 1 0 884 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3163
timestamp 1677677812
transform 1 0 908 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3235
timestamp 1677677812
transform 1 0 900 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3662
timestamp 1677677812
transform 1 0 908 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3217
timestamp 1677677812
transform 1 0 924 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3748
timestamp 1677677812
transform 1 0 924 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3523
timestamp 1677677812
transform 1 0 948 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3194
timestamp 1677677812
transform 1 0 948 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3663
timestamp 1677677812
transform 1 0 948 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3551
timestamp 1677677812
transform 1 0 972 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3552
timestamp 1677677812
transform 1 0 1004 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3164
timestamp 1677677812
transform 1 0 1036 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3553
timestamp 1677677812
transform 1 0 1036 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3093
timestamp 1677677812
transform 1 0 1076 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3094
timestamp 1677677812
transform 1 0 1108 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3165
timestamp 1677677812
transform 1 0 1100 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3554
timestamp 1677677812
transform 1 0 1060 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3555
timestamp 1677677812
transform 1 0 1100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3664
timestamp 1677677812
transform 1 0 1140 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3236
timestamp 1677677812
transform 1 0 1140 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3749
timestamp 1677677812
transform 1 0 1164 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3268
timestamp 1677677812
transform 1 0 1164 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3134
timestamp 1677677812
transform 1 0 1180 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3269
timestamp 1677677812
transform 1 0 1180 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3556
timestamp 1677677812
transform 1 0 1196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3557
timestamp 1677677812
transform 1 0 1260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3558
timestamp 1677677812
transform 1 0 1276 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3195
timestamp 1677677812
transform 1 0 1284 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3665
timestamp 1677677812
transform 1 0 1252 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3666
timestamp 1677677812
transform 1 0 1276 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3667
timestamp 1677677812
transform 1 0 1284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3524
timestamp 1677677812
transform 1 0 1340 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3559
timestamp 1677677812
transform 1 0 1364 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3121
timestamp 1677677812
transform 1 0 1428 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3560
timestamp 1677677812
transform 1 0 1420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3561
timestamp 1677677812
transform 1 0 1452 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3196
timestamp 1677677812
transform 1 0 1500 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3668
timestamp 1677677812
transform 1 0 1412 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3218
timestamp 1677677812
transform 1 0 1420 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3669
timestamp 1677677812
transform 1 0 1500 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3237
timestamp 1677677812
transform 1 0 1484 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3670
timestamp 1677677812
transform 1 0 1516 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3238
timestamp 1677677812
transform 1 0 1524 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3562
timestamp 1677677812
transform 1 0 1548 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3166
timestamp 1677677812
transform 1 0 1564 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3167
timestamp 1677677812
transform 1 0 1580 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3563
timestamp 1677677812
transform 1 0 1564 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3564
timestamp 1677677812
transform 1 0 1588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3671
timestamp 1677677812
transform 1 0 1580 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3672
timestamp 1677677812
transform 1 0 1604 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3197
timestamp 1677677812
transform 1 0 1612 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3198
timestamp 1677677812
transform 1 0 1628 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3135
timestamp 1677677812
transform 1 0 1644 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3136
timestamp 1677677812
transform 1 0 1668 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3168
timestamp 1677677812
transform 1 0 1684 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3565
timestamp 1677677812
transform 1 0 1668 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3566
timestamp 1677677812
transform 1 0 1684 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3219
timestamp 1677677812
transform 1 0 1668 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3673
timestamp 1677677812
transform 1 0 1676 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3567
timestamp 1677677812
transform 1 0 1716 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3674
timestamp 1677677812
transform 1 0 1724 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3568
timestamp 1677677812
transform 1 0 1748 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3675
timestamp 1677677812
transform 1 0 1764 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3676
timestamp 1677677812
transform 1 0 1772 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3239
timestamp 1677677812
transform 1 0 1772 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3270
timestamp 1677677812
transform 1 0 1764 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3271
timestamp 1677677812
transform 1 0 1780 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3569
timestamp 1677677812
transform 1 0 1812 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3570
timestamp 1677677812
transform 1 0 1820 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3571
timestamp 1677677812
transform 1 0 1836 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3677
timestamp 1677677812
transform 1 0 1828 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3678
timestamp 1677677812
transform 1 0 1844 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3240
timestamp 1677677812
transform 1 0 1836 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3272
timestamp 1677677812
transform 1 0 1828 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3199
timestamp 1677677812
transform 1 0 1868 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3169
timestamp 1677677812
transform 1 0 1892 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3572
timestamp 1677677812
transform 1 0 1876 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3679
timestamp 1677677812
transform 1 0 1868 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3200
timestamp 1677677812
transform 1 0 1884 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3573
timestamp 1677677812
transform 1 0 1892 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3574
timestamp 1677677812
transform 1 0 1932 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3680
timestamp 1677677812
transform 1 0 1908 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3681
timestamp 1677677812
transform 1 0 1924 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3220
timestamp 1677677812
transform 1 0 1932 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3682
timestamp 1677677812
transform 1 0 1940 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3241
timestamp 1677677812
transform 1 0 1916 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3273
timestamp 1677677812
transform 1 0 1924 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3242
timestamp 1677677812
transform 1 0 1956 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3170
timestamp 1677677812
transform 1 0 1972 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3575
timestamp 1677677812
transform 1 0 1972 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3122
timestamp 1677677812
transform 1 0 2012 0 1 3045
box -3 -3 3 3
use M2_M1  M2_M1_3576
timestamp 1677677812
transform 1 0 2012 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3683
timestamp 1677677812
transform 1 0 1988 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3684
timestamp 1677677812
transform 1 0 2004 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3243
timestamp 1677677812
transform 1 0 2012 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3685
timestamp 1677677812
transform 1 0 2036 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3274
timestamp 1677677812
transform 1 0 2036 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3123
timestamp 1677677812
transform 1 0 2052 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3124
timestamp 1677677812
transform 1 0 2092 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3125
timestamp 1677677812
transform 1 0 2180 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3171
timestamp 1677677812
transform 1 0 2084 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3172
timestamp 1677677812
transform 1 0 2156 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3173
timestamp 1677677812
transform 1 0 2196 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3577
timestamp 1677677812
transform 1 0 2068 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3578
timestamp 1677677812
transform 1 0 2084 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3579
timestamp 1677677812
transform 1 0 2100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3580
timestamp 1677677812
transform 1 0 2156 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3581
timestamp 1677677812
transform 1 0 2196 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3686
timestamp 1677677812
transform 1 0 2060 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3687
timestamp 1677677812
transform 1 0 2076 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3688
timestamp 1677677812
transform 1 0 2092 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3689
timestamp 1677677812
transform 1 0 2180 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3690
timestamp 1677677812
transform 1 0 2196 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3244
timestamp 1677677812
transform 1 0 2068 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3245
timestamp 1677677812
transform 1 0 2084 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3275
timestamp 1677677812
transform 1 0 2076 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3126
timestamp 1677677812
transform 1 0 2236 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3137
timestamp 1677677812
transform 1 0 2228 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3582
timestamp 1677677812
transform 1 0 2220 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3246
timestamp 1677677812
transform 1 0 2228 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3095
timestamp 1677677812
transform 1 0 2292 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3174
timestamp 1677677812
transform 1 0 2284 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3583
timestamp 1677677812
transform 1 0 2268 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3584
timestamp 1677677812
transform 1 0 2276 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3691
timestamp 1677677812
transform 1 0 2260 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3247
timestamp 1677677812
transform 1 0 2260 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3692
timestamp 1677677812
transform 1 0 2284 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3693
timestamp 1677677812
transform 1 0 2292 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3096
timestamp 1677677812
transform 1 0 2308 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3138
timestamp 1677677812
transform 1 0 2332 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3175
timestamp 1677677812
transform 1 0 2308 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3585
timestamp 1677677812
transform 1 0 2316 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3586
timestamp 1677677812
transform 1 0 2332 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3694
timestamp 1677677812
transform 1 0 2332 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3097
timestamp 1677677812
transform 1 0 2348 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3139
timestamp 1677677812
transform 1 0 2372 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3587
timestamp 1677677812
transform 1 0 2364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3588
timestamp 1677677812
transform 1 0 2372 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3589
timestamp 1677677812
transform 1 0 2388 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3201
timestamp 1677677812
transform 1 0 2396 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3590
timestamp 1677677812
transform 1 0 2404 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3695
timestamp 1677677812
transform 1 0 2356 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3221
timestamp 1677677812
transform 1 0 2364 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3696
timestamp 1677677812
transform 1 0 2372 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3222
timestamp 1677677812
transform 1 0 2388 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3591
timestamp 1677677812
transform 1 0 2420 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3697
timestamp 1677677812
transform 1 0 2420 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3098
timestamp 1677677812
transform 1 0 2444 0 1 3065
box -3 -3 3 3
use M3_M2  M3_M2_3106
timestamp 1677677812
transform 1 0 2524 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3592
timestamp 1677677812
transform 1 0 2492 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3593
timestamp 1677677812
transform 1 0 2500 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3594
timestamp 1677677812
transform 1 0 2516 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3595
timestamp 1677677812
transform 1 0 2540 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3140
timestamp 1677677812
transform 1 0 2548 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3698
timestamp 1677677812
transform 1 0 2508 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3699
timestamp 1677677812
transform 1 0 2524 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3700
timestamp 1677677812
transform 1 0 2532 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3223
timestamp 1677677812
transform 1 0 2540 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3107
timestamp 1677677812
transform 1 0 2612 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3176
timestamp 1677677812
transform 1 0 2604 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3177
timestamp 1677677812
transform 1 0 2644 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3596
timestamp 1677677812
transform 1 0 2604 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3597
timestamp 1677677812
transform 1 0 2612 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3598
timestamp 1677677812
transform 1 0 2644 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3202
timestamp 1677677812
transform 1 0 2692 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3224
timestamp 1677677812
transform 1 0 2620 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3701
timestamp 1677677812
transform 1 0 2692 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3141
timestamp 1677677812
transform 1 0 2708 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3702
timestamp 1677677812
transform 1 0 2708 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3599
timestamp 1677677812
transform 1 0 2796 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3225
timestamp 1677677812
transform 1 0 2796 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3525
timestamp 1677677812
transform 1 0 2828 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3178
timestamp 1677677812
transform 1 0 2836 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3203
timestamp 1677677812
transform 1 0 2828 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3703
timestamp 1677677812
transform 1 0 2836 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3750
timestamp 1677677812
transform 1 0 2828 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3179
timestamp 1677677812
transform 1 0 2860 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3600
timestamp 1677677812
transform 1 0 2860 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3226
timestamp 1677677812
transform 1 0 2852 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3227
timestamp 1677677812
transform 1 0 2868 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3751
timestamp 1677677812
transform 1 0 2852 0 1 2995
box -2 -2 2 2
use M2_M1  M2_M1_3752
timestamp 1677677812
transform 1 0 2860 0 1 2995
box -2 -2 2 2
use M3_M2  M3_M2_3276
timestamp 1677677812
transform 1 0 2860 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3180
timestamp 1677677812
transform 1 0 2892 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3181
timestamp 1677677812
transform 1 0 2908 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3099
timestamp 1677677812
transform 1 0 2932 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3526
timestamp 1677677812
transform 1 0 2932 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3601
timestamp 1677677812
transform 1 0 2916 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3704
timestamp 1677677812
transform 1 0 2908 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3204
timestamp 1677677812
transform 1 0 2924 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3705
timestamp 1677677812
transform 1 0 2924 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3100
timestamp 1677677812
transform 1 0 2972 0 1 3065
box -3 -3 3 3
use M2_M1  M2_M1_3527
timestamp 1677677812
transform 1 0 2996 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3602
timestamp 1677677812
transform 1 0 3004 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3205
timestamp 1677677812
transform 1 0 3012 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3706
timestamp 1677677812
transform 1 0 3012 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3182
timestamp 1677677812
transform 1 0 3028 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3603
timestamp 1677677812
transform 1 0 3028 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3604
timestamp 1677677812
transform 1 0 3044 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3707
timestamp 1677677812
transform 1 0 3036 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3248
timestamp 1677677812
transform 1 0 3036 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3142
timestamp 1677677812
transform 1 0 3100 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3605
timestamp 1677677812
transform 1 0 3100 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3606
timestamp 1677677812
transform 1 0 3132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3708
timestamp 1677677812
transform 1 0 3092 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3709
timestamp 1677677812
transform 1 0 3180 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3249
timestamp 1677677812
transform 1 0 3132 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3250
timestamp 1677677812
transform 1 0 3180 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3143
timestamp 1677677812
transform 1 0 3244 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3183
timestamp 1677677812
transform 1 0 3220 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3607
timestamp 1677677812
transform 1 0 3220 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3206
timestamp 1677677812
transform 1 0 3228 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3608
timestamp 1677677812
transform 1 0 3236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3710
timestamp 1677677812
transform 1 0 3212 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3711
timestamp 1677677812
transform 1 0 3228 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3228
timestamp 1677677812
transform 1 0 3236 0 1 3005
box -3 -3 3 3
use M2_M1  M2_M1_3712
timestamp 1677677812
transform 1 0 3244 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3251
timestamp 1677677812
transform 1 0 3228 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3609
timestamp 1677677812
transform 1 0 3308 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3713
timestamp 1677677812
transform 1 0 3284 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3229
timestamp 1677677812
transform 1 0 3308 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3252
timestamp 1677677812
transform 1 0 3284 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3207
timestamp 1677677812
transform 1 0 3388 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3610
timestamp 1677677812
transform 1 0 3396 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3528
timestamp 1677677812
transform 1 0 3412 0 1 3025
box -2 -2 2 2
use M2_M1  M2_M1_3522
timestamp 1677677812
transform 1 0 3436 0 1 3035
box -2 -2 2 2
use M2_M1  M2_M1_3611
timestamp 1677677812
transform 1 0 3444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3529
timestamp 1677677812
transform 1 0 3468 0 1 3025
box -2 -2 2 2
use M3_M2  M3_M2_3108
timestamp 1677677812
transform 1 0 3492 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3109
timestamp 1677677812
transform 1 0 3524 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3144
timestamp 1677677812
transform 1 0 3548 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3612
timestamp 1677677812
transform 1 0 3532 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3714
timestamp 1677677812
transform 1 0 3484 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3253
timestamp 1677677812
transform 1 0 3532 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3208
timestamp 1677677812
transform 1 0 3572 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3613
timestamp 1677677812
transform 1 0 3580 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3614
timestamp 1677677812
transform 1 0 3588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3615
timestamp 1677677812
transform 1 0 3604 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3715
timestamp 1677677812
transform 1 0 3572 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3716
timestamp 1677677812
transform 1 0 3596 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3717
timestamp 1677677812
transform 1 0 3612 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3254
timestamp 1677677812
transform 1 0 3596 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3277
timestamp 1677677812
transform 1 0 3588 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3718
timestamp 1677677812
transform 1 0 3636 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3184
timestamp 1677677812
transform 1 0 3660 0 1 3025
box -3 -3 3 3
use M3_M2  M3_M2_3145
timestamp 1677677812
transform 1 0 3676 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3616
timestamp 1677677812
transform 1 0 3676 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3209
timestamp 1677677812
transform 1 0 3700 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3617
timestamp 1677677812
transform 1 0 3708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3719
timestamp 1677677812
transform 1 0 3684 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3720
timestamp 1677677812
transform 1 0 3700 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3255
timestamp 1677677812
transform 1 0 3684 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3210
timestamp 1677677812
transform 1 0 3740 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3110
timestamp 1677677812
transform 1 0 3756 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3111
timestamp 1677677812
transform 1 0 3788 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3112
timestamp 1677677812
transform 1 0 3836 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3618
timestamp 1677677812
transform 1 0 3780 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3721
timestamp 1677677812
transform 1 0 3756 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3256
timestamp 1677677812
transform 1 0 3780 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3278
timestamp 1677677812
transform 1 0 3836 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3127
timestamp 1677677812
transform 1 0 3868 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3146
timestamp 1677677812
transform 1 0 3860 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3619
timestamp 1677677812
transform 1 0 3860 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3620
timestamp 1677677812
transform 1 0 3868 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3113
timestamp 1677677812
transform 1 0 3884 0 1 3055
box -3 -3 3 3
use M2_M1  M2_M1_3722
timestamp 1677677812
transform 1 0 3884 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3128
timestamp 1677677812
transform 1 0 3924 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3114
timestamp 1677677812
transform 1 0 3948 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3147
timestamp 1677677812
transform 1 0 3940 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3621
timestamp 1677677812
transform 1 0 3988 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3622
timestamp 1677677812
transform 1 0 4036 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3723
timestamp 1677677812
transform 1 0 3940 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3230
timestamp 1677677812
transform 1 0 3988 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3231
timestamp 1677677812
transform 1 0 4020 0 1 3005
box -3 -3 3 3
use M3_M2  M3_M2_3279
timestamp 1677677812
transform 1 0 3940 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3724
timestamp 1677677812
transform 1 0 4052 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3725
timestamp 1677677812
transform 1 0 4076 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3129
timestamp 1677677812
transform 1 0 4092 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3115
timestamp 1677677812
transform 1 0 4108 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3148
timestamp 1677677812
transform 1 0 4116 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3726
timestamp 1677677812
transform 1 0 4108 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3623
timestamp 1677677812
transform 1 0 4132 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3624
timestamp 1677677812
transform 1 0 4148 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3727
timestamp 1677677812
transform 1 0 4140 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3728
timestamp 1677677812
transform 1 0 4156 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3729
timestamp 1677677812
transform 1 0 4164 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3257
timestamp 1677677812
transform 1 0 4132 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3280
timestamp 1677677812
transform 1 0 4156 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3116
timestamp 1677677812
transform 1 0 4180 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3185
timestamp 1677677812
transform 1 0 4180 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3625
timestamp 1677677812
transform 1 0 4180 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3211
timestamp 1677677812
transform 1 0 4188 0 1 3015
box -3 -3 3 3
use M2_M1  M2_M1_3626
timestamp 1677677812
transform 1 0 4196 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3186
timestamp 1677677812
transform 1 0 4236 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3627
timestamp 1677677812
transform 1 0 4236 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3730
timestamp 1677677812
transform 1 0 4228 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3628
timestamp 1677677812
transform 1 0 4260 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3731
timestamp 1677677812
transform 1 0 4292 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3117
timestamp 1677677812
transform 1 0 4356 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3130
timestamp 1677677812
transform 1 0 4340 0 1 3045
box -3 -3 3 3
use M3_M2  M3_M2_3149
timestamp 1677677812
transform 1 0 4348 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3187
timestamp 1677677812
transform 1 0 4324 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3629
timestamp 1677677812
transform 1 0 4324 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3630
timestamp 1677677812
transform 1 0 4340 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3631
timestamp 1677677812
transform 1 0 4356 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3632
timestamp 1677677812
transform 1 0 4364 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3732
timestamp 1677677812
transform 1 0 4324 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3258
timestamp 1677677812
transform 1 0 4364 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3212
timestamp 1677677812
transform 1 0 4380 0 1 3015
box -3 -3 3 3
use M3_M2  M3_M2_3150
timestamp 1677677812
transform 1 0 4428 0 1 3035
box -3 -3 3 3
use M3_M2  M3_M2_3188
timestamp 1677677812
transform 1 0 4412 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3633
timestamp 1677677812
transform 1 0 4412 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3634
timestamp 1677677812
transform 1 0 4428 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3635
timestamp 1677677812
transform 1 0 4444 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3733
timestamp 1677677812
transform 1 0 4396 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3734
timestamp 1677677812
transform 1 0 4404 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3735
timestamp 1677677812
transform 1 0 4420 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3736
timestamp 1677677812
transform 1 0 4436 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3259
timestamp 1677677812
transform 1 0 4396 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3260
timestamp 1677677812
transform 1 0 4428 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3281
timestamp 1677677812
transform 1 0 4436 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3636
timestamp 1677677812
transform 1 0 4476 0 1 3015
box -2 -2 2 2
use M3_M2  M3_M2_3151
timestamp 1677677812
transform 1 0 4492 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3737
timestamp 1677677812
transform 1 0 4484 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3738
timestamp 1677677812
transform 1 0 4500 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3118
timestamp 1677677812
transform 1 0 4532 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3152
timestamp 1677677812
transform 1 0 4540 0 1 3035
box -3 -3 3 3
use M2_M1  M2_M1_3637
timestamp 1677677812
transform 1 0 4540 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3739
timestamp 1677677812
transform 1 0 4532 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3740
timestamp 1677677812
transform 1 0 4548 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3741
timestamp 1677677812
transform 1 0 4556 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3119
timestamp 1677677812
transform 1 0 4620 0 1 3055
box -3 -3 3 3
use M3_M2  M3_M2_3189
timestamp 1677677812
transform 1 0 4628 0 1 3025
box -3 -3 3 3
use M2_M1  M2_M1_3638
timestamp 1677677812
transform 1 0 4588 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3639
timestamp 1677677812
transform 1 0 4604 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3640
timestamp 1677677812
transform 1 0 4620 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3641
timestamp 1677677812
transform 1 0 4628 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3742
timestamp 1677677812
transform 1 0 4596 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3261
timestamp 1677677812
transform 1 0 4596 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3262
timestamp 1677677812
transform 1 0 4628 0 1 2995
box -3 -3 3 3
use M2_M1  M2_M1_3642
timestamp 1677677812
transform 1 0 4652 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3643
timestamp 1677677812
transform 1 0 4692 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3644
timestamp 1677677812
transform 1 0 4708 0 1 3015
box -2 -2 2 2
use M2_M1  M2_M1_3743
timestamp 1677677812
transform 1 0 4660 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3744
timestamp 1677677812
transform 1 0 4668 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3745
timestamp 1677677812
transform 1 0 4684 0 1 3005
box -2 -2 2 2
use M2_M1  M2_M1_3746
timestamp 1677677812
transform 1 0 4700 0 1 3005
box -2 -2 2 2
use M3_M2  M3_M2_3263
timestamp 1677677812
transform 1 0 4660 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3264
timestamp 1677677812
transform 1 0 4692 0 1 2995
box -3 -3 3 3
use M3_M2  M3_M2_3282
timestamp 1677677812
transform 1 0 4676 0 1 2985
box -3 -3 3 3
use M3_M2  M3_M2_3283
timestamp 1677677812
transform 1 0 4700 0 1 2985
box -3 -3 3 3
use M2_M1  M2_M1_3753
timestamp 1677677812
transform 1 0 4772 0 1 2995
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_34
timestamp 1677677812
transform 1 0 48 0 1 2970
box -10 -3 10 3
use FILL  FILL_3796
timestamp 1677677812
transform 1 0 72 0 1 2970
box -8 -3 16 105
use FILL  FILL_3797
timestamp 1677677812
transform 1 0 80 0 1 2970
box -8 -3 16 105
use FILL  FILL_3798
timestamp 1677677812
transform 1 0 88 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_269
timestamp 1677677812
transform 1 0 96 0 1 2970
box -9 -3 26 105
use AOI22X1  AOI22X1_163
timestamp 1677677812
transform -1 0 152 0 1 2970
box -8 -3 46 105
use FILL  FILL_3799
timestamp 1677677812
transform 1 0 152 0 1 2970
box -8 -3 16 105
use FILL  FILL_3800
timestamp 1677677812
transform 1 0 160 0 1 2970
box -8 -3 16 105
use FILL  FILL_3801
timestamp 1677677812
transform 1 0 168 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3284
timestamp 1677677812
transform 1 0 196 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_155
timestamp 1677677812
transform -1 0 216 0 1 2970
box -8 -3 46 105
use FILL  FILL_3802
timestamp 1677677812
transform 1 0 216 0 1 2970
box -8 -3 16 105
use FILL  FILL_3803
timestamp 1677677812
transform 1 0 224 0 1 2970
box -8 -3 16 105
use FILL  FILL_3804
timestamp 1677677812
transform 1 0 232 0 1 2970
box -8 -3 16 105
use FILL  FILL_3805
timestamp 1677677812
transform 1 0 240 0 1 2970
box -8 -3 16 105
use FILL  FILL_3806
timestamp 1677677812
transform 1 0 248 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_156
timestamp 1677677812
transform -1 0 296 0 1 2970
box -8 -3 46 105
use FILL  FILL_3807
timestamp 1677677812
transform 1 0 296 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_237
timestamp 1677677812
transform 1 0 304 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_270
timestamp 1677677812
transform -1 0 416 0 1 2970
box -9 -3 26 105
use FILL  FILL_3808
timestamp 1677677812
transform 1 0 416 0 1 2970
box -8 -3 16 105
use FILL  FILL_3809
timestamp 1677677812
transform 1 0 424 0 1 2970
box -8 -3 16 105
use FILL  FILL_3812
timestamp 1677677812
transform 1 0 432 0 1 2970
box -8 -3 16 105
use FILL  FILL_3814
timestamp 1677677812
transform 1 0 440 0 1 2970
box -8 -3 16 105
use FILL  FILL_3816
timestamp 1677677812
transform 1 0 448 0 1 2970
box -8 -3 16 105
use FILL  FILL_3818
timestamp 1677677812
transform 1 0 456 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_241
timestamp 1677677812
transform 1 0 464 0 1 2970
box -8 -3 104 105
use FILL  FILL_3820
timestamp 1677677812
transform 1 0 560 0 1 2970
box -8 -3 16 105
use FILL  FILL_3821
timestamp 1677677812
transform 1 0 568 0 1 2970
box -8 -3 16 105
use FILL  FILL_3822
timestamp 1677677812
transform 1 0 576 0 1 2970
box -8 -3 16 105
use FILL  FILL_3823
timestamp 1677677812
transform 1 0 584 0 1 2970
box -8 -3 16 105
use FILL  FILL_3830
timestamp 1677677812
transform 1 0 592 0 1 2970
box -8 -3 16 105
use FILL  FILL_3832
timestamp 1677677812
transform 1 0 600 0 1 2970
box -8 -3 16 105
use FILL  FILL_3834
timestamp 1677677812
transform 1 0 608 0 1 2970
box -8 -3 16 105
use FILL  FILL_3836
timestamp 1677677812
transform 1 0 616 0 1 2970
box -8 -3 16 105
use FILL  FILL_3838
timestamp 1677677812
transform 1 0 624 0 1 2970
box -8 -3 16 105
use FILL  FILL_3840
timestamp 1677677812
transform 1 0 632 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_157
timestamp 1677677812
transform 1 0 640 0 1 2970
box -8 -3 46 105
use FILL  FILL_3841
timestamp 1677677812
transform 1 0 680 0 1 2970
box -8 -3 16 105
use FILL  FILL_3844
timestamp 1677677812
transform 1 0 688 0 1 2970
box -8 -3 16 105
use FILL  FILL_3846
timestamp 1677677812
transform 1 0 696 0 1 2970
box -8 -3 16 105
use FILL  FILL_3848
timestamp 1677677812
transform 1 0 704 0 1 2970
box -8 -3 16 105
use FILL  FILL_3850
timestamp 1677677812
transform 1 0 712 0 1 2970
box -8 -3 16 105
use FILL  FILL_3851
timestamp 1677677812
transform 1 0 720 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_272
timestamp 1677677812
transform -1 0 744 0 1 2970
box -9 -3 26 105
use FILL  FILL_3852
timestamp 1677677812
transform 1 0 744 0 1 2970
box -8 -3 16 105
use FILL  FILL_3853
timestamp 1677677812
transform 1 0 752 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3285
timestamp 1677677812
transform 1 0 772 0 1 2975
box -3 -3 3 3
use FILL  FILL_3854
timestamp 1677677812
transform 1 0 760 0 1 2970
box -8 -3 16 105
use FILL  FILL_3855
timestamp 1677677812
transform 1 0 768 0 1 2970
box -8 -3 16 105
use FILL  FILL_3856
timestamp 1677677812
transform 1 0 776 0 1 2970
box -8 -3 16 105
use FILL  FILL_3857
timestamp 1677677812
transform 1 0 784 0 1 2970
box -8 -3 16 105
use FILL  FILL_3858
timestamp 1677677812
transform 1 0 792 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_39
timestamp 1677677812
transform 1 0 800 0 1 2970
box -8 -3 32 105
use FILL  FILL_3859
timestamp 1677677812
transform 1 0 824 0 1 2970
box -8 -3 16 105
use FILL  FILL_3863
timestamp 1677677812
transform 1 0 832 0 1 2970
box -8 -3 16 105
use FILL  FILL_3865
timestamp 1677677812
transform 1 0 840 0 1 2970
box -8 -3 16 105
use FILL  FILL_3866
timestamp 1677677812
transform 1 0 848 0 1 2970
box -8 -3 16 105
use FILL  FILL_3867
timestamp 1677677812
transform 1 0 856 0 1 2970
box -8 -3 16 105
use FILL  FILL_3869
timestamp 1677677812
transform 1 0 864 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_83
timestamp 1677677812
transform 1 0 872 0 1 2970
box -8 -3 34 105
use FILL  FILL_3871
timestamp 1677677812
transform 1 0 904 0 1 2970
box -8 -3 16 105
use FILL  FILL_3877
timestamp 1677677812
transform 1 0 912 0 1 2970
box -8 -3 16 105
use FILL  FILL_3879
timestamp 1677677812
transform 1 0 920 0 1 2970
box -8 -3 16 105
use FILL  FILL_3881
timestamp 1677677812
transform 1 0 928 0 1 2970
box -8 -3 16 105
use FILL  FILL_3882
timestamp 1677677812
transform 1 0 936 0 1 2970
box -8 -3 16 105
use FILL  FILL_3883
timestamp 1677677812
transform 1 0 944 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_40
timestamp 1677677812
transform 1 0 952 0 1 2970
box -8 -3 32 105
use FILL  FILL_3884
timestamp 1677677812
transform 1 0 976 0 1 2970
box -8 -3 16 105
use FILL  FILL_3889
timestamp 1677677812
transform 1 0 984 0 1 2970
box -8 -3 16 105
use FILL  FILL_3891
timestamp 1677677812
transform 1 0 992 0 1 2970
box -8 -3 16 105
use FILL  FILL_3893
timestamp 1677677812
transform 1 0 1000 0 1 2970
box -8 -3 16 105
use FILL  FILL_3895
timestamp 1677677812
transform 1 0 1008 0 1 2970
box -8 -3 16 105
use FILL  FILL_3897
timestamp 1677677812
transform 1 0 1016 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_274
timestamp 1677677812
transform 1 0 1024 0 1 2970
box -9 -3 26 105
use FILL  FILL_3898
timestamp 1677677812
transform 1 0 1040 0 1 2970
box -8 -3 16 105
use FILL  FILL_3899
timestamp 1677677812
transform 1 0 1048 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_243
timestamp 1677677812
transform -1 0 1152 0 1 2970
box -8 -3 104 105
use FILL  FILL_3900
timestamp 1677677812
transform 1 0 1152 0 1 2970
box -8 -3 16 105
use FILL  FILL_3901
timestamp 1677677812
transform 1 0 1160 0 1 2970
box -8 -3 16 105
use FILL  FILL_3902
timestamp 1677677812
transform 1 0 1168 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_42
timestamp 1677677812
transform 1 0 1176 0 1 2970
box -8 -3 32 105
use FILL  FILL_3903
timestamp 1677677812
transform 1 0 1200 0 1 2970
box -8 -3 16 105
use FILL  FILL_3918
timestamp 1677677812
transform 1 0 1208 0 1 2970
box -8 -3 16 105
use FILL  FILL_3920
timestamp 1677677812
transform 1 0 1216 0 1 2970
box -8 -3 16 105
use FILL  FILL_3922
timestamp 1677677812
transform 1 0 1224 0 1 2970
box -8 -3 16 105
use FILL  FILL_3924
timestamp 1677677812
transform 1 0 1232 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_169
timestamp 1677677812
transform 1 0 1240 0 1 2970
box -8 -3 46 105
use FILL  FILL_3926
timestamp 1677677812
transform 1 0 1280 0 1 2970
box -8 -3 16 105
use FILL  FILL_3927
timestamp 1677677812
transform 1 0 1288 0 1 2970
box -8 -3 16 105
use FILL  FILL_3928
timestamp 1677677812
transform 1 0 1296 0 1 2970
box -8 -3 16 105
use FILL  FILL_3933
timestamp 1677677812
transform 1 0 1304 0 1 2970
box -8 -3 16 105
use FILL  FILL_3935
timestamp 1677677812
transform 1 0 1312 0 1 2970
box -8 -3 16 105
use FILL  FILL_3937
timestamp 1677677812
transform 1 0 1320 0 1 2970
box -8 -3 16 105
use FILL  FILL_3939
timestamp 1677677812
transform 1 0 1328 0 1 2970
box -8 -3 16 105
use FILL  FILL_3941
timestamp 1677677812
transform 1 0 1336 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_85
timestamp 1677677812
transform -1 0 1376 0 1 2970
box -8 -3 34 105
use FILL  FILL_3943
timestamp 1677677812
transform 1 0 1376 0 1 2970
box -8 -3 16 105
use FILL  FILL_3945
timestamp 1677677812
transform 1 0 1384 0 1 2970
box -8 -3 16 105
use FILL  FILL_3947
timestamp 1677677812
transform 1 0 1392 0 1 2970
box -8 -3 16 105
use FILL  FILL_3949
timestamp 1677677812
transform 1 0 1400 0 1 2970
box -8 -3 16 105
use FILL  FILL_3951
timestamp 1677677812
transform 1 0 1408 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_244
timestamp 1677677812
transform -1 0 1512 0 1 2970
box -8 -3 104 105
use FILL  FILL_3952
timestamp 1677677812
transform 1 0 1512 0 1 2970
box -8 -3 16 105
use FILL  FILL_3953
timestamp 1677677812
transform 1 0 1520 0 1 2970
box -8 -3 16 105
use FILL  FILL_3954
timestamp 1677677812
transform 1 0 1528 0 1 2970
box -8 -3 16 105
use FILL  FILL_3955
timestamp 1677677812
transform 1 0 1536 0 1 2970
box -8 -3 16 105
use FILL  FILL_3956
timestamp 1677677812
transform 1 0 1544 0 1 2970
box -8 -3 16 105
use FILL  FILL_3957
timestamp 1677677812
transform 1 0 1552 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_159
timestamp 1677677812
transform 1 0 1560 0 1 2970
box -8 -3 46 105
use FILL  FILL_3958
timestamp 1677677812
transform 1 0 1600 0 1 2970
box -8 -3 16 105
use FILL  FILL_3968
timestamp 1677677812
transform 1 0 1608 0 1 2970
box -8 -3 16 105
use FILL  FILL_3970
timestamp 1677677812
transform 1 0 1616 0 1 2970
box -8 -3 16 105
use FILL  FILL_3971
timestamp 1677677812
transform 1 0 1624 0 1 2970
box -8 -3 16 105
use FILL  FILL_3972
timestamp 1677677812
transform 1 0 1632 0 1 2970
box -8 -3 16 105
use FILL  FILL_3974
timestamp 1677677812
transform 1 0 1640 0 1 2970
box -8 -3 16 105
use FILL  FILL_3976
timestamp 1677677812
transform 1 0 1648 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3286
timestamp 1677677812
transform 1 0 1684 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_160
timestamp 1677677812
transform -1 0 1696 0 1 2970
box -8 -3 46 105
use FILL  FILL_3977
timestamp 1677677812
transform 1 0 1696 0 1 2970
box -8 -3 16 105
use FILL  FILL_3983
timestamp 1677677812
transform 1 0 1704 0 1 2970
box -8 -3 16 105
use FILL  FILL_3984
timestamp 1677677812
transform 1 0 1712 0 1 2970
box -8 -3 16 105
use FILL  FILL_3985
timestamp 1677677812
transform 1 0 1720 0 1 2970
box -8 -3 16 105
use FILL  FILL_3986
timestamp 1677677812
transform 1 0 1728 0 1 2970
box -8 -3 16 105
use FILL  FILL_3987
timestamp 1677677812
transform 1 0 1736 0 1 2970
box -8 -3 16 105
use BUFX2  BUFX2_28
timestamp 1677677812
transform 1 0 1744 0 1 2970
box -5 -3 28 105
use INVX2  INVX2_277
timestamp 1677677812
transform 1 0 1768 0 1 2970
box -9 -3 26 105
use FILL  FILL_3990
timestamp 1677677812
transform 1 0 1784 0 1 2970
box -8 -3 16 105
use FILL  FILL_3991
timestamp 1677677812
transform 1 0 1792 0 1 2970
box -8 -3 16 105
use FILL  FILL_3992
timestamp 1677677812
transform 1 0 1800 0 1 2970
box -8 -3 16 105
use FILL  FILL_3993
timestamp 1677677812
transform 1 0 1808 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_170
timestamp 1677677812
transform 1 0 1816 0 1 2970
box -8 -3 46 105
use FILL  FILL_3994
timestamp 1677677812
transform 1 0 1856 0 1 2970
box -8 -3 16 105
use FILL  FILL_3998
timestamp 1677677812
transform 1 0 1864 0 1 2970
box -8 -3 16 105
use FILL  FILL_4000
timestamp 1677677812
transform 1 0 1872 0 1 2970
box -8 -3 16 105
use FILL  FILL_4002
timestamp 1677677812
transform 1 0 1880 0 1 2970
box -8 -3 16 105
use FILL  FILL_4004
timestamp 1677677812
transform 1 0 1888 0 1 2970
box -8 -3 16 105
use FILL  FILL_4005
timestamp 1677677812
transform 1 0 1896 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3287
timestamp 1677677812
transform 1 0 1916 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_161
timestamp 1677677812
transform 1 0 1904 0 1 2970
box -8 -3 46 105
use FILL  FILL_4006
timestamp 1677677812
transform 1 0 1944 0 1 2970
box -8 -3 16 105
use FILL  FILL_4010
timestamp 1677677812
transform 1 0 1952 0 1 2970
box -8 -3 16 105
use FILL  FILL_4012
timestamp 1677677812
transform 1 0 1960 0 1 2970
box -8 -3 16 105
use FILL  FILL_4013
timestamp 1677677812
transform 1 0 1968 0 1 2970
box -8 -3 16 105
use FILL  FILL_4014
timestamp 1677677812
transform 1 0 1976 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3288
timestamp 1677677812
transform 1 0 2020 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_162
timestamp 1677677812
transform 1 0 1984 0 1 2970
box -8 -3 46 105
use FILL  FILL_4015
timestamp 1677677812
transform 1 0 2024 0 1 2970
box -8 -3 16 105
use FILL  FILL_4016
timestamp 1677677812
transform 1 0 2032 0 1 2970
box -8 -3 16 105
use FILL  FILL_4017
timestamp 1677677812
transform 1 0 2040 0 1 2970
box -8 -3 16 105
use FILL  FILL_4018
timestamp 1677677812
transform 1 0 2048 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3289
timestamp 1677677812
transform 1 0 2076 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_163
timestamp 1677677812
transform -1 0 2096 0 1 2970
box -8 -3 46 105
use M3_M2  M3_M2_3290
timestamp 1677677812
transform 1 0 2124 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3291
timestamp 1677677812
transform 1 0 2140 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3292
timestamp 1677677812
transform 1 0 2172 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3293
timestamp 1677677812
transform 1 0 2196 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_247
timestamp 1677677812
transform -1 0 2192 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_278
timestamp 1677677812
transform 1 0 2192 0 1 2970
box -9 -3 26 105
use FILL  FILL_4019
timestamp 1677677812
transform 1 0 2208 0 1 2970
box -8 -3 16 105
use BUFX2  BUFX2_29
timestamp 1677677812
transform 1 0 2216 0 1 2970
box -5 -3 28 105
use FILL  FILL_4035
timestamp 1677677812
transform 1 0 2240 0 1 2970
box -8 -3 16 105
use FILL  FILL_4036
timestamp 1677677812
transform 1 0 2248 0 1 2970
box -8 -3 16 105
use FILL  FILL_4037
timestamp 1677677812
transform 1 0 2256 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_280
timestamp 1677677812
transform -1 0 2280 0 1 2970
box -9 -3 26 105
use FILL  FILL_4038
timestamp 1677677812
transform 1 0 2280 0 1 2970
box -8 -3 16 105
use FILL  FILL_4039
timestamp 1677677812
transform 1 0 2288 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3294
timestamp 1677677812
transform 1 0 2332 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_175
timestamp 1677677812
transform -1 0 2336 0 1 2970
box -8 -3 46 105
use FILL  FILL_4040
timestamp 1677677812
transform 1 0 2336 0 1 2970
box -8 -3 16 105
use FILL  FILL_4045
timestamp 1677677812
transform 1 0 2344 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3295
timestamp 1677677812
transform 1 0 2372 0 1 2975
box -3 -3 3 3
use INVX2  INVX2_281
timestamp 1677677812
transform 1 0 2352 0 1 2970
box -9 -3 26 105
use M3_M2  M3_M2_3296
timestamp 1677677812
transform 1 0 2396 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_176
timestamp 1677677812
transform 1 0 2368 0 1 2970
box -8 -3 46 105
use FILL  FILL_4047
timestamp 1677677812
transform 1 0 2408 0 1 2970
box -8 -3 16 105
use FILL  FILL_4056
timestamp 1677677812
transform 1 0 2416 0 1 2970
box -8 -3 16 105
use FILL  FILL_4058
timestamp 1677677812
transform 1 0 2424 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_282
timestamp 1677677812
transform 1 0 2432 0 1 2970
box -9 -3 26 105
use FILL  FILL_4060
timestamp 1677677812
transform 1 0 2448 0 1 2970
box -8 -3 16 105
use FILL  FILL_4061
timestamp 1677677812
transform 1 0 2456 0 1 2970
box -8 -3 16 105
use FILL  FILL_4062
timestamp 1677677812
transform 1 0 2464 0 1 2970
box -8 -3 16 105
use FILL  FILL_4063
timestamp 1677677812
transform 1 0 2472 0 1 2970
box -8 -3 16 105
use FILL  FILL_4064
timestamp 1677677812
transform 1 0 2480 0 1 2970
box -8 -3 16 105
use FILL  FILL_4065
timestamp 1677677812
transform 1 0 2488 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_177
timestamp 1677677812
transform 1 0 2496 0 1 2970
box -8 -3 46 105
use FILL  FILL_4066
timestamp 1677677812
transform 1 0 2536 0 1 2970
box -8 -3 16 105
use FILL  FILL_4067
timestamp 1677677812
transform 1 0 2544 0 1 2970
box -8 -3 16 105
use FILL  FILL_4068
timestamp 1677677812
transform 1 0 2552 0 1 2970
box -8 -3 16 105
use FILL  FILL_4073
timestamp 1677677812
transform 1 0 2560 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_283
timestamp 1677677812
transform 1 0 2568 0 1 2970
box -9 -3 26 105
use FILL  FILL_4075
timestamp 1677677812
transform 1 0 2584 0 1 2970
box -8 -3 16 105
use FILL  FILL_4076
timestamp 1677677812
transform 1 0 2592 0 1 2970
box -8 -3 16 105
use FILL  FILL_4077
timestamp 1677677812
transform 1 0 2600 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_250
timestamp 1677677812
transform -1 0 2704 0 1 2970
box -8 -3 104 105
use FILL  FILL_4078
timestamp 1677677812
transform 1 0 2704 0 1 2970
box -8 -3 16 105
use FILL  FILL_4079
timestamp 1677677812
transform 1 0 2712 0 1 2970
box -8 -3 16 105
use FILL  FILL_4080
timestamp 1677677812
transform 1 0 2720 0 1 2970
box -8 -3 16 105
use FILL  FILL_4081
timestamp 1677677812
transform 1 0 2728 0 1 2970
box -8 -3 16 105
use FILL  FILL_4082
timestamp 1677677812
transform 1 0 2736 0 1 2970
box -8 -3 16 105
use FILL  FILL_4083
timestamp 1677677812
transform 1 0 2744 0 1 2970
box -8 -3 16 105
use FILL  FILL_4084
timestamp 1677677812
transform 1 0 2752 0 1 2970
box -8 -3 16 105
use FILL  FILL_4085
timestamp 1677677812
transform 1 0 2760 0 1 2970
box -8 -3 16 105
use FILL  FILL_4086
timestamp 1677677812
transform 1 0 2768 0 1 2970
box -8 -3 16 105
use FILL  FILL_4094
timestamp 1677677812
transform 1 0 2776 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_88
timestamp 1677677812
transform 1 0 2784 0 1 2970
box -8 -3 34 105
use M3_M2  M3_M2_3297
timestamp 1677677812
transform 1 0 2828 0 1 2975
box -3 -3 3 3
use FILL  FILL_4096
timestamp 1677677812
transform 1 0 2816 0 1 2970
box -8 -3 16 105
use FILL  FILL_4102
timestamp 1677677812
transform 1 0 2824 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_43
timestamp 1677677812
transform 1 0 2832 0 1 2970
box -8 -3 32 105
use FILL  FILL_4103
timestamp 1677677812
transform 1 0 2856 0 1 2970
box -8 -3 16 105
use FILL  FILL_4106
timestamp 1677677812
transform 1 0 2864 0 1 2970
box -8 -3 16 105
use FILL  FILL_4107
timestamp 1677677812
transform 1 0 2872 0 1 2970
box -8 -3 16 105
use FILL  FILL_4108
timestamp 1677677812
transform 1 0 2880 0 1 2970
box -8 -3 16 105
use FILL  FILL_4109
timestamp 1677677812
transform 1 0 2888 0 1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_45
timestamp 1677677812
transform 1 0 2896 0 1 2970
box -8 -3 32 105
use FILL  FILL_4110
timestamp 1677677812
transform 1 0 2920 0 1 2970
box -8 -3 16 105
use FILL  FILL_4115
timestamp 1677677812
transform 1 0 2928 0 1 2970
box -8 -3 16 105
use FILL  FILL_4116
timestamp 1677677812
transform 1 0 2936 0 1 2970
box -8 -3 16 105
use FILL  FILL_4117
timestamp 1677677812
transform 1 0 2944 0 1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_90
timestamp 1677677812
transform -1 0 2984 0 1 2970
box -8 -3 34 105
use FILL  FILL_4118
timestamp 1677677812
transform 1 0 2984 0 1 2970
box -8 -3 16 105
use FILL  FILL_4119
timestamp 1677677812
transform 1 0 2992 0 1 2970
box -8 -3 16 105
use FILL  FILL_4120
timestamp 1677677812
transform 1 0 3000 0 1 2970
box -8 -3 16 105
use FILL  FILL_4121
timestamp 1677677812
transform 1 0 3008 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_164
timestamp 1677677812
transform 1 0 3016 0 1 2970
box -8 -3 46 105
use FILL  FILL_4122
timestamp 1677677812
transform 1 0 3056 0 1 2970
box -8 -3 16 105
use FILL  FILL_4132
timestamp 1677677812
transform 1 0 3064 0 1 2970
box -8 -3 16 105
use FILL  FILL_4134
timestamp 1677677812
transform 1 0 3072 0 1 2970
box -8 -3 16 105
use FILL  FILL_4136
timestamp 1677677812
transform 1 0 3080 0 1 2970
box -8 -3 16 105
use FILL  FILL_4137
timestamp 1677677812
transform 1 0 3088 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_252
timestamp 1677677812
transform -1 0 3192 0 1 2970
box -8 -3 104 105
use FILL  FILL_4138
timestamp 1677677812
transform 1 0 3192 0 1 2970
box -8 -3 16 105
use FILL  FILL_4152
timestamp 1677677812
transform 1 0 3200 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_165
timestamp 1677677812
transform 1 0 3208 0 1 2970
box -8 -3 46 105
use FILL  FILL_4154
timestamp 1677677812
transform 1 0 3248 0 1 2970
box -8 -3 16 105
use FILL  FILL_4161
timestamp 1677677812
transform 1 0 3256 0 1 2970
box -8 -3 16 105
use FILL  FILL_4163
timestamp 1677677812
transform 1 0 3264 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3298
timestamp 1677677812
transform 1 0 3308 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3299
timestamp 1677677812
transform 1 0 3332 0 1 2975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_253
timestamp 1677677812
transform 1 0 3272 0 1 2970
box -8 -3 104 105
use FILL  FILL_4165
timestamp 1677677812
transform 1 0 3368 0 1 2970
box -8 -3 16 105
use FILL  FILL_4166
timestamp 1677677812
transform 1 0 3376 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_286
timestamp 1677677812
transform 1 0 3384 0 1 2970
box -9 -3 26 105
use FILL  FILL_4167
timestamp 1677677812
transform 1 0 3400 0 1 2970
box -8 -3 16 105
use FILL  FILL_4168
timestamp 1677677812
transform 1 0 3408 0 1 2970
box -8 -3 16 105
use FILL  FILL_4169
timestamp 1677677812
transform 1 0 3416 0 1 2970
box -8 -3 16 105
use NAND3X1  NAND3X1_23
timestamp 1677677812
transform -1 0 3456 0 1 2970
box -8 -3 40 105
use FILL  FILL_4170
timestamp 1677677812
transform 1 0 3456 0 1 2970
box -8 -3 16 105
use FILL  FILL_4181
timestamp 1677677812
transform 1 0 3464 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_255
timestamp 1677677812
transform 1 0 3472 0 1 2970
box -8 -3 104 105
use FILL  FILL_4183
timestamp 1677677812
transform 1 0 3568 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3300
timestamp 1677677812
transform 1 0 3612 0 1 2975
box -3 -3 3 3
use OAI22X1  OAI22X1_167
timestamp 1677677812
transform 1 0 3576 0 1 2970
box -8 -3 46 105
use FILL  FILL_4192
timestamp 1677677812
transform 1 0 3616 0 1 2970
box -8 -3 16 105
use FILL  FILL_4193
timestamp 1677677812
transform 1 0 3624 0 1 2970
box -8 -3 16 105
use FILL  FILL_4194
timestamp 1677677812
transform 1 0 3632 0 1 2970
box -8 -3 16 105
use FILL  FILL_4195
timestamp 1677677812
transform 1 0 3640 0 1 2970
box -8 -3 16 105
use FILL  FILL_4200
timestamp 1677677812
transform 1 0 3648 0 1 2970
box -8 -3 16 105
use FILL  FILL_4202
timestamp 1677677812
transform 1 0 3656 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_169
timestamp 1677677812
transform -1 0 3704 0 1 2970
box -8 -3 46 105
use FILL  FILL_4203
timestamp 1677677812
transform 1 0 3704 0 1 2970
box -8 -3 16 105
use FILL  FILL_4204
timestamp 1677677812
transform 1 0 3712 0 1 2970
box -8 -3 16 105
use FILL  FILL_4205
timestamp 1677677812
transform 1 0 3720 0 1 2970
box -8 -3 16 105
use FILL  FILL_4206
timestamp 1677677812
transform 1 0 3728 0 1 2970
box -8 -3 16 105
use FILL  FILL_4207
timestamp 1677677812
transform 1 0 3736 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_256
timestamp 1677677812
transform 1 0 3744 0 1 2970
box -8 -3 104 105
use FILL  FILL_4208
timestamp 1677677812
transform 1 0 3840 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_288
timestamp 1677677812
transform 1 0 3848 0 1 2970
box -9 -3 26 105
use BUFX2  BUFX2_30
timestamp 1677677812
transform 1 0 3864 0 1 2970
box -5 -3 28 105
use FILL  FILL_4221
timestamp 1677677812
transform 1 0 3888 0 1 2970
box -8 -3 16 105
use FILL  FILL_4222
timestamp 1677677812
transform 1 0 3896 0 1 2970
box -8 -3 16 105
use FILL  FILL_4223
timestamp 1677677812
transform 1 0 3904 0 1 2970
box -8 -3 16 105
use FILL  FILL_4224
timestamp 1677677812
transform 1 0 3912 0 1 2970
box -8 -3 16 105
use FILL  FILL_4225
timestamp 1677677812
transform 1 0 3920 0 1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_258
timestamp 1677677812
transform 1 0 3928 0 1 2970
box -8 -3 104 105
use INVX2  INVX2_289
timestamp 1677677812
transform 1 0 4024 0 1 2970
box -9 -3 26 105
use FILL  FILL_4226
timestamp 1677677812
transform 1 0 4040 0 1 2970
box -8 -3 16 105
use FILL  FILL_4242
timestamp 1677677812
transform 1 0 4048 0 1 2970
box -8 -3 16 105
use BUFX2  BUFX2_31
timestamp 1677677812
transform 1 0 4056 0 1 2970
box -5 -3 28 105
use FILL  FILL_4244
timestamp 1677677812
transform 1 0 4080 0 1 2970
box -8 -3 16 105
use FILL  FILL_4245
timestamp 1677677812
transform 1 0 4088 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3301
timestamp 1677677812
transform 1 0 4108 0 1 2975
box -3 -3 3 3
use FILL  FILL_4246
timestamp 1677677812
transform 1 0 4096 0 1 2970
box -8 -3 16 105
use FILL  FILL_4247
timestamp 1677677812
transform 1 0 4104 0 1 2970
box -8 -3 16 105
use FILL  FILL_4248
timestamp 1677677812
transform 1 0 4112 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_171
timestamp 1677677812
transform 1 0 4120 0 1 2970
box -8 -3 46 105
use FILL  FILL_4249
timestamp 1677677812
transform 1 0 4160 0 1 2970
box -8 -3 16 105
use FILL  FILL_4250
timestamp 1677677812
transform 1 0 4168 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3302
timestamp 1677677812
transform 1 0 4188 0 1 2975
box -3 -3 3 3
use M3_M2  M3_M2_3303
timestamp 1677677812
transform 1 0 4212 0 1 2975
box -3 -3 3 3
use AOI22X1  AOI22X1_180
timestamp 1677677812
transform -1 0 4216 0 1 2970
box -8 -3 46 105
use FILL  FILL_4251
timestamp 1677677812
transform 1 0 4216 0 1 2970
box -8 -3 16 105
use FILL  FILL_4252
timestamp 1677677812
transform 1 0 4224 0 1 2970
box -8 -3 16 105
use FILL  FILL_4253
timestamp 1677677812
transform 1 0 4232 0 1 2970
box -8 -3 16 105
use FILL  FILL_4254
timestamp 1677677812
transform 1 0 4240 0 1 2970
box -8 -3 16 105
use FILL  FILL_4255
timestamp 1677677812
transform 1 0 4248 0 1 2970
box -8 -3 16 105
use FILL  FILL_4256
timestamp 1677677812
transform 1 0 4256 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3304
timestamp 1677677812
transform 1 0 4284 0 1 2975
box -3 -3 3 3
use BUFX2  BUFX2_32
timestamp 1677677812
transform 1 0 4264 0 1 2970
box -5 -3 28 105
use FILL  FILL_4264
timestamp 1677677812
transform 1 0 4288 0 1 2970
box -8 -3 16 105
use FILL  FILL_4269
timestamp 1677677812
transform 1 0 4296 0 1 2970
box -8 -3 16 105
use FILL  FILL_4270
timestamp 1677677812
transform 1 0 4304 0 1 2970
box -8 -3 16 105
use FILL  FILL_4271
timestamp 1677677812
transform 1 0 4312 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_181
timestamp 1677677812
transform 1 0 4320 0 1 2970
box -8 -3 46 105
use FILL  FILL_4272
timestamp 1677677812
transform 1 0 4360 0 1 2970
box -8 -3 16 105
use FILL  FILL_4277
timestamp 1677677812
transform 1 0 4368 0 1 2970
box -8 -3 16 105
use FILL  FILL_4278
timestamp 1677677812
transform 1 0 4376 0 1 2970
box -8 -3 16 105
use FILL  FILL_4279
timestamp 1677677812
transform 1 0 4384 0 1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3305
timestamp 1677677812
transform 1 0 4404 0 1 2975
box -3 -3 3 3
use FILL  FILL_4280
timestamp 1677677812
transform 1 0 4392 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_174
timestamp 1677677812
transform 1 0 4400 0 1 2970
box -8 -3 46 105
use FILL  FILL_4281
timestamp 1677677812
transform 1 0 4440 0 1 2970
box -8 -3 16 105
use FILL  FILL_4282
timestamp 1677677812
transform 1 0 4448 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_291
timestamp 1677677812
transform -1 0 4472 0 1 2970
box -9 -3 26 105
use FILL  FILL_4283
timestamp 1677677812
transform 1 0 4472 0 1 2970
box -8 -3 16 105
use FILL  FILL_4284
timestamp 1677677812
transform 1 0 4480 0 1 2970
box -8 -3 16 105
use FILL  FILL_4285
timestamp 1677677812
transform 1 0 4488 0 1 2970
box -8 -3 16 105
use FILL  FILL_4288
timestamp 1677677812
transform 1 0 4496 0 1 2970
box -8 -3 16 105
use FILL  FILL_4289
timestamp 1677677812
transform 1 0 4504 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_175
timestamp 1677677812
transform 1 0 4512 0 1 2970
box -8 -3 46 105
use FILL  FILL_4290
timestamp 1677677812
transform 1 0 4552 0 1 2970
box -8 -3 16 105
use FILL  FILL_4291
timestamp 1677677812
transform 1 0 4560 0 1 2970
box -8 -3 16 105
use FILL  FILL_4292
timestamp 1677677812
transform 1 0 4568 0 1 2970
box -8 -3 16 105
use FILL  FILL_4293
timestamp 1677677812
transform 1 0 4576 0 1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_182
timestamp 1677677812
transform 1 0 4584 0 1 2970
box -8 -3 46 105
use FILL  FILL_4294
timestamp 1677677812
transform 1 0 4624 0 1 2970
box -8 -3 16 105
use FILL  FILL_4295
timestamp 1677677812
transform 1 0 4632 0 1 2970
box -8 -3 16 105
use FILL  FILL_4300
timestamp 1677677812
transform 1 0 4640 0 1 2970
box -8 -3 16 105
use FILL  FILL_4301
timestamp 1677677812
transform 1 0 4648 0 1 2970
box -8 -3 16 105
use FILL  FILL_4302
timestamp 1677677812
transform 1 0 4656 0 1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_176
timestamp 1677677812
transform 1 0 4664 0 1 2970
box -8 -3 46 105
use FILL  FILL_4303
timestamp 1677677812
transform 1 0 4704 0 1 2970
box -8 -3 16 105
use FILL  FILL_4304
timestamp 1677677812
transform 1 0 4712 0 1 2970
box -8 -3 16 105
use FILL  FILL_4305
timestamp 1677677812
transform 1 0 4720 0 1 2970
box -8 -3 16 105
use INVX2  INVX2_294
timestamp 1677677812
transform -1 0 4744 0 1 2970
box -9 -3 26 105
use FILL  FILL_4306
timestamp 1677677812
transform 1 0 4744 0 1 2970
box -8 -3 16 105
use FILL  FILL_4307
timestamp 1677677812
transform 1 0 4752 0 1 2970
box -8 -3 16 105
use FILL  FILL_4308
timestamp 1677677812
transform 1 0 4760 0 1 2970
box -8 -3 16 105
use FILL  FILL_4309
timestamp 1677677812
transform 1 0 4768 0 1 2970
box -8 -3 16 105
use FILL  FILL_4310
timestamp 1677677812
transform 1 0 4776 0 1 2970
box -8 -3 16 105
use FILL  FILL_4311
timestamp 1677677812
transform 1 0 4784 0 1 2970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_35
timestamp 1677677812
transform 1 0 4819 0 1 2970
box -10 -3 10 3
use M2_M1  M2_M1_3760
timestamp 1677677812
transform 1 0 84 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3306
timestamp 1677677812
transform 1 0 172 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3843
timestamp 1677677812
transform 1 0 108 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3844
timestamp 1677677812
transform 1 0 164 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3315
timestamp 1677677812
transform 1 0 188 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3316
timestamp 1677677812
transform 1 0 252 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3307
timestamp 1677677812
transform 1 0 308 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3308
timestamp 1677677812
transform 1 0 340 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3317
timestamp 1677677812
transform 1 0 356 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3346
timestamp 1677677812
transform 1 0 404 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3761
timestamp 1677677812
transform 1 0 188 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3762
timestamp 1677677812
transform 1 0 276 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3763
timestamp 1677677812
transform 1 0 300 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3764
timestamp 1677677812
transform 1 0 308 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3765
timestamp 1677677812
transform 1 0 324 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3845
timestamp 1677677812
transform 1 0 236 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3846
timestamp 1677677812
transform 1 0 268 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3847
timestamp 1677677812
transform 1 0 276 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3848
timestamp 1677677812
transform 1 0 292 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3439
timestamp 1677677812
transform 1 0 236 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3440
timestamp 1677677812
transform 1 0 268 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3366
timestamp 1677677812
transform 1 0 372 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3367
timestamp 1677677812
transform 1 0 412 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3849
timestamp 1677677812
transform 1 0 372 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3850
timestamp 1677677812
transform 1 0 404 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3851
timestamp 1677677812
transform 1 0 412 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3441
timestamp 1677677812
transform 1 0 308 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3468
timestamp 1677677812
transform 1 0 300 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3469
timestamp 1677677812
transform 1 0 332 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3393
timestamp 1677677812
transform 1 0 436 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3318
timestamp 1677677812
transform 1 0 476 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3347
timestamp 1677677812
transform 1 0 492 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3766
timestamp 1677677812
transform 1 0 468 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3767
timestamp 1677677812
transform 1 0 476 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3768
timestamp 1677677812
transform 1 0 492 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3852
timestamp 1677677812
transform 1 0 468 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3394
timestamp 1677677812
transform 1 0 476 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3853
timestamp 1677677812
transform 1 0 484 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3854
timestamp 1677677812
transform 1 0 500 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3416
timestamp 1677677812
transform 1 0 468 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3769
timestamp 1677677812
transform 1 0 532 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3855
timestamp 1677677812
transform 1 0 540 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3417
timestamp 1677677812
transform 1 0 540 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3470
timestamp 1677677812
transform 1 0 532 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3770
timestamp 1677677812
transform 1 0 572 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3856
timestamp 1677677812
transform 1 0 564 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3857
timestamp 1677677812
transform 1 0 580 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3442
timestamp 1677677812
transform 1 0 604 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3319
timestamp 1677677812
transform 1 0 628 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3320
timestamp 1677677812
transform 1 0 652 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3348
timestamp 1677677812
transform 1 0 668 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3771
timestamp 1677677812
transform 1 0 652 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3772
timestamp 1677677812
transform 1 0 668 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3858
timestamp 1677677812
transform 1 0 644 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3859
timestamp 1677677812
transform 1 0 660 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3395
timestamp 1677677812
transform 1 0 684 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3773
timestamp 1677677812
transform 1 0 724 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3368
timestamp 1677677812
transform 1 0 772 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3396
timestamp 1677677812
transform 1 0 724 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3369
timestamp 1677677812
transform 1 0 812 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3860
timestamp 1677677812
transform 1 0 772 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3861
timestamp 1677677812
transform 1 0 804 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3862
timestamp 1677677812
transform 1 0 812 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3471
timestamp 1677677812
transform 1 0 812 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3774
timestamp 1677677812
transform 1 0 836 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3321
timestamp 1677677812
transform 1 0 868 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3758
timestamp 1677677812
transform 1 0 868 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3443
timestamp 1677677812
transform 1 0 868 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3349
timestamp 1677677812
transform 1 0 1004 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3863
timestamp 1677677812
transform 1 0 1004 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3309
timestamp 1677677812
transform 1 0 1036 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3775
timestamp 1677677812
transform 1 0 1028 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3864
timestamp 1677677812
transform 1 0 1036 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3776
timestamp 1677677812
transform 1 0 1060 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3865
timestamp 1677677812
transform 1 0 1068 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3777
timestamp 1677677812
transform 1 0 1084 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3778
timestamp 1677677812
transform 1 0 1092 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3866
timestamp 1677677812
transform 1 0 1092 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3418
timestamp 1677677812
transform 1 0 1092 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3444
timestamp 1677677812
transform 1 0 1092 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3867
timestamp 1677677812
transform 1 0 1148 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3419
timestamp 1677677812
transform 1 0 1148 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3868
timestamp 1677677812
transform 1 0 1172 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3869
timestamp 1677677812
transform 1 0 1188 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3445
timestamp 1677677812
transform 1 0 1188 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3870
timestamp 1677677812
transform 1 0 1228 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3779
timestamp 1677677812
transform 1 0 1260 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3350
timestamp 1677677812
transform 1 0 1308 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3780
timestamp 1677677812
transform 1 0 1308 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3781
timestamp 1677677812
transform 1 0 1316 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3936
timestamp 1677677812
transform 1 0 1324 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3446
timestamp 1677677812
transform 1 0 1324 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3472
timestamp 1677677812
transform 1 0 1316 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3370
timestamp 1677677812
transform 1 0 1340 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3937
timestamp 1677677812
transform 1 0 1340 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3322
timestamp 1677677812
transform 1 0 1364 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3871
timestamp 1677677812
transform 1 0 1364 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3782
timestamp 1677677812
transform 1 0 1380 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3371
timestamp 1677677812
transform 1 0 1388 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3783
timestamp 1677677812
transform 1 0 1404 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3397
timestamp 1677677812
transform 1 0 1396 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3938
timestamp 1677677812
transform 1 0 1388 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3447
timestamp 1677677812
transform 1 0 1404 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3462
timestamp 1677677812
transform 1 0 1404 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3323
timestamp 1677677812
transform 1 0 1444 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3872
timestamp 1677677812
transform 1 0 1444 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3351
timestamp 1677677812
transform 1 0 1492 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3784
timestamp 1677677812
transform 1 0 1492 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3352
timestamp 1677677812
transform 1 0 1588 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3785
timestamp 1677677812
transform 1 0 1508 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3372
timestamp 1677677812
transform 1 0 1556 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3373
timestamp 1677677812
transform 1 0 1580 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3398
timestamp 1677677812
transform 1 0 1508 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3873
timestamp 1677677812
transform 1 0 1556 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3353
timestamp 1677677812
transform 1 0 1628 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3874
timestamp 1677677812
transform 1 0 1628 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3786
timestamp 1677677812
transform 1 0 1660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3875
timestamp 1677677812
transform 1 0 1668 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3787
timestamp 1677677812
transform 1 0 1684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3876
timestamp 1677677812
transform 1 0 1748 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3788
timestamp 1677677812
transform 1 0 1772 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3877
timestamp 1677677812
transform 1 0 1812 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3399
timestamp 1677677812
transform 1 0 1836 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3420
timestamp 1677677812
transform 1 0 1796 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3473
timestamp 1677677812
transform 1 0 1804 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3474
timestamp 1677677812
transform 1 0 1828 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3789
timestamp 1677677812
transform 1 0 1860 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3400
timestamp 1677677812
transform 1 0 1860 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3374
timestamp 1677677812
transform 1 0 1876 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3878
timestamp 1677677812
transform 1 0 1868 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3879
timestamp 1677677812
transform 1 0 1876 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3324
timestamp 1677677812
transform 1 0 1900 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3325
timestamp 1677677812
transform 1 0 1932 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3790
timestamp 1677677812
transform 1 0 1908 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3791
timestamp 1677677812
transform 1 0 1924 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3792
timestamp 1677677812
transform 1 0 1932 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3880
timestamp 1677677812
transform 1 0 1916 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3881
timestamp 1677677812
transform 1 0 1956 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3375
timestamp 1677677812
transform 1 0 1980 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3882
timestamp 1677677812
transform 1 0 1980 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3401
timestamp 1677677812
transform 1 0 1988 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3354
timestamp 1677677812
transform 1 0 2004 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3326
timestamp 1677677812
transform 1 0 2036 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3793
timestamp 1677677812
transform 1 0 2012 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3794
timestamp 1677677812
transform 1 0 2020 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3795
timestamp 1677677812
transform 1 0 2036 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3402
timestamp 1677677812
transform 1 0 2020 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3883
timestamp 1677677812
transform 1 0 2028 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3376
timestamp 1677677812
transform 1 0 2068 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3884
timestamp 1677677812
transform 1 0 2060 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3885
timestamp 1677677812
transform 1 0 2068 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3327
timestamp 1677677812
transform 1 0 2108 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3796
timestamp 1677677812
transform 1 0 2092 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3797
timestamp 1677677812
transform 1 0 2108 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3798
timestamp 1677677812
transform 1 0 2116 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3886
timestamp 1677677812
transform 1 0 2100 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3421
timestamp 1677677812
transform 1 0 2084 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3403
timestamp 1677677812
transform 1 0 2116 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3887
timestamp 1677677812
transform 1 0 2124 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3377
timestamp 1677677812
transform 1 0 2140 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3888
timestamp 1677677812
transform 1 0 2140 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3422
timestamp 1677677812
transform 1 0 2140 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3328
timestamp 1677677812
transform 1 0 2180 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3799
timestamp 1677677812
transform 1 0 2180 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3889
timestamp 1677677812
transform 1 0 2172 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3378
timestamp 1677677812
transform 1 0 2196 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3890
timestamp 1677677812
transform 1 0 2196 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3404
timestamp 1677677812
transform 1 0 2204 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3463
timestamp 1677677812
transform 1 0 2196 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3464
timestamp 1677677812
transform 1 0 2220 0 1 2895
box -3 -3 3 3
use M2_M1  M2_M1_3800
timestamp 1677677812
transform 1 0 2236 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3379
timestamp 1677677812
transform 1 0 2260 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3891
timestamp 1677677812
transform 1 0 2260 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3892
timestamp 1677677812
transform 1 0 2316 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3423
timestamp 1677677812
transform 1 0 2276 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3465
timestamp 1677677812
transform 1 0 2252 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3329
timestamp 1677677812
transform 1 0 2332 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3448
timestamp 1677677812
transform 1 0 2340 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3754
timestamp 1677677812
transform 1 0 2380 0 1 2955
box -2 -2 2 2
use M3_M2  M3_M2_3424
timestamp 1677677812
transform 1 0 2404 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3755
timestamp 1677677812
transform 1 0 2420 0 1 2955
box -2 -2 2 2
use M2_M1  M2_M1_3893
timestamp 1677677812
transform 1 0 2444 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3330
timestamp 1677677812
transform 1 0 2508 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3380
timestamp 1677677812
transform 1 0 2476 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3801
timestamp 1677677812
transform 1 0 2540 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3894
timestamp 1677677812
transform 1 0 2492 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3449
timestamp 1677677812
transform 1 0 2540 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3331
timestamp 1677677812
transform 1 0 2556 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3802
timestamp 1677677812
transform 1 0 2556 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3895
timestamp 1677677812
transform 1 0 2564 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3332
timestamp 1677677812
transform 1 0 2612 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3803
timestamp 1677677812
transform 1 0 2604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3804
timestamp 1677677812
transform 1 0 2612 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3896
timestamp 1677677812
transform 1 0 2596 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3405
timestamp 1677677812
transform 1 0 2604 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3897
timestamp 1677677812
transform 1 0 2620 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3450
timestamp 1677677812
transform 1 0 2636 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3898
timestamp 1677677812
transform 1 0 2668 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3425
timestamp 1677677812
transform 1 0 2668 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3805
timestamp 1677677812
transform 1 0 2684 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3899
timestamp 1677677812
transform 1 0 2708 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3406
timestamp 1677677812
transform 1 0 2756 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3759
timestamp 1677677812
transform 1 0 2772 0 1 2945
box -2 -2 2 2
use M3_M2  M3_M2_3381
timestamp 1677677812
transform 1 0 2772 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3900
timestamp 1677677812
transform 1 0 2764 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3426
timestamp 1677677812
transform 1 0 2708 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3333
timestamp 1677677812
transform 1 0 2844 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3355
timestamp 1677677812
transform 1 0 2852 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3806
timestamp 1677677812
transform 1 0 2836 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3807
timestamp 1677677812
transform 1 0 2844 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3901
timestamp 1677677812
transform 1 0 2844 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3902
timestamp 1677677812
transform 1 0 2868 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3427
timestamp 1677677812
transform 1 0 2868 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3939
timestamp 1677677812
transform 1 0 2892 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3451
timestamp 1677677812
transform 1 0 2900 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3808
timestamp 1677677812
transform 1 0 2916 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3809
timestamp 1677677812
transform 1 0 2924 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3903
timestamp 1677677812
transform 1 0 2916 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3407
timestamp 1677677812
transform 1 0 2924 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3428
timestamp 1677677812
transform 1 0 2916 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3452
timestamp 1677677812
transform 1 0 2932 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3810
timestamp 1677677812
transform 1 0 2956 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3940
timestamp 1677677812
transform 1 0 2972 0 1 2915
box -2 -2 2 2
use M3_M2  M3_M2_3453
timestamp 1677677812
transform 1 0 2972 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3904
timestamp 1677677812
transform 1 0 3004 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3905
timestamp 1677677812
transform 1 0 3044 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3475
timestamp 1677677812
transform 1 0 3060 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3476
timestamp 1677677812
transform 1 0 3076 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3811
timestamp 1677677812
transform 1 0 3100 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3429
timestamp 1677677812
transform 1 0 3092 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3466
timestamp 1677677812
transform 1 0 3180 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3430
timestamp 1677677812
transform 1 0 3204 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3454
timestamp 1677677812
transform 1 0 3308 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3334
timestamp 1677677812
transform 1 0 3364 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3335
timestamp 1677677812
transform 1 0 3380 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3356
timestamp 1677677812
transform 1 0 3380 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3812
timestamp 1677677812
transform 1 0 3332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3906
timestamp 1677677812
transform 1 0 3380 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3431
timestamp 1677677812
transform 1 0 3332 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3455
timestamp 1677677812
transform 1 0 3324 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3467
timestamp 1677677812
transform 1 0 3332 0 1 2895
box -3 -3 3 3
use M3_M2  M3_M2_3310
timestamp 1677677812
transform 1 0 3436 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3813
timestamp 1677677812
transform 1 0 3444 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3336
timestamp 1677677812
transform 1 0 3468 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3814
timestamp 1677677812
transform 1 0 3468 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3337
timestamp 1677677812
transform 1 0 3508 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3357
timestamp 1677677812
transform 1 0 3500 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3382
timestamp 1677677812
transform 1 0 3492 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3815
timestamp 1677677812
transform 1 0 3500 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3907
timestamp 1677677812
transform 1 0 3484 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3908
timestamp 1677677812
transform 1 0 3492 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3909
timestamp 1677677812
transform 1 0 3508 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3456
timestamp 1677677812
transform 1 0 3508 0 1 2905
box -3 -3 3 3
use M2_M1  M2_M1_3816
timestamp 1677677812
transform 1 0 3540 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3383
timestamp 1677677812
transform 1 0 3548 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3408
timestamp 1677677812
transform 1 0 3556 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3457
timestamp 1677677812
transform 1 0 3564 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3384
timestamp 1677677812
transform 1 0 3588 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3311
timestamp 1677677812
transform 1 0 3612 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3338
timestamp 1677677812
transform 1 0 3604 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3358
timestamp 1677677812
transform 1 0 3620 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3817
timestamp 1677677812
transform 1 0 3596 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3818
timestamp 1677677812
transform 1 0 3604 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3819
timestamp 1677677812
transform 1 0 3620 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3820
timestamp 1677677812
transform 1 0 3636 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3409
timestamp 1677677812
transform 1 0 3596 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3910
timestamp 1677677812
transform 1 0 3612 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3911
timestamp 1677677812
transform 1 0 3628 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3410
timestamp 1677677812
transform 1 0 3636 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3312
timestamp 1677677812
transform 1 0 3652 0 1 2965
box -3 -3 3 3
use M2_M1  M2_M1_3912
timestamp 1677677812
transform 1 0 3668 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3313
timestamp 1677677812
transform 1 0 3708 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3339
timestamp 1677677812
transform 1 0 3716 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3340
timestamp 1677677812
transform 1 0 3756 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3359
timestamp 1677677812
transform 1 0 3708 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3821
timestamp 1677677812
transform 1 0 3756 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3913
timestamp 1677677812
transform 1 0 3708 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3914
timestamp 1677677812
transform 1 0 3884 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3822
timestamp 1677677812
transform 1 0 3900 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3385
timestamp 1677677812
transform 1 0 3908 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3915
timestamp 1677677812
transform 1 0 3908 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3916
timestamp 1677677812
transform 1 0 3924 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3756
timestamp 1677677812
transform 1 0 3940 0 1 2955
box -2 -2 2 2
use M2_M1  M2_M1_3757
timestamp 1677677812
transform 1 0 3972 0 1 2955
box -2 -2 2 2
use M2_M1  M2_M1_3823
timestamp 1677677812
transform 1 0 3956 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3824
timestamp 1677677812
transform 1 0 3964 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3477
timestamp 1677677812
transform 1 0 3964 0 1 2885
box -3 -3 3 3
use M2_M1  M2_M1_3825
timestamp 1677677812
transform 1 0 4020 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3386
timestamp 1677677812
transform 1 0 4028 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3826
timestamp 1677677812
transform 1 0 4036 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3917
timestamp 1677677812
transform 1 0 4012 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3918
timestamp 1677677812
transform 1 0 4028 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3478
timestamp 1677677812
transform 1 0 4044 0 1 2885
box -3 -3 3 3
use M3_M2  M3_M2_3360
timestamp 1677677812
transform 1 0 4132 0 1 2945
box -3 -3 3 3
use M3_M2  M3_M2_3361
timestamp 1677677812
transform 1 0 4148 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3827
timestamp 1677677812
transform 1 0 4164 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3919
timestamp 1677677812
transform 1 0 4084 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3920
timestamp 1677677812
transform 1 0 4140 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3432
timestamp 1677677812
transform 1 0 4164 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3828
timestamp 1677677812
transform 1 0 4188 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3314
timestamp 1677677812
transform 1 0 4212 0 1 2965
box -3 -3 3 3
use M3_M2  M3_M2_3341
timestamp 1677677812
transform 1 0 4220 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3362
timestamp 1677677812
transform 1 0 4236 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3829
timestamp 1677677812
transform 1 0 4220 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3387
timestamp 1677677812
transform 1 0 4228 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3830
timestamp 1677677812
transform 1 0 4236 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3831
timestamp 1677677812
transform 1 0 4244 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3921
timestamp 1677677812
transform 1 0 4212 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3922
timestamp 1677677812
transform 1 0 4228 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3411
timestamp 1677677812
transform 1 0 4236 0 1 2925
box -3 -3 3 3
use M3_M2  M3_M2_3458
timestamp 1677677812
transform 1 0 4212 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3388
timestamp 1677677812
transform 1 0 4252 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3923
timestamp 1677677812
transform 1 0 4252 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3342
timestamp 1677677812
transform 1 0 4268 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3832
timestamp 1677677812
transform 1 0 4284 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3363
timestamp 1677677812
transform 1 0 4332 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3833
timestamp 1677677812
transform 1 0 4316 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3389
timestamp 1677677812
transform 1 0 4324 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3834
timestamp 1677677812
transform 1 0 4332 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3924
timestamp 1677677812
transform 1 0 4308 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3925
timestamp 1677677812
transform 1 0 4324 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3459
timestamp 1677677812
transform 1 0 4308 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3390
timestamp 1677677812
transform 1 0 4356 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3926
timestamp 1677677812
transform 1 0 4356 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3343
timestamp 1677677812
transform 1 0 4404 0 1 2955
box -3 -3 3 3
use M2_M1  M2_M1_3835
timestamp 1677677812
transform 1 0 4388 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3836
timestamp 1677677812
transform 1 0 4404 0 1 2935
box -2 -2 2 2
use M3_M2  M3_M2_3412
timestamp 1677677812
transform 1 0 4388 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3927
timestamp 1677677812
transform 1 0 4428 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3413
timestamp 1677677812
transform 1 0 4436 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3928
timestamp 1677677812
transform 1 0 4484 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3433
timestamp 1677677812
transform 1 0 4404 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3434
timestamp 1677677812
transform 1 0 4428 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3435
timestamp 1677677812
transform 1 0 4468 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3460
timestamp 1677677812
transform 1 0 4444 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3461
timestamp 1677677812
transform 1 0 4476 0 1 2905
box -3 -3 3 3
use M3_M2  M3_M2_3364
timestamp 1677677812
transform 1 0 4548 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3837
timestamp 1677677812
transform 1 0 4508 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3929
timestamp 1677677812
transform 1 0 4532 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3436
timestamp 1677677812
transform 1 0 4540 0 1 2915
box -3 -3 3 3
use M2_M1  M2_M1_3930
timestamp 1677677812
transform 1 0 4628 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3344
timestamp 1677677812
transform 1 0 4684 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3345
timestamp 1677677812
transform 1 0 4716 0 1 2955
box -3 -3 3 3
use M3_M2  M3_M2_3365
timestamp 1677677812
transform 1 0 4692 0 1 2945
box -3 -3 3 3
use M2_M1  M2_M1_3838
timestamp 1677677812
transform 1 0 4644 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3839
timestamp 1677677812
transform 1 0 4660 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3840
timestamp 1677677812
transform 1 0 4676 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3841
timestamp 1677677812
transform 1 0 4692 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3842
timestamp 1677677812
transform 1 0 4780 0 1 2935
box -2 -2 2 2
use M2_M1  M2_M1_3931
timestamp 1677677812
transform 1 0 4652 0 1 2925
box -2 -2 2 2
use M2_M1  M2_M1_3932
timestamp 1677677812
transform 1 0 4668 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3437
timestamp 1677677812
transform 1 0 4668 0 1 2915
box -3 -3 3 3
use M3_M2  M3_M2_3391
timestamp 1677677812
transform 1 0 4788 0 1 2935
box -3 -3 3 3
use M3_M2  M3_M2_3392
timestamp 1677677812
transform 1 0 4804 0 1 2935
box -3 -3 3 3
use M2_M1  M2_M1_3933
timestamp 1677677812
transform 1 0 4716 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3414
timestamp 1677677812
transform 1 0 4764 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3934
timestamp 1677677812
transform 1 0 4772 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3415
timestamp 1677677812
transform 1 0 4780 0 1 2925
box -3 -3 3 3
use M2_M1  M2_M1_3935
timestamp 1677677812
transform 1 0 4788 0 1 2925
box -2 -2 2 2
use M3_M2  M3_M2_3438
timestamp 1677677812
transform 1 0 4788 0 1 2915
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_36
timestamp 1677677812
transform 1 0 24 0 1 2870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_238
timestamp 1677677812
transform 1 0 72 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3810
timestamp 1677677812
transform 1 0 168 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_239
timestamp 1677677812
transform 1 0 176 0 -1 2970
box -8 -3 104 105
use AOI22X1  AOI22X1_164
timestamp 1677677812
transform -1 0 312 0 -1 2970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_240
timestamp 1677677812
transform 1 0 312 0 -1 2970
box -8 -3 104 105
use INVX2  INVX2_271
timestamp 1677677812
transform -1 0 424 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3811
timestamp 1677677812
transform 1 0 424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3813
timestamp 1677677812
transform 1 0 432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3815
timestamp 1677677812
transform 1 0 440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3817
timestamp 1677677812
transform 1 0 448 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3819
timestamp 1677677812
transform 1 0 456 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_165
timestamp 1677677812
transform 1 0 464 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3824
timestamp 1677677812
transform 1 0 504 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3825
timestamp 1677677812
transform 1 0 512 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3826
timestamp 1677677812
transform 1 0 520 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3827
timestamp 1677677812
transform 1 0 528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3828
timestamp 1677677812
transform 1 0 536 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_166
timestamp 1677677812
transform 1 0 544 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3829
timestamp 1677677812
transform 1 0 584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3831
timestamp 1677677812
transform 1 0 592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3833
timestamp 1677677812
transform 1 0 600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3835
timestamp 1677677812
transform 1 0 608 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3837
timestamp 1677677812
transform 1 0 616 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3839
timestamp 1677677812
transform 1 0 624 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_158
timestamp 1677677812
transform 1 0 632 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3842
timestamp 1677677812
transform 1 0 672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3843
timestamp 1677677812
transform 1 0 680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3845
timestamp 1677677812
transform 1 0 688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3847
timestamp 1677677812
transform 1 0 696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3849
timestamp 1677677812
transform 1 0 704 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_242
timestamp 1677677812
transform 1 0 712 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3860
timestamp 1677677812
transform 1 0 808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3861
timestamp 1677677812
transform 1 0 816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3862
timestamp 1677677812
transform 1 0 824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3864
timestamp 1677677812
transform 1 0 832 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3479
timestamp 1677677812
transform 1 0 868 0 1 2875
box -3 -3 3 3
use INVX2  INVX2_273
timestamp 1677677812
transform 1 0 840 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3868
timestamp 1677677812
transform 1 0 856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3870
timestamp 1677677812
transform 1 0 864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3872
timestamp 1677677812
transform 1 0 872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3873
timestamp 1677677812
transform 1 0 880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3874
timestamp 1677677812
transform 1 0 888 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3875
timestamp 1677677812
transform 1 0 896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3876
timestamp 1677677812
transform 1 0 904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3878
timestamp 1677677812
transform 1 0 912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3880
timestamp 1677677812
transform 1 0 920 0 -1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_41
timestamp 1677677812
transform 1 0 928 0 -1 2970
box -8 -3 32 105
use FILL  FILL_3885
timestamp 1677677812
transform 1 0 952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3886
timestamp 1677677812
transform 1 0 960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3887
timestamp 1677677812
transform 1 0 968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3888
timestamp 1677677812
transform 1 0 976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3890
timestamp 1677677812
transform 1 0 984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3892
timestamp 1677677812
transform 1 0 992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3894
timestamp 1677677812
transform 1 0 1000 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3896
timestamp 1677677812
transform 1 0 1008 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_167
timestamp 1677677812
transform 1 0 1016 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3904
timestamp 1677677812
transform 1 0 1056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3905
timestamp 1677677812
transform 1 0 1064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3906
timestamp 1677677812
transform 1 0 1072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3907
timestamp 1677677812
transform 1 0 1080 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3908
timestamp 1677677812
transform 1 0 1088 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3909
timestamp 1677677812
transform 1 0 1096 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3910
timestamp 1677677812
transform 1 0 1104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3911
timestamp 1677677812
transform 1 0 1112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3912
timestamp 1677677812
transform 1 0 1120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3913
timestamp 1677677812
transform 1 0 1128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3914
timestamp 1677677812
transform 1 0 1136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3915
timestamp 1677677812
transform 1 0 1144 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_168
timestamp 1677677812
transform 1 0 1152 0 -1 2970
box -8 -3 46 105
use FILL  FILL_3916
timestamp 1677677812
transform 1 0 1192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3917
timestamp 1677677812
transform 1 0 1200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3919
timestamp 1677677812
transform 1 0 1208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3921
timestamp 1677677812
transform 1 0 1216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3923
timestamp 1677677812
transform 1 0 1224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3925
timestamp 1677677812
transform 1 0 1232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3929
timestamp 1677677812
transform 1 0 1240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3930
timestamp 1677677812
transform 1 0 1248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3931
timestamp 1677677812
transform 1 0 1256 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_84
timestamp 1677677812
transform 1 0 1264 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3932
timestamp 1677677812
transform 1 0 1296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3934
timestamp 1677677812
transform 1 0 1304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3936
timestamp 1677677812
transform 1 0 1312 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3938
timestamp 1677677812
transform 1 0 1320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3940
timestamp 1677677812
transform 1 0 1328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3942
timestamp 1677677812
transform 1 0 1336 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_86
timestamp 1677677812
transform -1 0 1376 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3944
timestamp 1677677812
transform 1 0 1376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3946
timestamp 1677677812
transform 1 0 1384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3948
timestamp 1677677812
transform 1 0 1392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3950
timestamp 1677677812
transform 1 0 1400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3959
timestamp 1677677812
transform 1 0 1408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3960
timestamp 1677677812
transform 1 0 1416 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_87
timestamp 1677677812
transform -1 0 1456 0 -1 2970
box -8 -3 34 105
use FILL  FILL_3961
timestamp 1677677812
transform 1 0 1456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3962
timestamp 1677677812
transform 1 0 1464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3963
timestamp 1677677812
transform 1 0 1472 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3964
timestamp 1677677812
transform 1 0 1480 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3965
timestamp 1677677812
transform 1 0 1488 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_245
timestamp 1677677812
transform 1 0 1496 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3966
timestamp 1677677812
transform 1 0 1592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3967
timestamp 1677677812
transform 1 0 1600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3969
timestamp 1677677812
transform 1 0 1608 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_275
timestamp 1677677812
transform 1 0 1616 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3973
timestamp 1677677812
transform 1 0 1632 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3975
timestamp 1677677812
transform 1 0 1640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3978
timestamp 1677677812
transform 1 0 1648 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_276
timestamp 1677677812
transform 1 0 1656 0 -1 2970
box -9 -3 26 105
use FILL  FILL_3979
timestamp 1677677812
transform 1 0 1672 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3980
timestamp 1677677812
transform 1 0 1680 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3981
timestamp 1677677812
transform 1 0 1688 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3982
timestamp 1677677812
transform 1 0 1696 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3988
timestamp 1677677812
transform 1 0 1704 0 -1 2970
box -8 -3 16 105
use BUFX2  BUFX2_27
timestamp 1677677812
transform -1 0 1736 0 -1 2970
box -5 -3 28 105
use FILL  FILL_3989
timestamp 1677677812
transform 1 0 1736 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3995
timestamp 1677677812
transform 1 0 1744 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3996
timestamp 1677677812
transform 1 0 1752 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_246
timestamp 1677677812
transform 1 0 1760 0 -1 2970
box -8 -3 104 105
use FILL  FILL_3997
timestamp 1677677812
transform 1 0 1856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_3999
timestamp 1677677812
transform 1 0 1864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4001
timestamp 1677677812
transform 1 0 1872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4003
timestamp 1677677812
transform 1 0 1880 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4007
timestamp 1677677812
transform 1 0 1888 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_171
timestamp 1677677812
transform -1 0 1936 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4008
timestamp 1677677812
transform 1 0 1936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4009
timestamp 1677677812
transform 1 0 1944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4011
timestamp 1677677812
transform 1 0 1952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4020
timestamp 1677677812
transform 1 0 1960 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_279
timestamp 1677677812
transform -1 0 1984 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4021
timestamp 1677677812
transform 1 0 1984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4022
timestamp 1677677812
transform 1 0 1992 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4023
timestamp 1677677812
transform 1 0 2000 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_172
timestamp 1677677812
transform -1 0 2048 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4024
timestamp 1677677812
transform 1 0 2048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4025
timestamp 1677677812
transform 1 0 2056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4026
timestamp 1677677812
transform 1 0 2064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4027
timestamp 1677677812
transform 1 0 2072 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3480
timestamp 1677677812
transform 1 0 2124 0 1 2875
box -3 -3 3 3
use AOI22X1  AOI22X1_173
timestamp 1677677812
transform -1 0 2120 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4028
timestamp 1677677812
transform 1 0 2120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4029
timestamp 1677677812
transform 1 0 2128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4030
timestamp 1677677812
transform 1 0 2136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4031
timestamp 1677677812
transform 1 0 2144 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_174
timestamp 1677677812
transform -1 0 2192 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4032
timestamp 1677677812
transform 1 0 2192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4033
timestamp 1677677812
transform 1 0 2200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4034
timestamp 1677677812
transform 1 0 2208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4041
timestamp 1677677812
transform 1 0 2216 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_248
timestamp 1677677812
transform 1 0 2224 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4042
timestamp 1677677812
transform 1 0 2320 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4043
timestamp 1677677812
transform 1 0 2328 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4044
timestamp 1677677812
transform 1 0 2336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4046
timestamp 1677677812
transform 1 0 2344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4048
timestamp 1677677812
transform 1 0 2352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4049
timestamp 1677677812
transform 1 0 2360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4050
timestamp 1677677812
transform 1 0 2368 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4051
timestamp 1677677812
transform 1 0 2376 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4052
timestamp 1677677812
transform 1 0 2384 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4053
timestamp 1677677812
transform 1 0 2392 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4054
timestamp 1677677812
transform 1 0 2400 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4055
timestamp 1677677812
transform 1 0 2408 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4057
timestamp 1677677812
transform 1 0 2416 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4059
timestamp 1677677812
transform 1 0 2424 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4069
timestamp 1677677812
transform 1 0 2432 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4070
timestamp 1677677812
transform 1 0 2440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4071
timestamp 1677677812
transform 1 0 2448 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3481
timestamp 1677677812
transform 1 0 2500 0 1 2875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_249
timestamp 1677677812
transform -1 0 2552 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4072
timestamp 1677677812
transform 1 0 2552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4074
timestamp 1677677812
transform 1 0 2560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4087
timestamp 1677677812
transform 1 0 2568 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_178
timestamp 1677677812
transform 1 0 2576 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4088
timestamp 1677677812
transform 1 0 2616 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4089
timestamp 1677677812
transform 1 0 2624 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4090
timestamp 1677677812
transform 1 0 2632 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_284
timestamp 1677677812
transform 1 0 2640 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4091
timestamp 1677677812
transform 1 0 2656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4092
timestamp 1677677812
transform 1 0 2664 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_251
timestamp 1677677812
transform 1 0 2672 0 -1 2970
box -8 -3 104 105
use M3_M2  M3_M2_3482
timestamp 1677677812
transform 1 0 2780 0 1 2875
box -3 -3 3 3
use FILL  FILL_4093
timestamp 1677677812
transform 1 0 2768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4095
timestamp 1677677812
transform 1 0 2776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4097
timestamp 1677677812
transform 1 0 2784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4098
timestamp 1677677812
transform 1 0 2792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4099
timestamp 1677677812
transform 1 0 2800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4100
timestamp 1677677812
transform 1 0 2808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4101
timestamp 1677677812
transform 1 0 2816 0 -1 2970
box -8 -3 16 105
use NOR2X1  NOR2X1_44
timestamp 1677677812
transform 1 0 2824 0 -1 2970
box -8 -3 32 105
use FILL  FILL_4104
timestamp 1677677812
transform 1 0 2848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4105
timestamp 1677677812
transform 1 0 2856 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_89
timestamp 1677677812
transform 1 0 2864 0 -1 2970
box -8 -3 34 105
use FILL  FILL_4111
timestamp 1677677812
transform 1 0 2896 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4112
timestamp 1677677812
transform 1 0 2904 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4113
timestamp 1677677812
transform 1 0 2912 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4114
timestamp 1677677812
transform 1 0 2920 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_91
timestamp 1677677812
transform 1 0 2928 0 -1 2970
box -8 -3 34 105
use FILL  FILL_4123
timestamp 1677677812
transform 1 0 2960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4124
timestamp 1677677812
transform 1 0 2968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4125
timestamp 1677677812
transform 1 0 2976 0 -1 2970
box -8 -3 16 105
use OAI21X1  OAI21X1_92
timestamp 1677677812
transform -1 0 3016 0 -1 2970
box -8 -3 34 105
use FILL  FILL_4126
timestamp 1677677812
transform 1 0 3016 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4127
timestamp 1677677812
transform 1 0 3024 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4128
timestamp 1677677812
transform 1 0 3032 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4129
timestamp 1677677812
transform 1 0 3040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4130
timestamp 1677677812
transform 1 0 3048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4131
timestamp 1677677812
transform 1 0 3056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4133
timestamp 1677677812
transform 1 0 3064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4135
timestamp 1677677812
transform 1 0 3072 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4139
timestamp 1677677812
transform 1 0 3080 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_285
timestamp 1677677812
transform -1 0 3104 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4140
timestamp 1677677812
transform 1 0 3104 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4141
timestamp 1677677812
transform 1 0 3112 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4142
timestamp 1677677812
transform 1 0 3120 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4143
timestamp 1677677812
transform 1 0 3128 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4144
timestamp 1677677812
transform 1 0 3136 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4145
timestamp 1677677812
transform 1 0 3144 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4146
timestamp 1677677812
transform 1 0 3152 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4147
timestamp 1677677812
transform 1 0 3160 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4148
timestamp 1677677812
transform 1 0 3168 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4149
timestamp 1677677812
transform 1 0 3176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4150
timestamp 1677677812
transform 1 0 3184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4151
timestamp 1677677812
transform 1 0 3192 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4153
timestamp 1677677812
transform 1 0 3200 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4155
timestamp 1677677812
transform 1 0 3208 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4156
timestamp 1677677812
transform 1 0 3216 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4157
timestamp 1677677812
transform 1 0 3224 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4158
timestamp 1677677812
transform 1 0 3232 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4159
timestamp 1677677812
transform 1 0 3240 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4160
timestamp 1677677812
transform 1 0 3248 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4162
timestamp 1677677812
transform 1 0 3256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4164
timestamp 1677677812
transform 1 0 3264 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4171
timestamp 1677677812
transform 1 0 3272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4172
timestamp 1677677812
transform 1 0 3280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4173
timestamp 1677677812
transform 1 0 3288 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4174
timestamp 1677677812
transform 1 0 3296 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4175
timestamp 1677677812
transform 1 0 3304 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4176
timestamp 1677677812
transform 1 0 3312 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_254
timestamp 1677677812
transform 1 0 3320 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4177
timestamp 1677677812
transform 1 0 3416 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_287
timestamp 1677677812
transform 1 0 3424 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4178
timestamp 1677677812
transform 1 0 3440 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4179
timestamp 1677677812
transform 1 0 3448 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4180
timestamp 1677677812
transform 1 0 3456 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4182
timestamp 1677677812
transform 1 0 3464 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4184
timestamp 1677677812
transform 1 0 3472 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_166
timestamp 1677677812
transform 1 0 3480 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4185
timestamp 1677677812
transform 1 0 3520 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4186
timestamp 1677677812
transform 1 0 3528 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4187
timestamp 1677677812
transform 1 0 3536 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4188
timestamp 1677677812
transform 1 0 3544 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4189
timestamp 1677677812
transform 1 0 3552 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4190
timestamp 1677677812
transform 1 0 3560 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4191
timestamp 1677677812
transform 1 0 3568 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4196
timestamp 1677677812
transform 1 0 3576 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4197
timestamp 1677677812
transform 1 0 3584 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4198
timestamp 1677677812
transform 1 0 3592 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_168
timestamp 1677677812
transform 1 0 3600 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4199
timestamp 1677677812
transform 1 0 3640 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4201
timestamp 1677677812
transform 1 0 3648 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4209
timestamp 1677677812
transform 1 0 3656 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4210
timestamp 1677677812
transform 1 0 3664 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_257
timestamp 1677677812
transform -1 0 3768 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4211
timestamp 1677677812
transform 1 0 3768 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4212
timestamp 1677677812
transform 1 0 3776 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4213
timestamp 1677677812
transform 1 0 3784 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4214
timestamp 1677677812
transform 1 0 3792 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4215
timestamp 1677677812
transform 1 0 3800 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4216
timestamp 1677677812
transform 1 0 3808 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4217
timestamp 1677677812
transform 1 0 3816 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4218
timestamp 1677677812
transform 1 0 3824 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4219
timestamp 1677677812
transform 1 0 3832 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4220
timestamp 1677677812
transform 1 0 3840 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4227
timestamp 1677677812
transform 1 0 3848 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4228
timestamp 1677677812
transform 1 0 3856 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4229
timestamp 1677677812
transform 1 0 3864 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4230
timestamp 1677677812
transform 1 0 3872 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4231
timestamp 1677677812
transform 1 0 3880 0 -1 2970
box -8 -3 16 105
use AOI22X1  AOI22X1_179
timestamp 1677677812
transform 1 0 3888 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4232
timestamp 1677677812
transform 1 0 3928 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4233
timestamp 1677677812
transform 1 0 3936 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4234
timestamp 1677677812
transform 1 0 3944 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4235
timestamp 1677677812
transform 1 0 3952 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4236
timestamp 1677677812
transform 1 0 3960 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4237
timestamp 1677677812
transform 1 0 3968 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4238
timestamp 1677677812
transform 1 0 3976 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4239
timestamp 1677677812
transform 1 0 3984 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4240
timestamp 1677677812
transform 1 0 3992 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_170
timestamp 1677677812
transform 1 0 4000 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4241
timestamp 1677677812
transform 1 0 4040 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4243
timestamp 1677677812
transform 1 0 4048 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4257
timestamp 1677677812
transform 1 0 4056 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4258
timestamp 1677677812
transform 1 0 4064 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4259
timestamp 1677677812
transform 1 0 4072 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_259
timestamp 1677677812
transform -1 0 4176 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4260
timestamp 1677677812
transform 1 0 4176 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4261
timestamp 1677677812
transform 1 0 4184 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4262
timestamp 1677677812
transform 1 0 4192 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_172
timestamp 1677677812
transform 1 0 4200 0 -1 2970
box -8 -3 46 105
use INVX2  INVX2_290
timestamp 1677677812
transform 1 0 4240 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4263
timestamp 1677677812
transform 1 0 4256 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4265
timestamp 1677677812
transform 1 0 4264 0 -1 2970
box -8 -3 16 105
use M3_M2  M3_M2_3483
timestamp 1677677812
transform 1 0 4284 0 1 2875
box -3 -3 3 3
use FILL  FILL_4266
timestamp 1677677812
transform 1 0 4272 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4267
timestamp 1677677812
transform 1 0 4280 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4268
timestamp 1677677812
transform 1 0 4288 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_173
timestamp 1677677812
transform 1 0 4296 0 -1 2970
box -8 -3 46 105
use FILL  FILL_4273
timestamp 1677677812
transform 1 0 4336 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4274
timestamp 1677677812
transform 1 0 4344 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4275
timestamp 1677677812
transform 1 0 4352 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4276
timestamp 1677677812
transform 1 0 4360 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4286
timestamp 1677677812
transform 1 0 4368 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_292
timestamp 1677677812
transform -1 0 4392 0 -1 2970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_260
timestamp 1677677812
transform 1 0 4392 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4287
timestamp 1677677812
transform 1 0 4488 0 -1 2970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_261
timestamp 1677677812
transform 1 0 4496 0 -1 2970
box -8 -3 104 105
use FILL  FILL_4296
timestamp 1677677812
transform 1 0 4592 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4297
timestamp 1677677812
transform 1 0 4600 0 -1 2970
box -8 -3 16 105
use FILL  FILL_4298
timestamp 1677677812
transform 1 0 4608 0 -1 2970
box -8 -3 16 105
use INVX2  INVX2_293
timestamp 1677677812
transform 1 0 4616 0 -1 2970
box -9 -3 26 105
use FILL  FILL_4299
timestamp 1677677812
transform 1 0 4632 0 -1 2970
box -8 -3 16 105
use OAI22X1  OAI22X1_177
timestamp 1677677812
transform 1 0 4640 0 -1 2970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_262
timestamp 1677677812
transform 1 0 4680 0 -1 2970
box -8 -3 104 105
use INVX2  INVX2_295
timestamp 1677677812
transform 1 0 4776 0 -1 2970
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_37
timestamp 1677677812
transform 1 0 4843 0 1 2870
box -10 -3 10 3
use M3_M2  M3_M2_3491
timestamp 1677677812
transform 1 0 84 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3953
timestamp 1677677812
transform 1 0 108 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3954
timestamp 1677677812
transform 1 0 164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3955
timestamp 1677677812
transform 1 0 204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3956
timestamp 1677677812
transform 1 0 260 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3957
timestamp 1677677812
transform 1 0 268 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4044
timestamp 1677677812
transform 1 0 84 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4045
timestamp 1677677812
transform 1 0 180 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3598
timestamp 1677677812
transform 1 0 180 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3615
timestamp 1677677812
transform 1 0 212 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4046
timestamp 1677677812
transform 1 0 292 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3616
timestamp 1677677812
transform 1 0 292 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3492
timestamp 1677677812
transform 1 0 308 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3526
timestamp 1677677812
transform 1 0 356 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3527
timestamp 1677677812
transform 1 0 396 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3958
timestamp 1677677812
transform 1 0 356 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3959
timestamp 1677677812
transform 1 0 388 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3960
timestamp 1677677812
transform 1 0 396 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4047
timestamp 1677677812
transform 1 0 308 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3617
timestamp 1677677812
transform 1 0 308 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3618
timestamp 1677677812
transform 1 0 348 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4048
timestamp 1677677812
transform 1 0 396 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3507
timestamp 1677677812
transform 1 0 524 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3528
timestamp 1677677812
transform 1 0 492 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3529
timestamp 1677677812
transform 1 0 532 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3961
timestamp 1677677812
transform 1 0 492 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3962
timestamp 1677677812
transform 1 0 524 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3963
timestamp 1677677812
transform 1 0 532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4049
timestamp 1677677812
transform 1 0 444 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3599
timestamp 1677677812
transform 1 0 444 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4050
timestamp 1677677812
transform 1 0 564 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3508
timestamp 1677677812
transform 1 0 572 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3530
timestamp 1677677812
transform 1 0 580 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3964
timestamp 1677677812
transform 1 0 580 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3493
timestamp 1677677812
transform 1 0 628 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3965
timestamp 1677677812
transform 1 0 644 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3565
timestamp 1677677812
transform 1 0 668 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4051
timestamp 1677677812
transform 1 0 668 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3619
timestamp 1677677812
transform 1 0 620 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3509
timestamp 1677677812
transform 1 0 692 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3531
timestamp 1677677812
transform 1 0 692 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4052
timestamp 1677677812
transform 1 0 692 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3966
timestamp 1677677812
transform 1 0 708 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3510
timestamp 1677677812
transform 1 0 724 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4053
timestamp 1677677812
transform 1 0 740 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3600
timestamp 1677677812
transform 1 0 756 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3620
timestamp 1677677812
transform 1 0 756 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3967
timestamp 1677677812
transform 1 0 772 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3968
timestamp 1677677812
transform 1 0 796 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4054
timestamp 1677677812
transform 1 0 804 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3944
timestamp 1677677812
transform 1 0 812 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3532
timestamp 1677677812
transform 1 0 852 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3969
timestamp 1677677812
transform 1 0 836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4055
timestamp 1677677812
transform 1 0 852 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3970
timestamp 1677677812
transform 1 0 868 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3566
timestamp 1677677812
transform 1 0 876 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3533
timestamp 1677677812
transform 1 0 900 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3971
timestamp 1677677812
transform 1 0 908 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4056
timestamp 1677677812
transform 1 0 964 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3503
timestamp 1677677812
transform 1 0 1004 0 1 2845
box -3 -3 3 3
use M3_M2  M3_M2_3511
timestamp 1677677812
transform 1 0 996 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3534
timestamp 1677677812
transform 1 0 1012 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3972
timestamp 1677677812
transform 1 0 996 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3973
timestamp 1677677812
transform 1 0 1012 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4057
timestamp 1677677812
transform 1 0 1004 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3581
timestamp 1677677812
transform 1 0 1012 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3484
timestamp 1677677812
transform 1 0 1052 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3974
timestamp 1677677812
transform 1 0 1044 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4058
timestamp 1677677812
transform 1 0 1100 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3567
timestamp 1677677812
transform 1 0 1132 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4059
timestamp 1677677812
transform 1 0 1132 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3535
timestamp 1677677812
transform 1 0 1148 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3975
timestamp 1677677812
transform 1 0 1148 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3494
timestamp 1677677812
transform 1 0 1212 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3536
timestamp 1677677812
transform 1 0 1196 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3568
timestamp 1677677812
transform 1 0 1172 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_3976
timestamp 1677677812
transform 1 0 1196 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4060
timestamp 1677677812
transform 1 0 1172 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3977
timestamp 1677677812
transform 1 0 1260 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3537
timestamp 1677677812
transform 1 0 1348 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3538
timestamp 1677677812
transform 1 0 1380 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3485
timestamp 1677677812
transform 1 0 1412 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3512
timestamp 1677677812
transform 1 0 1404 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3513
timestamp 1677677812
transform 1 0 1420 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3486
timestamp 1677677812
transform 1 0 1468 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3539
timestamp 1677677812
transform 1 0 1460 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3978
timestamp 1677677812
transform 1 0 1460 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4061
timestamp 1677677812
transform 1 0 1452 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4062
timestamp 1677677812
transform 1 0 1468 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4063
timestamp 1677677812
transform 1 0 1484 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4064
timestamp 1677677812
transform 1 0 1500 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3979
timestamp 1677677812
transform 1 0 1548 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3540
timestamp 1677677812
transform 1 0 1620 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3980
timestamp 1677677812
transform 1 0 1620 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4065
timestamp 1677677812
transform 1 0 1572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3981
timestamp 1677677812
transform 1 0 1660 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3541
timestamp 1677677812
transform 1 0 1676 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4066
timestamp 1677677812
transform 1 0 1684 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3514
timestamp 1677677812
transform 1 0 1708 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3982
timestamp 1677677812
transform 1 0 1708 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3983
timestamp 1677677812
transform 1 0 1724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4067
timestamp 1677677812
transform 1 0 1716 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3487
timestamp 1677677812
transform 1 0 1756 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3488
timestamp 1677677812
transform 1 0 1780 0 1 2865
box -3 -3 3 3
use M3_M2  M3_M2_3495
timestamp 1677677812
transform 1 0 1748 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3496
timestamp 1677677812
transform 1 0 1788 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3497
timestamp 1677677812
transform 1 0 1820 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_4068
timestamp 1677677812
transform 1 0 1740 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3515
timestamp 1677677812
transform 1 0 1820 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3542
timestamp 1677677812
transform 1 0 1804 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3543
timestamp 1677677812
transform 1 0 1844 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3984
timestamp 1677677812
transform 1 0 1804 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3985
timestamp 1677677812
transform 1 0 1836 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3986
timestamp 1677677812
transform 1 0 1844 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4069
timestamp 1677677812
transform 1 0 1756 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3582
timestamp 1677677812
transform 1 0 1780 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3583
timestamp 1677677812
transform 1 0 1804 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3601
timestamp 1677677812
transform 1 0 1780 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3621
timestamp 1677677812
transform 1 0 1756 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3498
timestamp 1677677812
transform 1 0 1892 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_4070
timestamp 1677677812
transform 1 0 1900 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3544
timestamp 1677677812
transform 1 0 2060 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3545
timestamp 1677677812
transform 1 0 2100 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3987
timestamp 1677677812
transform 1 0 1956 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3988
timestamp 1677677812
transform 1 0 1996 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3989
timestamp 1677677812
transform 1 0 2060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3990
timestamp 1677677812
transform 1 0 2092 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3991
timestamp 1677677812
transform 1 0 2100 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4071
timestamp 1677677812
transform 1 0 1916 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3622
timestamp 1677677812
transform 1 0 1916 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4072
timestamp 1677677812
transform 1 0 2012 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4073
timestamp 1677677812
transform 1 0 2100 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3602
timestamp 1677677812
transform 1 0 2108 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3623
timestamp 1677677812
transform 1 0 2012 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3624
timestamp 1677677812
transform 1 0 2100 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4074
timestamp 1677677812
transform 1 0 2124 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_3992
timestamp 1677677812
transform 1 0 2140 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3625
timestamp 1677677812
transform 1 0 2132 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3993
timestamp 1677677812
transform 1 0 2172 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3994
timestamp 1677677812
transform 1 0 2188 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4075
timestamp 1677677812
transform 1 0 2180 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3626
timestamp 1677677812
transform 1 0 2188 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_3995
timestamp 1677677812
transform 1 0 2284 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4076
timestamp 1677677812
transform 1 0 2276 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3546
timestamp 1677677812
transform 1 0 2316 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3996
timestamp 1677677812
transform 1 0 2364 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3997
timestamp 1677677812
transform 1 0 2380 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_3998
timestamp 1677677812
transform 1 0 2396 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3584
timestamp 1677677812
transform 1 0 2364 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4077
timestamp 1677677812
transform 1 0 2372 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3569
timestamp 1677677812
transform 1 0 2404 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4078
timestamp 1677677812
transform 1 0 2404 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3547
timestamp 1677677812
transform 1 0 2420 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4079
timestamp 1677677812
transform 1 0 2420 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3548
timestamp 1677677812
transform 1 0 2436 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3570
timestamp 1677677812
transform 1 0 2444 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3549
timestamp 1677677812
transform 1 0 2484 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3999
timestamp 1677677812
transform 1 0 2468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4000
timestamp 1677677812
transform 1 0 2484 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3571
timestamp 1677677812
transform 1 0 2492 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4001
timestamp 1677677812
transform 1 0 2500 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4080
timestamp 1677677812
transform 1 0 2476 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4081
timestamp 1677677812
transform 1 0 2492 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3627
timestamp 1677677812
transform 1 0 2484 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3585
timestamp 1677677812
transform 1 0 2500 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4082
timestamp 1677677812
transform 1 0 2540 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4002
timestamp 1677677812
transform 1 0 2564 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3572
timestamp 1677677812
transform 1 0 2572 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4083
timestamp 1677677812
transform 1 0 2556 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4084
timestamp 1677677812
transform 1 0 2572 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4085
timestamp 1677677812
transform 1 0 2580 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3628
timestamp 1677677812
transform 1 0 2548 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3629
timestamp 1677677812
transform 1 0 2580 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4003
timestamp 1677677812
transform 1 0 2596 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4004
timestamp 1677677812
transform 1 0 2612 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3550
timestamp 1677677812
transform 1 0 2644 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4005
timestamp 1677677812
transform 1 0 2644 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3551
timestamp 1677677812
transform 1 0 2684 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4006
timestamp 1677677812
transform 1 0 2684 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3573
timestamp 1677677812
transform 1 0 2732 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4007
timestamp 1677677812
transform 1 0 2740 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4086
timestamp 1677677812
transform 1 0 2660 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4116
timestamp 1677677812
transform 1 0 2748 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3630
timestamp 1677677812
transform 1 0 2748 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3574
timestamp 1677677812
transform 1 0 2788 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4087
timestamp 1677677812
transform 1 0 2780 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4088
timestamp 1677677812
transform 1 0 2788 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4008
timestamp 1677677812
transform 1 0 2812 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3586
timestamp 1677677812
transform 1 0 2812 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3499
timestamp 1677677812
transform 1 0 2836 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_4009
timestamp 1677677812
transform 1 0 2828 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4089
timestamp 1677677812
transform 1 0 2844 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3489
timestamp 1677677812
transform 1 0 2860 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_3945
timestamp 1677677812
transform 1 0 2860 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3575
timestamp 1677677812
transform 1 0 2860 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4117
timestamp 1677677812
transform 1 0 2852 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3576
timestamp 1677677812
transform 1 0 2892 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4090
timestamp 1677677812
transform 1 0 2884 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4091
timestamp 1677677812
transform 1 0 2892 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3552
timestamp 1677677812
transform 1 0 2924 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3516
timestamp 1677677812
transform 1 0 2940 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3946
timestamp 1677677812
transform 1 0 2932 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4010
timestamp 1677677812
transform 1 0 2924 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3587
timestamp 1677677812
transform 1 0 2916 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3517
timestamp 1677677812
transform 1 0 2964 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3553
timestamp 1677677812
transform 1 0 2956 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4011
timestamp 1677677812
transform 1 0 2948 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3588
timestamp 1677677812
transform 1 0 2948 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3589
timestamp 1677677812
transform 1 0 2996 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4092
timestamp 1677677812
transform 1 0 3012 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4118
timestamp 1677677812
transform 1 0 3004 0 1 2795
box -2 -2 2 2
use M3_M2  M3_M2_3554
timestamp 1677677812
transform 1 0 3028 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4012
timestamp 1677677812
transform 1 0 3028 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3555
timestamp 1677677812
transform 1 0 3068 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4013
timestamp 1677677812
transform 1 0 3044 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3577
timestamp 1677677812
transform 1 0 3060 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4014
timestamp 1677677812
transform 1 0 3068 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4093
timestamp 1677677812
transform 1 0 3052 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4094
timestamp 1677677812
transform 1 0 3076 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3518
timestamp 1677677812
transform 1 0 3204 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4015
timestamp 1677677812
transform 1 0 3164 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4095
timestamp 1677677812
transform 1 0 3116 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3603
timestamp 1677677812
transform 1 0 3164 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3556
timestamp 1677677812
transform 1 0 3212 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4016
timestamp 1677677812
transform 1 0 3212 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4096
timestamp 1677677812
transform 1 0 3220 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3519
timestamp 1677677812
transform 1 0 3252 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3557
timestamp 1677677812
transform 1 0 3252 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4017
timestamp 1677677812
transform 1 0 3252 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4018
timestamp 1677677812
transform 1 0 3268 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3558
timestamp 1677677812
transform 1 0 3332 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4019
timestamp 1677677812
transform 1 0 3340 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4097
timestamp 1677677812
transform 1 0 3244 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4098
timestamp 1677677812
transform 1 0 3260 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4099
timestamp 1677677812
transform 1 0 3276 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4100
timestamp 1677677812
transform 1 0 3292 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3604
timestamp 1677677812
transform 1 0 3260 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3590
timestamp 1677677812
transform 1 0 3340 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3631
timestamp 1677677812
transform 1 0 3284 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3632
timestamp 1677677812
transform 1 0 3324 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3605
timestamp 1677677812
transform 1 0 3380 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4020
timestamp 1677677812
transform 1 0 3404 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4021
timestamp 1677677812
transform 1 0 3428 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3606
timestamp 1677677812
transform 1 0 3428 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3578
timestamp 1677677812
transform 1 0 3444 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4101
timestamp 1677677812
transform 1 0 3500 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3520
timestamp 1677677812
transform 1 0 3564 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4022
timestamp 1677677812
transform 1 0 3564 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4023
timestamp 1677677812
transform 1 0 3580 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4024
timestamp 1677677812
transform 1 0 3596 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3607
timestamp 1677677812
transform 1 0 3604 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_3947
timestamp 1677677812
transform 1 0 3628 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3591
timestamp 1677677812
transform 1 0 3628 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3559
timestamp 1677677812
transform 1 0 3644 0 1 2825
box -3 -3 3 3
use M3_M2  M3_M2_3521
timestamp 1677677812
transform 1 0 3660 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4102
timestamp 1677677812
transform 1 0 3668 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3504
timestamp 1677677812
transform 1 0 3716 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3941
timestamp 1677677812
transform 1 0 3716 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3948
timestamp 1677677812
transform 1 0 3700 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3560
timestamp 1677677812
transform 1 0 3708 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_3949
timestamp 1677677812
transform 1 0 3732 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3608
timestamp 1677677812
transform 1 0 3764 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3500
timestamp 1677677812
transform 1 0 3796 0 1 2855
box -3 -3 3 3
use M2_M1  M2_M1_3942
timestamp 1677677812
transform 1 0 3796 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_4025
timestamp 1677677812
transform 1 0 3804 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3579
timestamp 1677677812
transform 1 0 3812 0 1 2815
box -3 -3 3 3
use M3_M2  M3_M2_3609
timestamp 1677677812
transform 1 0 3844 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3505
timestamp 1677677812
transform 1 0 3868 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3950
timestamp 1677677812
transform 1 0 3908 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3592
timestamp 1677677812
transform 1 0 3964 0 1 2805
box -3 -3 3 3
use M2_M1  M2_M1_4026
timestamp 1677677812
transform 1 0 4012 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4027
timestamp 1677677812
transform 1 0 4060 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4103
timestamp 1677677812
transform 1 0 3980 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3593
timestamp 1677677812
transform 1 0 4012 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3610
timestamp 1677677812
transform 1 0 4044 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4104
timestamp 1677677812
transform 1 0 4084 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3594
timestamp 1677677812
transform 1 0 4092 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3490
timestamp 1677677812
transform 1 0 4108 0 1 2865
box -3 -3 3 3
use M2_M1  M2_M1_4028
timestamp 1677677812
transform 1 0 4132 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3595
timestamp 1677677812
transform 1 0 4132 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3561
timestamp 1677677812
transform 1 0 4156 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4029
timestamp 1677677812
transform 1 0 4204 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4030
timestamp 1677677812
transform 1 0 4236 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4105
timestamp 1677677812
transform 1 0 4156 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3506
timestamp 1677677812
transform 1 0 4252 0 1 2845
box -3 -3 3 3
use M2_M1  M2_M1_3943
timestamp 1677677812
transform 1 0 4284 0 1 2835
box -2 -2 2 2
use M2_M1  M2_M1_3951
timestamp 1677677812
transform 1 0 4276 0 1 2825
box -2 -2 2 2
use M2_M1  M2_M1_4031
timestamp 1677677812
transform 1 0 4292 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3596
timestamp 1677677812
transform 1 0 4284 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3522
timestamp 1677677812
transform 1 0 4316 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_3952
timestamp 1677677812
transform 1 0 4316 0 1 2825
box -2 -2 2 2
use M3_M2  M3_M2_3501
timestamp 1677677812
transform 1 0 4348 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3523
timestamp 1677677812
transform 1 0 4372 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3524
timestamp 1677677812
transform 1 0 4388 0 1 2835
box -3 -3 3 3
use M3_M2  M3_M2_3562
timestamp 1677677812
transform 1 0 4348 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4032
timestamp 1677677812
transform 1 0 4372 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4106
timestamp 1677677812
transform 1 0 4348 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3611
timestamp 1677677812
transform 1 0 4420 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4033
timestamp 1677677812
transform 1 0 4436 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4034
timestamp 1677677812
transform 1 0 4444 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4035
timestamp 1677677812
transform 1 0 4452 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4036
timestamp 1677677812
transform 1 0 4468 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4119
timestamp 1677677812
transform 1 0 4436 0 1 2785
box -2 -2 2 2
use M2_M1  M2_M1_4107
timestamp 1677677812
transform 1 0 4460 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4108
timestamp 1677677812
transform 1 0 4476 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4109
timestamp 1677677812
transform 1 0 4484 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3612
timestamp 1677677812
transform 1 0 4476 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3633
timestamp 1677677812
transform 1 0 4452 0 1 2785
box -3 -3 3 3
use M2_M1  M2_M1_4037
timestamp 1677677812
transform 1 0 4492 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3502
timestamp 1677677812
transform 1 0 4508 0 1 2855
box -3 -3 3 3
use M3_M2  M3_M2_3525
timestamp 1677677812
transform 1 0 4556 0 1 2835
box -3 -3 3 3
use M2_M1  M2_M1_4038
timestamp 1677677812
transform 1 0 4532 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4039
timestamp 1677677812
transform 1 0 4556 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4110
timestamp 1677677812
transform 1 0 4524 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3597
timestamp 1677677812
transform 1 0 4532 0 1 2805
box -3 -3 3 3
use M3_M2  M3_M2_3580
timestamp 1677677812
transform 1 0 4564 0 1 2815
box -3 -3 3 3
use M2_M1  M2_M1_4040
timestamp 1677677812
transform 1 0 4572 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4111
timestamp 1677677812
transform 1 0 4540 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4112
timestamp 1677677812
transform 1 0 4556 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4113
timestamp 1677677812
transform 1 0 4564 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3613
timestamp 1677677812
transform 1 0 4548 0 1 2795
box -3 -3 3 3
use M3_M2  M3_M2_3634
timestamp 1677677812
transform 1 0 4548 0 1 2785
box -3 -3 3 3
use M3_M2  M3_M2_3614
timestamp 1677677812
transform 1 0 4588 0 1 2795
box -3 -3 3 3
use M2_M1  M2_M1_4041
timestamp 1677677812
transform 1 0 4620 0 1 2815
box -2 -2 2 2
use M3_M2  M3_M2_3563
timestamp 1677677812
transform 1 0 4660 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4114
timestamp 1677677812
transform 1 0 4668 0 1 2805
box -2 -2 2 2
use M3_M2  M3_M2_3564
timestamp 1677677812
transform 1 0 4724 0 1 2825
box -3 -3 3 3
use M2_M1  M2_M1_4042
timestamp 1677677812
transform 1 0 4724 0 1 2815
box -2 -2 2 2
use M2_M1  M2_M1_4115
timestamp 1677677812
transform 1 0 4700 0 1 2805
box -2 -2 2 2
use M2_M1  M2_M1_4043
timestamp 1677677812
transform 1 0 4804 0 1 2815
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_38
timestamp 1677677812
transform 1 0 48 0 1 2770
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_263
timestamp 1677677812
transform 1 0 72 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_264
timestamp 1677677812
transform 1 0 168 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_296
timestamp 1677677812
transform -1 0 280 0 1 2770
box -9 -3 26 105
use FILL  FILL_4312
timestamp 1677677812
transform 1 0 280 0 1 2770
box -8 -3 16 105
use FILL  FILL_4313
timestamp 1677677812
transform 1 0 288 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3635
timestamp 1677677812
transform 1 0 388 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_265
timestamp 1677677812
transform 1 0 296 0 1 2770
box -8 -3 104 105
use M3_M2  M3_M2_3636
timestamp 1677677812
transform 1 0 404 0 1 2775
box -3 -3 3 3
use FILL  FILL_4314
timestamp 1677677812
transform 1 0 392 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_297
timestamp 1677677812
transform 1 0 400 0 1 2770
box -9 -3 26 105
use FILL  FILL_4315
timestamp 1677677812
transform 1 0 416 0 1 2770
box -8 -3 16 105
use FILL  FILL_4334
timestamp 1677677812
transform 1 0 424 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_266
timestamp 1677677812
transform 1 0 432 0 1 2770
box -8 -3 104 105
use FILL  FILL_4336
timestamp 1677677812
transform 1 0 528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4338
timestamp 1677677812
transform 1 0 536 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_301
timestamp 1677677812
transform -1 0 560 0 1 2770
box -9 -3 26 105
use FILL  FILL_4339
timestamp 1677677812
transform 1 0 560 0 1 2770
box -8 -3 16 105
use FILL  FILL_4344
timestamp 1677677812
transform 1 0 568 0 1 2770
box -8 -3 16 105
use FILL  FILL_4346
timestamp 1677677812
transform 1 0 576 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_268
timestamp 1677677812
transform -1 0 680 0 1 2770
box -8 -3 104 105
use FILL  FILL_4347
timestamp 1677677812
transform 1 0 680 0 1 2770
box -8 -3 16 105
use FILL  FILL_4357
timestamp 1677677812
transform 1 0 688 0 1 2770
box -8 -3 16 105
use FILL  FILL_4358
timestamp 1677677812
transform 1 0 696 0 1 2770
box -8 -3 16 105
use FILL  FILL_4359
timestamp 1677677812
transform 1 0 704 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_93
timestamp 1677677812
transform 1 0 712 0 1 2770
box -8 -3 34 105
use FILL  FILL_4360
timestamp 1677677812
transform 1 0 744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4367
timestamp 1677677812
transform 1 0 752 0 1 2770
box -8 -3 16 105
use FILL  FILL_4368
timestamp 1677677812
transform 1 0 760 0 1 2770
box -8 -3 16 105
use FILL  FILL_4369
timestamp 1677677812
transform 1 0 768 0 1 2770
box -8 -3 16 105
use FILL  FILL_4370
timestamp 1677677812
transform 1 0 776 0 1 2770
box -8 -3 16 105
use FILL  FILL_4371
timestamp 1677677812
transform 1 0 784 0 1 2770
box -8 -3 16 105
use FILL  FILL_4372
timestamp 1677677812
transform 1 0 792 0 1 2770
box -8 -3 16 105
use FILL  FILL_4373
timestamp 1677677812
transform 1 0 800 0 1 2770
box -8 -3 16 105
use FILL  FILL_4376
timestamp 1677677812
transform 1 0 808 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3637
timestamp 1677677812
transform 1 0 852 0 1 2775
box -3 -3 3 3
use AOI22X1  AOI22X1_187
timestamp 1677677812
transform -1 0 856 0 1 2770
box -8 -3 46 105
use FILL  FILL_4377
timestamp 1677677812
transform 1 0 856 0 1 2770
box -8 -3 16 105
use FILL  FILL_4385
timestamp 1677677812
transform 1 0 864 0 1 2770
box -8 -3 16 105
use FILL  FILL_4386
timestamp 1677677812
transform 1 0 872 0 1 2770
box -8 -3 16 105
use FILL  FILL_4387
timestamp 1677677812
transform 1 0 880 0 1 2770
box -8 -3 16 105
use FILL  FILL_4388
timestamp 1677677812
transform 1 0 888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4389
timestamp 1677677812
transform 1 0 896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4390
timestamp 1677677812
transform 1 0 904 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_303
timestamp 1677677812
transform -1 0 928 0 1 2770
box -9 -3 26 105
use FILL  FILL_4391
timestamp 1677677812
transform 1 0 928 0 1 2770
box -8 -3 16 105
use FILL  FILL_4392
timestamp 1677677812
transform 1 0 936 0 1 2770
box -8 -3 16 105
use FILL  FILL_4393
timestamp 1677677812
transform 1 0 944 0 1 2770
box -8 -3 16 105
use FILL  FILL_4394
timestamp 1677677812
transform 1 0 952 0 1 2770
box -8 -3 16 105
use FILL  FILL_4395
timestamp 1677677812
transform 1 0 960 0 1 2770
box -8 -3 16 105
use FILL  FILL_4397
timestamp 1677677812
transform 1 0 968 0 1 2770
box -8 -3 16 105
use FILL  FILL_4399
timestamp 1677677812
transform 1 0 976 0 1 2770
box -8 -3 16 105
use FILL  FILL_4401
timestamp 1677677812
transform 1 0 984 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_188
timestamp 1677677812
transform 1 0 992 0 1 2770
box -8 -3 46 105
use FILL  FILL_4403
timestamp 1677677812
transform 1 0 1032 0 1 2770
box -8 -3 16 105
use FILL  FILL_4407
timestamp 1677677812
transform 1 0 1040 0 1 2770
box -8 -3 16 105
use FILL  FILL_4409
timestamp 1677677812
transform 1 0 1048 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3638
timestamp 1677677812
transform 1 0 1068 0 1 2775
box -3 -3 3 3
use FILL  FILL_4411
timestamp 1677677812
transform 1 0 1056 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3639
timestamp 1677677812
transform 1 0 1084 0 1 2775
box -3 -3 3 3
use FILL  FILL_4412
timestamp 1677677812
transform 1 0 1064 0 1 2770
box -8 -3 16 105
use FILL  FILL_4413
timestamp 1677677812
transform 1 0 1072 0 1 2770
box -8 -3 16 105
use FILL  FILL_4414
timestamp 1677677812
transform 1 0 1080 0 1 2770
box -8 -3 16 105
use FILL  FILL_4415
timestamp 1677677812
transform 1 0 1088 0 1 2770
box -8 -3 16 105
use FILL  FILL_4416
timestamp 1677677812
transform 1 0 1096 0 1 2770
box -8 -3 16 105
use FILL  FILL_4418
timestamp 1677677812
transform 1 0 1104 0 1 2770
box -8 -3 16 105
use FILL  FILL_4420
timestamp 1677677812
transform 1 0 1112 0 1 2770
box -8 -3 16 105
use FILL  FILL_4422
timestamp 1677677812
transform 1 0 1120 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3640
timestamp 1677677812
transform 1 0 1140 0 1 2775
box -3 -3 3 3
use INVX2  INVX2_304
timestamp 1677677812
transform 1 0 1128 0 1 2770
box -9 -3 26 105
use FILL  FILL_4424
timestamp 1677677812
transform 1 0 1144 0 1 2770
box -8 -3 16 105
use FILL  FILL_4425
timestamp 1677677812
transform 1 0 1152 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3641
timestamp 1677677812
transform 1 0 1172 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3642
timestamp 1677677812
transform 1 0 1188 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3643
timestamp 1677677812
transform 1 0 1220 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_270
timestamp 1677677812
transform 1 0 1160 0 1 2770
box -8 -3 104 105
use FILL  FILL_4426
timestamp 1677677812
transform 1 0 1256 0 1 2770
box -8 -3 16 105
use FILL  FILL_4427
timestamp 1677677812
transform 1 0 1264 0 1 2770
box -8 -3 16 105
use FILL  FILL_4428
timestamp 1677677812
transform 1 0 1272 0 1 2770
box -8 -3 16 105
use FILL  FILL_4429
timestamp 1677677812
transform 1 0 1280 0 1 2770
box -8 -3 16 105
use FILL  FILL_4430
timestamp 1677677812
transform 1 0 1288 0 1 2770
box -8 -3 16 105
use FILL  FILL_4431
timestamp 1677677812
transform 1 0 1296 0 1 2770
box -8 -3 16 105
use FILL  FILL_4432
timestamp 1677677812
transform 1 0 1304 0 1 2770
box -8 -3 16 105
use FILL  FILL_4440
timestamp 1677677812
transform 1 0 1312 0 1 2770
box -8 -3 16 105
use FILL  FILL_4442
timestamp 1677677812
transform 1 0 1320 0 1 2770
box -8 -3 16 105
use FILL  FILL_4443
timestamp 1677677812
transform 1 0 1328 0 1 2770
box -8 -3 16 105
use FILL  FILL_4444
timestamp 1677677812
transform 1 0 1336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4446
timestamp 1677677812
transform 1 0 1344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4448
timestamp 1677677812
transform 1 0 1352 0 1 2770
box -8 -3 16 105
use FILL  FILL_4450
timestamp 1677677812
transform 1 0 1360 0 1 2770
box -8 -3 16 105
use FILL  FILL_4452
timestamp 1677677812
transform 1 0 1368 0 1 2770
box -8 -3 16 105
use FILL  FILL_4453
timestamp 1677677812
transform 1 0 1376 0 1 2770
box -8 -3 16 105
use FILL  FILL_4454
timestamp 1677677812
transform 1 0 1384 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3644
timestamp 1677677812
transform 1 0 1404 0 1 2775
box -3 -3 3 3
use FILL  FILL_4455
timestamp 1677677812
transform 1 0 1392 0 1 2770
box -8 -3 16 105
use FILL  FILL_4456
timestamp 1677677812
transform 1 0 1400 0 1 2770
box -8 -3 16 105
use FILL  FILL_4457
timestamp 1677677812
transform 1 0 1408 0 1 2770
box -8 -3 16 105
use FILL  FILL_4460
timestamp 1677677812
transform 1 0 1416 0 1 2770
box -8 -3 16 105
use FILL  FILL_4462
timestamp 1677677812
transform 1 0 1424 0 1 2770
box -8 -3 16 105
use FILL  FILL_4464
timestamp 1677677812
transform 1 0 1432 0 1 2770
box -8 -3 16 105
use FILL  FILL_4466
timestamp 1677677812
transform 1 0 1440 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3645
timestamp 1677677812
transform 1 0 1468 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_180
timestamp 1677677812
transform -1 0 1488 0 1 2770
box -8 -3 46 105
use FILL  FILL_4467
timestamp 1677677812
transform 1 0 1488 0 1 2770
box -8 -3 16 105
use FILL  FILL_4468
timestamp 1677677812
transform 1 0 1496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4469
timestamp 1677677812
transform 1 0 1504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4470
timestamp 1677677812
transform 1 0 1512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4476
timestamp 1677677812
transform 1 0 1520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4478
timestamp 1677677812
transform 1 0 1528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4480
timestamp 1677677812
transform 1 0 1536 0 1 2770
box -8 -3 16 105
use FILL  FILL_4482
timestamp 1677677812
transform 1 0 1544 0 1 2770
box -8 -3 16 105
use FILL  FILL_4484
timestamp 1677677812
transform 1 0 1552 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3646
timestamp 1677677812
transform 1 0 1628 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_272
timestamp 1677677812
transform 1 0 1560 0 1 2770
box -8 -3 104 105
use FILL  FILL_4486
timestamp 1677677812
transform 1 0 1656 0 1 2770
box -8 -3 16 105
use FILL  FILL_4487
timestamp 1677677812
transform 1 0 1664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4488
timestamp 1677677812
transform 1 0 1672 0 1 2770
box -8 -3 16 105
use FILL  FILL_4489
timestamp 1677677812
transform 1 0 1680 0 1 2770
box -8 -3 16 105
use FILL  FILL_4490
timestamp 1677677812
transform 1 0 1688 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_182
timestamp 1677677812
transform -1 0 1736 0 1 2770
box -8 -3 46 105
use FILL  FILL_4491
timestamp 1677677812
transform 1 0 1736 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_273
timestamp 1677677812
transform 1 0 1744 0 1 2770
box -8 -3 104 105
use FILL  FILL_4492
timestamp 1677677812
transform 1 0 1840 0 1 2770
box -8 -3 16 105
use FILL  FILL_4493
timestamp 1677677812
transform 1 0 1848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4494
timestamp 1677677812
transform 1 0 1856 0 1 2770
box -8 -3 16 105
use FILL  FILL_4495
timestamp 1677677812
transform 1 0 1864 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_306
timestamp 1677677812
transform -1 0 1888 0 1 2770
box -9 -3 26 105
use FILL  FILL_4496
timestamp 1677677812
transform 1 0 1888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4497
timestamp 1677677812
transform 1 0 1896 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_274
timestamp 1677677812
transform 1 0 1904 0 1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_275
timestamp 1677677812
transform 1 0 2000 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_307
timestamp 1677677812
transform 1 0 2096 0 1 2770
box -9 -3 26 105
use FILL  FILL_4498
timestamp 1677677812
transform 1 0 2112 0 1 2770
box -8 -3 16 105
use FILL  FILL_4499
timestamp 1677677812
transform 1 0 2120 0 1 2770
box -8 -3 16 105
use FILL  FILL_4500
timestamp 1677677812
transform 1 0 2128 0 1 2770
box -8 -3 16 105
use FILL  FILL_4535
timestamp 1677677812
transform 1 0 2136 0 1 2770
box -8 -3 16 105
use FILL  FILL_4537
timestamp 1677677812
transform 1 0 2144 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_191
timestamp 1677677812
transform -1 0 2192 0 1 2770
box -8 -3 46 105
use FILL  FILL_4538
timestamp 1677677812
transform 1 0 2192 0 1 2770
box -8 -3 16 105
use FILL  FILL_4544
timestamp 1677677812
transform 1 0 2200 0 1 2770
box -8 -3 16 105
use FILL  FILL_4546
timestamp 1677677812
transform 1 0 2208 0 1 2770
box -8 -3 16 105
use FILL  FILL_4548
timestamp 1677677812
transform 1 0 2216 0 1 2770
box -8 -3 16 105
use FILL  FILL_4550
timestamp 1677677812
transform 1 0 2224 0 1 2770
box -8 -3 16 105
use FILL  FILL_4552
timestamp 1677677812
transform 1 0 2232 0 1 2770
box -8 -3 16 105
use FILL  FILL_4553
timestamp 1677677812
transform 1 0 2240 0 1 2770
box -8 -3 16 105
use FILL  FILL_4554
timestamp 1677677812
transform 1 0 2248 0 1 2770
box -8 -3 16 105
use FILL  FILL_4556
timestamp 1677677812
transform 1 0 2256 0 1 2770
box -8 -3 16 105
use FILL  FILL_4558
timestamp 1677677812
transform 1 0 2264 0 1 2770
box -8 -3 16 105
use FILL  FILL_4560
timestamp 1677677812
transform 1 0 2272 0 1 2770
box -8 -3 16 105
use FILL  FILL_4562
timestamp 1677677812
transform 1 0 2280 0 1 2770
box -8 -3 16 105
use FILL  FILL_4564
timestamp 1677677812
transform 1 0 2288 0 1 2770
box -8 -3 16 105
use FILL  FILL_4565
timestamp 1677677812
transform 1 0 2296 0 1 2770
box -8 -3 16 105
use FILL  FILL_4566
timestamp 1677677812
transform 1 0 2304 0 1 2770
box -8 -3 16 105
use FILL  FILL_4567
timestamp 1677677812
transform 1 0 2312 0 1 2770
box -8 -3 16 105
use FILL  FILL_4568
timestamp 1677677812
transform 1 0 2320 0 1 2770
box -8 -3 16 105
use FILL  FILL_4569
timestamp 1677677812
transform 1 0 2328 0 1 2770
box -8 -3 16 105
use FILL  FILL_4571
timestamp 1677677812
transform 1 0 2336 0 1 2770
box -8 -3 16 105
use FILL  FILL_4573
timestamp 1677677812
transform 1 0 2344 0 1 2770
box -8 -3 16 105
use FILL  FILL_4575
timestamp 1677677812
transform 1 0 2352 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_193
timestamp 1677677812
transform 1 0 2360 0 1 2770
box -8 -3 46 105
use FILL  FILL_4577
timestamp 1677677812
transform 1 0 2400 0 1 2770
box -8 -3 16 105
use FILL  FILL_4578
timestamp 1677677812
transform 1 0 2408 0 1 2770
box -8 -3 16 105
use FILL  FILL_4579
timestamp 1677677812
transform 1 0 2416 0 1 2770
box -8 -3 16 105
use FILL  FILL_4580
timestamp 1677677812
transform 1 0 2424 0 1 2770
box -8 -3 16 105
use FILL  FILL_4585
timestamp 1677677812
transform 1 0 2432 0 1 2770
box -8 -3 16 105
use FILL  FILL_4587
timestamp 1677677812
transform 1 0 2440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4589
timestamp 1677677812
transform 1 0 2448 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_184
timestamp 1677677812
transform -1 0 2496 0 1 2770
box -8 -3 46 105
use FILL  FILL_4590
timestamp 1677677812
transform 1 0 2496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4596
timestamp 1677677812
transform 1 0 2504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4598
timestamp 1677677812
transform 1 0 2512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4600
timestamp 1677677812
transform 1 0 2520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4602
timestamp 1677677812
transform 1 0 2528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4603
timestamp 1677677812
transform 1 0 2536 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_195
timestamp 1677677812
transform 1 0 2544 0 1 2770
box -8 -3 46 105
use FILL  FILL_4604
timestamp 1677677812
transform 1 0 2584 0 1 2770
box -8 -3 16 105
use FILL  FILL_4608
timestamp 1677677812
transform 1 0 2592 0 1 2770
box -8 -3 16 105
use FILL  FILL_4610
timestamp 1677677812
transform 1 0 2600 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_313
timestamp 1677677812
transform 1 0 2608 0 1 2770
box -9 -3 26 105
use FILL  FILL_4612
timestamp 1677677812
transform 1 0 2624 0 1 2770
box -8 -3 16 105
use FILL  FILL_4614
timestamp 1677677812
transform 1 0 2632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4616
timestamp 1677677812
transform 1 0 2640 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_278
timestamp 1677677812
transform 1 0 2648 0 1 2770
box -8 -3 104 105
use FILL  FILL_4618
timestamp 1677677812
transform 1 0 2744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4619
timestamp 1677677812
transform 1 0 2752 0 1 2770
box -8 -3 16 105
use FILL  FILL_4620
timestamp 1677677812
transform 1 0 2760 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_47
timestamp 1677677812
transform 1 0 2768 0 1 2770
box -8 -3 32 105
use FILL  FILL_4621
timestamp 1677677812
transform 1 0 2792 0 1 2770
box -8 -3 16 105
use FILL  FILL_4622
timestamp 1677677812
transform 1 0 2800 0 1 2770
box -8 -3 16 105
use FILL  FILL_4623
timestamp 1677677812
transform 1 0 2808 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_96
timestamp 1677677812
transform 1 0 2816 0 1 2770
box -8 -3 34 105
use FILL  FILL_4624
timestamp 1677677812
transform 1 0 2848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4627
timestamp 1677677812
transform 1 0 2856 0 1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_48
timestamp 1677677812
transform 1 0 2864 0 1 2770
box -8 -3 32 105
use FILL  FILL_4629
timestamp 1677677812
transform 1 0 2888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4630
timestamp 1677677812
transform 1 0 2896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4631
timestamp 1677677812
transform 1 0 2904 0 1 2770
box -8 -3 16 105
use FILL  FILL_4632
timestamp 1677677812
transform 1 0 2912 0 1 2770
box -8 -3 16 105
use FILL  FILL_4633
timestamp 1677677812
transform 1 0 2920 0 1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_97
timestamp 1677677812
transform -1 0 2960 0 1 2770
box -8 -3 34 105
use FILL  FILL_4634
timestamp 1677677812
transform 1 0 2960 0 1 2770
box -8 -3 16 105
use FILL  FILL_4644
timestamp 1677677812
transform 1 0 2968 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_315
timestamp 1677677812
transform -1 0 2992 0 1 2770
box -9 -3 26 105
use FILL  FILL_4645
timestamp 1677677812
transform 1 0 2992 0 1 2770
box -8 -3 16 105
use FILL  FILL_4646
timestamp 1677677812
transform 1 0 3000 0 1 2770
box -8 -3 16 105
use FILL  FILL_4647
timestamp 1677677812
transform 1 0 3008 0 1 2770
box -8 -3 16 105
use FILL  FILL_4650
timestamp 1677677812
transform 1 0 3016 0 1 2770
box -8 -3 16 105
use FILL  FILL_4652
timestamp 1677677812
transform 1 0 3024 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3647
timestamp 1677677812
transform 1 0 3060 0 1 2775
box -3 -3 3 3
use OAI22X1  OAI22X1_185
timestamp 1677677812
transform -1 0 3072 0 1 2770
box -8 -3 46 105
use FILL  FILL_4653
timestamp 1677677812
transform 1 0 3072 0 1 2770
box -8 -3 16 105
use FILL  FILL_4654
timestamp 1677677812
transform 1 0 3080 0 1 2770
box -8 -3 16 105
use FILL  FILL_4655
timestamp 1677677812
transform 1 0 3088 0 1 2770
box -8 -3 16 105
use FILL  FILL_4656
timestamp 1677677812
transform 1 0 3096 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_281
timestamp 1677677812
transform 1 0 3104 0 1 2770
box -8 -3 104 105
use INVX2  INVX2_316
timestamp 1677677812
transform 1 0 3200 0 1 2770
box -9 -3 26 105
use FILL  FILL_4657
timestamp 1677677812
transform 1 0 3216 0 1 2770
box -8 -3 16 105
use FILL  FILL_4658
timestamp 1677677812
transform 1 0 3224 0 1 2770
box -8 -3 16 105
use FILL  FILL_4659
timestamp 1677677812
transform 1 0 3232 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_186
timestamp 1677677812
transform -1 0 3280 0 1 2770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_282
timestamp 1677677812
transform 1 0 3280 0 1 2770
box -8 -3 104 105
use FILL  FILL_4660
timestamp 1677677812
transform 1 0 3376 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_319
timestamp 1677677812
transform 1 0 3384 0 1 2770
box -9 -3 26 105
use FILL  FILL_4685
timestamp 1677677812
transform 1 0 3400 0 1 2770
box -8 -3 16 105
use FILL  FILL_4689
timestamp 1677677812
transform 1 0 3408 0 1 2770
box -8 -3 16 105
use FILL  FILL_4691
timestamp 1677677812
transform 1 0 3416 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3648
timestamp 1677677812
transform 1 0 3436 0 1 2775
box -3 -3 3 3
use FILL  FILL_4693
timestamp 1677677812
transform 1 0 3424 0 1 2770
box -8 -3 16 105
use FILL  FILL_4695
timestamp 1677677812
transform 1 0 3432 0 1 2770
box -8 -3 16 105
use FILL  FILL_4697
timestamp 1677677812
transform 1 0 3440 0 1 2770
box -8 -3 16 105
use FILL  FILL_4699
timestamp 1677677812
transform 1 0 3448 0 1 2770
box -8 -3 16 105
use FILL  FILL_4701
timestamp 1677677812
transform 1 0 3456 0 1 2770
box -8 -3 16 105
use FILL  FILL_4703
timestamp 1677677812
transform 1 0 3464 0 1 2770
box -8 -3 16 105
use FILL  FILL_4704
timestamp 1677677812
transform 1 0 3472 0 1 2770
box -8 -3 16 105
use FILL  FILL_4705
timestamp 1677677812
transform 1 0 3480 0 1 2770
box -8 -3 16 105
use FILL  FILL_4706
timestamp 1677677812
transform 1 0 3488 0 1 2770
box -8 -3 16 105
use FILL  FILL_4707
timestamp 1677677812
transform 1 0 3496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4708
timestamp 1677677812
transform 1 0 3504 0 1 2770
box -8 -3 16 105
use FILL  FILL_4709
timestamp 1677677812
transform 1 0 3512 0 1 2770
box -8 -3 16 105
use FILL  FILL_4710
timestamp 1677677812
transform 1 0 3520 0 1 2770
box -8 -3 16 105
use FILL  FILL_4711
timestamp 1677677812
transform 1 0 3528 0 1 2770
box -8 -3 16 105
use FILL  FILL_4712
timestamp 1677677812
transform 1 0 3536 0 1 2770
box -8 -3 16 105
use FILL  FILL_4713
timestamp 1677677812
transform 1 0 3544 0 1 2770
box -8 -3 16 105
use FILL  FILL_4714
timestamp 1677677812
transform 1 0 3552 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_197
timestamp 1677677812
transform -1 0 3600 0 1 2770
box -8 -3 46 105
use FILL  FILL_4715
timestamp 1677677812
transform 1 0 3600 0 1 2770
box -8 -3 16 105
use FILL  FILL_4716
timestamp 1677677812
transform 1 0 3608 0 1 2770
box -8 -3 16 105
use FILL  FILL_4717
timestamp 1677677812
transform 1 0 3616 0 1 2770
box -8 -3 16 105
use FILL  FILL_4718
timestamp 1677677812
transform 1 0 3624 0 1 2770
box -8 -3 16 105
use FILL  FILL_4719
timestamp 1677677812
transform 1 0 3632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4720
timestamp 1677677812
transform 1 0 3640 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_320
timestamp 1677677812
transform -1 0 3664 0 1 2770
box -9 -3 26 105
use FILL  FILL_4721
timestamp 1677677812
transform 1 0 3664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4731
timestamp 1677677812
transform 1 0 3672 0 1 2770
box -8 -3 16 105
use FILL  FILL_4733
timestamp 1677677812
transform 1 0 3680 0 1 2770
box -8 -3 16 105
use FILL  FILL_4735
timestamp 1677677812
transform 1 0 3688 0 1 2770
box -8 -3 16 105
use FILL  FILL_4737
timestamp 1677677812
transform 1 0 3696 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_24
timestamp 1677677812
transform -1 0 3736 0 1 2770
box -8 -3 40 105
use FILL  FILL_4738
timestamp 1677677812
transform 1 0 3736 0 1 2770
box -8 -3 16 105
use FILL  FILL_4739
timestamp 1677677812
transform 1 0 3744 0 1 2770
box -8 -3 16 105
use FILL  FILL_4740
timestamp 1677677812
transform 1 0 3752 0 1 2770
box -8 -3 16 105
use FILL  FILL_4741
timestamp 1677677812
transform 1 0 3760 0 1 2770
box -8 -3 16 105
use FILL  FILL_4742
timestamp 1677677812
transform 1 0 3768 0 1 2770
box -8 -3 16 105
use FILL  FILL_4743
timestamp 1677677812
transform 1 0 3776 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_25
timestamp 1677677812
transform -1 0 3816 0 1 2770
box -8 -3 40 105
use FILL  FILL_4744
timestamp 1677677812
transform 1 0 3816 0 1 2770
box -8 -3 16 105
use FILL  FILL_4749
timestamp 1677677812
transform 1 0 3824 0 1 2770
box -8 -3 16 105
use FILL  FILL_4750
timestamp 1677677812
transform 1 0 3832 0 1 2770
box -8 -3 16 105
use FILL  FILL_4751
timestamp 1677677812
transform 1 0 3840 0 1 2770
box -8 -3 16 105
use FILL  FILL_4753
timestamp 1677677812
transform 1 0 3848 0 1 2770
box -8 -3 16 105
use FILL  FILL_4755
timestamp 1677677812
transform 1 0 3856 0 1 2770
box -8 -3 16 105
use FILL  FILL_4757
timestamp 1677677812
transform 1 0 3864 0 1 2770
box -8 -3 16 105
use FILL  FILL_4759
timestamp 1677677812
transform 1 0 3872 0 1 2770
box -8 -3 16 105
use FILL  FILL_4761
timestamp 1677677812
transform 1 0 3880 0 1 2770
box -8 -3 16 105
use FILL  FILL_4762
timestamp 1677677812
transform 1 0 3888 0 1 2770
box -8 -3 16 105
use FILL  FILL_4763
timestamp 1677677812
transform 1 0 3896 0 1 2770
box -8 -3 16 105
use FILL  FILL_4764
timestamp 1677677812
transform 1 0 3904 0 1 2770
box -8 -3 16 105
use FILL  FILL_4765
timestamp 1677677812
transform 1 0 3912 0 1 2770
box -8 -3 16 105
use FILL  FILL_4766
timestamp 1677677812
transform 1 0 3920 0 1 2770
box -8 -3 16 105
use FILL  FILL_4768
timestamp 1677677812
transform 1 0 3928 0 1 2770
box -8 -3 16 105
use FILL  FILL_4770
timestamp 1677677812
transform 1 0 3936 0 1 2770
box -8 -3 16 105
use FILL  FILL_4772
timestamp 1677677812
transform 1 0 3944 0 1 2770
box -8 -3 16 105
use FILL  FILL_4773
timestamp 1677677812
transform 1 0 3952 0 1 2770
box -8 -3 16 105
use FILL  FILL_4774
timestamp 1677677812
transform 1 0 3960 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3649
timestamp 1677677812
transform 1 0 4052 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_286
timestamp 1677677812
transform 1 0 3968 0 1 2770
box -8 -3 104 105
use FILL  FILL_4775
timestamp 1677677812
transform 1 0 4064 0 1 2770
box -8 -3 16 105
use FILL  FILL_4776
timestamp 1677677812
transform 1 0 4072 0 1 2770
box -8 -3 16 105
use FILL  FILL_4777
timestamp 1677677812
transform 1 0 4080 0 1 2770
box -8 -3 16 105
use INVX2  INVX2_322
timestamp 1677677812
transform 1 0 4088 0 1 2770
box -9 -3 26 105
use FILL  FILL_4778
timestamp 1677677812
transform 1 0 4104 0 1 2770
box -8 -3 16 105
use FILL  FILL_4788
timestamp 1677677812
transform 1 0 4112 0 1 2770
box -8 -3 16 105
use FILL  FILL_4790
timestamp 1677677812
transform 1 0 4120 0 1 2770
box -8 -3 16 105
use FILL  FILL_4791
timestamp 1677677812
transform 1 0 4128 0 1 2770
box -8 -3 16 105
use FILL  FILL_4792
timestamp 1677677812
transform 1 0 4136 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_287
timestamp 1677677812
transform 1 0 4144 0 1 2770
box -8 -3 104 105
use FILL  FILL_4793
timestamp 1677677812
transform 1 0 4240 0 1 2770
box -8 -3 16 105
use FILL  FILL_4794
timestamp 1677677812
transform 1 0 4248 0 1 2770
box -8 -3 16 105
use FILL  FILL_4798
timestamp 1677677812
transform 1 0 4256 0 1 2770
box -8 -3 16 105
use FILL  FILL_4800
timestamp 1677677812
transform 1 0 4264 0 1 2770
box -8 -3 16 105
use FILL  FILL_4801
timestamp 1677677812
transform 1 0 4272 0 1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_26
timestamp 1677677812
transform 1 0 4280 0 1 2770
box -8 -3 40 105
use FILL  FILL_4802
timestamp 1677677812
transform 1 0 4312 0 1 2770
box -8 -3 16 105
use FILL  FILL_4803
timestamp 1677677812
transform 1 0 4320 0 1 2770
box -8 -3 16 105
use FILL  FILL_4804
timestamp 1677677812
transform 1 0 4328 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3650
timestamp 1677677812
transform 1 0 4348 0 1 2775
box -3 -3 3 3
use M3_M2  M3_M2_3651
timestamp 1677677812
transform 1 0 4436 0 1 2775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_289
timestamp 1677677812
transform 1 0 4336 0 1 2770
box -8 -3 104 105
use FILL  FILL_4807
timestamp 1677677812
transform 1 0 4432 0 1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_192
timestamp 1677677812
transform 1 0 4440 0 1 2770
box -8 -3 46 105
use FILL  FILL_4808
timestamp 1677677812
transform 1 0 4480 0 1 2770
box -8 -3 16 105
use FILL  FILL_4809
timestamp 1677677812
transform 1 0 4488 0 1 2770
box -8 -3 16 105
use FILL  FILL_4810
timestamp 1677677812
transform 1 0 4496 0 1 2770
box -8 -3 16 105
use FILL  FILL_4811
timestamp 1677677812
transform 1 0 4504 0 1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_198
timestamp 1677677812
transform 1 0 4512 0 1 2770
box -8 -3 46 105
use AOI22X1  AOI22X1_199
timestamp 1677677812
transform 1 0 4552 0 1 2770
box -8 -3 46 105
use FILL  FILL_4820
timestamp 1677677812
transform 1 0 4592 0 1 2770
box -8 -3 16 105
use FILL  FILL_4822
timestamp 1677677812
transform 1 0 4600 0 1 2770
box -8 -3 16 105
use FILL  FILL_4824
timestamp 1677677812
transform 1 0 4608 0 1 2770
box -8 -3 16 105
use FILL  FILL_4825
timestamp 1677677812
transform 1 0 4616 0 1 2770
box -8 -3 16 105
use FILL  FILL_4826
timestamp 1677677812
transform 1 0 4624 0 1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3652
timestamp 1677677812
transform 1 0 4644 0 1 2775
box -3 -3 3 3
use FILL  FILL_4827
timestamp 1677677812
transform 1 0 4632 0 1 2770
box -8 -3 16 105
use FILL  FILL_4830
timestamp 1677677812
transform 1 0 4640 0 1 2770
box -8 -3 16 105
use FILL  FILL_4831
timestamp 1677677812
transform 1 0 4648 0 1 2770
box -8 -3 16 105
use FILL  FILL_4832
timestamp 1677677812
transform 1 0 4656 0 1 2770
box -8 -3 16 105
use FILL  FILL_4833
timestamp 1677677812
transform 1 0 4664 0 1 2770
box -8 -3 16 105
use FILL  FILL_4834
timestamp 1677677812
transform 1 0 4672 0 1 2770
box -8 -3 16 105
use FILL  FILL_4835
timestamp 1677677812
transform 1 0 4680 0 1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_291
timestamp 1677677812
transform 1 0 4688 0 1 2770
box -8 -3 104 105
use FILL  FILL_4836
timestamp 1677677812
transform 1 0 4784 0 1 2770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_39
timestamp 1677677812
transform 1 0 4819 0 1 2770
box -10 -3 10 3
use M2_M1  M2_M1_4122
timestamp 1677677812
transform 1 0 92 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3782
timestamp 1677677812
transform 1 0 92 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4213
timestamp 1677677812
transform 1 0 108 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3690
timestamp 1677677812
transform 1 0 132 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4123
timestamp 1677677812
transform 1 0 132 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4124
timestamp 1677677812
transform 1 0 148 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4214
timestamp 1677677812
transform 1 0 124 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4215
timestamp 1677677812
transform 1 0 140 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3750
timestamp 1677677812
transform 1 0 148 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3691
timestamp 1677677812
transform 1 0 164 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4216
timestamp 1677677812
transform 1 0 156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3783
timestamp 1677677812
transform 1 0 140 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3812
timestamp 1677677812
transform 1 0 124 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3733
timestamp 1677677812
transform 1 0 180 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4125
timestamp 1677677812
transform 1 0 188 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4217
timestamp 1677677812
transform 1 0 180 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3784
timestamp 1677677812
transform 1 0 188 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4218
timestamp 1677677812
transform 1 0 204 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3734
timestamp 1677677812
transform 1 0 220 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4219
timestamp 1677677812
transform 1 0 220 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3845
timestamp 1677677812
transform 1 0 220 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3670
timestamp 1677677812
transform 1 0 236 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4126
timestamp 1677677812
transform 1 0 236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4127
timestamp 1677677812
transform 1 0 260 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4220
timestamp 1677677812
transform 1 0 244 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3785
timestamp 1677677812
transform 1 0 244 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3671
timestamp 1677677812
transform 1 0 324 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3692
timestamp 1677677812
transform 1 0 316 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4128
timestamp 1677677812
transform 1 0 300 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4129
timestamp 1677677812
transform 1 0 316 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4130
timestamp 1677677812
transform 1 0 324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4221
timestamp 1677677812
transform 1 0 284 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4222
timestamp 1677677812
transform 1 0 292 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4223
timestamp 1677677812
transform 1 0 308 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3786
timestamp 1677677812
transform 1 0 284 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3838
timestamp 1677677812
transform 1 0 292 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4224
timestamp 1677677812
transform 1 0 324 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3787
timestamp 1677677812
transform 1 0 324 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3839
timestamp 1677677812
transform 1 0 324 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4131
timestamp 1677677812
transform 1 0 348 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3751
timestamp 1677677812
transform 1 0 348 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3788
timestamp 1677677812
transform 1 0 348 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3672
timestamp 1677677812
transform 1 0 364 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3673
timestamp 1677677812
transform 1 0 404 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4132
timestamp 1677677812
transform 1 0 404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4225
timestamp 1677677812
transform 1 0 372 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4226
timestamp 1677677812
transform 1 0 388 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4227
timestamp 1677677812
transform 1 0 404 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3789
timestamp 1677677812
transform 1 0 372 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3813
timestamp 1677677812
transform 1 0 404 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3790
timestamp 1677677812
transform 1 0 420 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4133
timestamp 1677677812
transform 1 0 444 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4228
timestamp 1677677812
transform 1 0 468 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3791
timestamp 1677677812
transform 1 0 476 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3840
timestamp 1677677812
transform 1 0 476 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4229
timestamp 1677677812
transform 1 0 540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4230
timestamp 1677677812
transform 1 0 620 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3653
timestamp 1677677812
transform 1 0 652 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3674
timestamp 1677677812
transform 1 0 668 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3693
timestamp 1677677812
transform 1 0 644 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3694
timestamp 1677677812
transform 1 0 676 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4134
timestamp 1677677812
transform 1 0 652 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4135
timestamp 1677677812
transform 1 0 668 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4231
timestamp 1677677812
transform 1 0 660 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4232
timestamp 1677677812
transform 1 0 676 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3752
timestamp 1677677812
transform 1 0 692 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3792
timestamp 1677677812
transform 1 0 716 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3675
timestamp 1677677812
transform 1 0 796 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4136
timestamp 1677677812
transform 1 0 764 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4137
timestamp 1677677812
transform 1 0 772 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4233
timestamp 1677677812
transform 1 0 756 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3753
timestamp 1677677812
transform 1 0 772 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4138
timestamp 1677677812
transform 1 0 804 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4234
timestamp 1677677812
transform 1 0 780 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4235
timestamp 1677677812
transform 1 0 796 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3793
timestamp 1677677812
transform 1 0 772 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3846
timestamp 1677677812
transform 1 0 796 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4139
timestamp 1677677812
transform 1 0 852 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4140
timestamp 1677677812
transform 1 0 876 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3754
timestamp 1677677812
transform 1 0 876 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4236
timestamp 1677677812
transform 1 0 908 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3755
timestamp 1677677812
transform 1 0 924 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3847
timestamp 1677677812
transform 1 0 884 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3848
timestamp 1677677812
transform 1 0 940 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3654
timestamp 1677677812
transform 1 0 972 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4120
timestamp 1677677812
transform 1 0 972 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3756
timestamp 1677677812
transform 1 0 964 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3794
timestamp 1677677812
transform 1 0 972 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3841
timestamp 1677677812
transform 1 0 964 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4141
timestamp 1677677812
transform 1 0 988 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4237
timestamp 1677677812
transform 1 0 996 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3814
timestamp 1677677812
transform 1 0 996 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3655
timestamp 1677677812
transform 1 0 1044 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4142
timestamp 1677677812
transform 1 0 1036 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3849
timestamp 1677677812
transform 1 0 1036 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3695
timestamp 1677677812
transform 1 0 1052 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3656
timestamp 1677677812
transform 1 0 1076 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4143
timestamp 1677677812
transform 1 0 1060 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4144
timestamp 1677677812
transform 1 0 1068 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4145
timestamp 1677677812
transform 1 0 1084 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4238
timestamp 1677677812
transform 1 0 1052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4239
timestamp 1677677812
transform 1 0 1060 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3757
timestamp 1677677812
transform 1 0 1068 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4240
timestamp 1677677812
transform 1 0 1076 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4241
timestamp 1677677812
transform 1 0 1092 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3795
timestamp 1677677812
transform 1 0 1060 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3815
timestamp 1677677812
transform 1 0 1084 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3850
timestamp 1677677812
transform 1 0 1060 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4242
timestamp 1677677812
transform 1 0 1140 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3696
timestamp 1677677812
transform 1 0 1172 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4146
timestamp 1677677812
transform 1 0 1172 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3758
timestamp 1677677812
transform 1 0 1196 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4316
timestamp 1677677812
transform 1 0 1196 0 1 2715
box -2 -2 2 2
use M3_M2  M3_M2_3816
timestamp 1677677812
transform 1 0 1188 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3657
timestamp 1677677812
transform 1 0 1276 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3658
timestamp 1677677812
transform 1 0 1300 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4147
timestamp 1677677812
transform 1 0 1220 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3735
timestamp 1677677812
transform 1 0 1268 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4243
timestamp 1677677812
transform 1 0 1268 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3817
timestamp 1677677812
transform 1 0 1212 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4148
timestamp 1677677812
transform 1 0 1340 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3759
timestamp 1677677812
transform 1 0 1340 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4244
timestamp 1677677812
transform 1 0 1348 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4317
timestamp 1677677812
transform 1 0 1380 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4245
timestamp 1677677812
transform 1 0 1404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4149
timestamp 1677677812
transform 1 0 1420 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3818
timestamp 1677677812
transform 1 0 1420 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4150
timestamp 1677677812
transform 1 0 1452 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3736
timestamp 1677677812
transform 1 0 1460 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4246
timestamp 1677677812
transform 1 0 1444 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3760
timestamp 1677677812
transform 1 0 1452 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4151
timestamp 1677677812
transform 1 0 1492 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4247
timestamp 1677677812
transform 1 0 1484 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4248
timestamp 1677677812
transform 1 0 1500 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3819
timestamp 1677677812
transform 1 0 1484 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3697
timestamp 1677677812
transform 1 0 1572 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3761
timestamp 1677677812
transform 1 0 1580 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3698
timestamp 1677677812
transform 1 0 1612 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3762
timestamp 1677677812
transform 1 0 1604 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4152
timestamp 1677677812
transform 1 0 1628 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4249
timestamp 1677677812
transform 1 0 1628 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3820
timestamp 1677677812
transform 1 0 1628 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3699
timestamp 1677677812
transform 1 0 1660 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4153
timestamp 1677677812
transform 1 0 1660 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3763
timestamp 1677677812
transform 1 0 1684 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4250
timestamp 1677677812
transform 1 0 1708 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3821
timestamp 1677677812
transform 1 0 1724 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3851
timestamp 1677677812
transform 1 0 1724 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3852
timestamp 1677677812
transform 1 0 1804 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4251
timestamp 1677677812
transform 1 0 1820 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3700
timestamp 1677677812
transform 1 0 1852 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3701
timestamp 1677677812
transform 1 0 1876 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3702
timestamp 1677677812
transform 1 0 1932 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4154
timestamp 1677677812
transform 1 0 1852 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3737
timestamp 1677677812
transform 1 0 1900 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3738
timestamp 1677677812
transform 1 0 1940 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4252
timestamp 1677677812
transform 1 0 1900 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4253
timestamp 1677677812
transform 1 0 1932 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4254
timestamp 1677677812
transform 1 0 1940 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3822
timestamp 1677677812
transform 1 0 1852 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3823
timestamp 1677677812
transform 1 0 1892 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3764
timestamp 1677677812
transform 1 0 1980 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3676
timestamp 1677677812
transform 1 0 2004 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3703
timestamp 1677677812
transform 1 0 2036 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4155
timestamp 1677677812
transform 1 0 2012 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4156
timestamp 1677677812
transform 1 0 2020 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4157
timestamp 1677677812
transform 1 0 2036 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4255
timestamp 1677677812
transform 1 0 2004 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4256
timestamp 1677677812
transform 1 0 2028 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4257
timestamp 1677677812
transform 1 0 2052 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4258
timestamp 1677677812
transform 1 0 2068 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3853
timestamp 1677677812
transform 1 0 2068 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4158
timestamp 1677677812
transform 1 0 2108 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4159
timestamp 1677677812
transform 1 0 2124 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4259
timestamp 1677677812
transform 1 0 2100 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4260
timestamp 1677677812
transform 1 0 2116 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3739
timestamp 1677677812
transform 1 0 2132 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4160
timestamp 1677677812
transform 1 0 2172 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3677
timestamp 1677677812
transform 1 0 2188 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4261
timestamp 1677677812
transform 1 0 2180 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3659
timestamp 1677677812
transform 1 0 2212 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3678
timestamp 1677677812
transform 1 0 2236 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4161
timestamp 1677677812
transform 1 0 2236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4162
timestamp 1677677812
transform 1 0 2268 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4262
timestamp 1677677812
transform 1 0 2260 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4263
timestamp 1677677812
transform 1 0 2284 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3796
timestamp 1677677812
transform 1 0 2284 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3679
timestamp 1677677812
transform 1 0 2308 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4163
timestamp 1677677812
transform 1 0 2316 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4164
timestamp 1677677812
transform 1 0 2324 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4264
timestamp 1677677812
transform 1 0 2308 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4265
timestamp 1677677812
transform 1 0 2324 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3797
timestamp 1677677812
transform 1 0 2316 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3854
timestamp 1677677812
transform 1 0 2324 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3660
timestamp 1677677812
transform 1 0 2380 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3680
timestamp 1677677812
transform 1 0 2372 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4165
timestamp 1677677812
transform 1 0 2372 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4266
timestamp 1677677812
transform 1 0 2364 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3855
timestamp 1677677812
transform 1 0 2356 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3661
timestamp 1677677812
transform 1 0 2428 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3681
timestamp 1677677812
transform 1 0 2420 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3704
timestamp 1677677812
transform 1 0 2404 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4166
timestamp 1677677812
transform 1 0 2388 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4167
timestamp 1677677812
transform 1 0 2396 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4168
timestamp 1677677812
transform 1 0 2420 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3765
timestamp 1677677812
transform 1 0 2396 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4267
timestamp 1677677812
transform 1 0 2404 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4268
timestamp 1677677812
transform 1 0 2420 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3798
timestamp 1677677812
transform 1 0 2420 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3705
timestamp 1677677812
transform 1 0 2444 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4169
timestamp 1677677812
transform 1 0 2444 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3766
timestamp 1677677812
transform 1 0 2444 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3662
timestamp 1677677812
transform 1 0 2468 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4170
timestamp 1677677812
transform 1 0 2484 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4269
timestamp 1677677812
transform 1 0 2524 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4171
timestamp 1677677812
transform 1 0 2540 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4172
timestamp 1677677812
transform 1 0 2556 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4173
timestamp 1677677812
transform 1 0 2564 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4270
timestamp 1677677812
transform 1 0 2548 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3824
timestamp 1677677812
transform 1 0 2556 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4271
timestamp 1677677812
transform 1 0 2596 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3799
timestamp 1677677812
transform 1 0 2588 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3767
timestamp 1677677812
transform 1 0 2628 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3800
timestamp 1677677812
transform 1 0 2628 0 1 2715
box -3 -3 3 3
use M2_M1  M2_M1_4272
timestamp 1677677812
transform 1 0 2644 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3801
timestamp 1677677812
transform 1 0 2644 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3706
timestamp 1677677812
transform 1 0 2660 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4174
timestamp 1677677812
transform 1 0 2660 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3768
timestamp 1677677812
transform 1 0 2660 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3663
timestamp 1677677812
transform 1 0 2804 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3707
timestamp 1677677812
transform 1 0 2756 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3708
timestamp 1677677812
transform 1 0 2804 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4175
timestamp 1677677812
transform 1 0 2756 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4273
timestamp 1677677812
transform 1 0 2684 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4274
timestamp 1677677812
transform 1 0 2740 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4275
timestamp 1677677812
transform 1 0 2788 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3802
timestamp 1677677812
transform 1 0 2684 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3825
timestamp 1677677812
transform 1 0 2740 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3856
timestamp 1677677812
transform 1 0 2780 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3664
timestamp 1677677812
transform 1 0 2852 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4276
timestamp 1677677812
transform 1 0 2844 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4277
timestamp 1677677812
transform 1 0 2852 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4176
timestamp 1677677812
transform 1 0 2884 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3826
timestamp 1677677812
transform 1 0 2884 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3682
timestamp 1677677812
transform 1 0 2908 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4177
timestamp 1677677812
transform 1 0 2916 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4318
timestamp 1677677812
transform 1 0 2932 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4278
timestamp 1677677812
transform 1 0 2996 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4279
timestamp 1677677812
transform 1 0 3012 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3665
timestamp 1677677812
transform 1 0 3036 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4178
timestamp 1677677812
transform 1 0 3036 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3827
timestamp 1677677812
transform 1 0 3028 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3709
timestamp 1677677812
transform 1 0 3052 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3710
timestamp 1677677812
transform 1 0 3076 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4179
timestamp 1677677812
transform 1 0 3124 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4280
timestamp 1677677812
transform 1 0 3076 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3711
timestamp 1677677812
transform 1 0 3172 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4180
timestamp 1677677812
transform 1 0 3172 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3712
timestamp 1677677812
transform 1 0 3196 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4181
timestamp 1677677812
transform 1 0 3196 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4281
timestamp 1677677812
transform 1 0 3196 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3828
timestamp 1677677812
transform 1 0 3196 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3666
timestamp 1677677812
transform 1 0 3212 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3713
timestamp 1677677812
transform 1 0 3212 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3714
timestamp 1677677812
transform 1 0 3228 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4182
timestamp 1677677812
transform 1 0 3220 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4183
timestamp 1677677812
transform 1 0 3236 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4184
timestamp 1677677812
transform 1 0 3252 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4282
timestamp 1677677812
transform 1 0 3228 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4283
timestamp 1677677812
transform 1 0 3244 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3803
timestamp 1677677812
transform 1 0 3236 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3829
timestamp 1677677812
transform 1 0 3244 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4185
timestamp 1677677812
transform 1 0 3268 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3769
timestamp 1677677812
transform 1 0 3268 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4284
timestamp 1677677812
transform 1 0 3276 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4121
timestamp 1677677812
transform 1 0 3300 0 1 2745
box -2 -2 2 2
use M3_M2  M3_M2_3740
timestamp 1677677812
transform 1 0 3300 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3770
timestamp 1677677812
transform 1 0 3364 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4285
timestamp 1677677812
transform 1 0 3380 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3771
timestamp 1677677812
transform 1 0 3404 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3857
timestamp 1677677812
transform 1 0 3412 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3715
timestamp 1677677812
transform 1 0 3452 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3683
timestamp 1677677812
transform 1 0 3500 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4186
timestamp 1677677812
transform 1 0 3476 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4286
timestamp 1677677812
transform 1 0 3516 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3804
timestamp 1677677812
transform 1 0 3516 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3805
timestamp 1677677812
transform 1 0 3548 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3830
timestamp 1677677812
transform 1 0 3468 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3831
timestamp 1677677812
transform 1 0 3524 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3858
timestamp 1677677812
transform 1 0 3492 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3741
timestamp 1677677812
transform 1 0 3564 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4287
timestamp 1677677812
transform 1 0 3580 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3859
timestamp 1677677812
transform 1 0 3572 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3716
timestamp 1677677812
transform 1 0 3596 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3684
timestamp 1677677812
transform 1 0 3644 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3717
timestamp 1677677812
transform 1 0 3612 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3718
timestamp 1677677812
transform 1 0 3636 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4187
timestamp 1677677812
transform 1 0 3612 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4188
timestamp 1677677812
transform 1 0 3628 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3742
timestamp 1677677812
transform 1 0 3636 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4189
timestamp 1677677812
transform 1 0 3644 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3772
timestamp 1677677812
transform 1 0 3612 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4288
timestamp 1677677812
transform 1 0 3620 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4289
timestamp 1677677812
transform 1 0 3636 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3719
timestamp 1677677812
transform 1 0 3660 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4290
timestamp 1677677812
transform 1 0 3652 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3720
timestamp 1677677812
transform 1 0 3724 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4190
timestamp 1677677812
transform 1 0 3724 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3743
timestamp 1677677812
transform 1 0 3772 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3773
timestamp 1677677812
transform 1 0 3748 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4291
timestamp 1677677812
transform 1 0 3772 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3721
timestamp 1677677812
transform 1 0 3836 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4191
timestamp 1677677812
transform 1 0 3844 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3722
timestamp 1677677812
transform 1 0 3876 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3744
timestamp 1677677812
transform 1 0 3892 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4192
timestamp 1677677812
transform 1 0 3900 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4292
timestamp 1677677812
transform 1 0 3884 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4293
timestamp 1677677812
transform 1 0 3892 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4294
timestamp 1677677812
transform 1 0 3908 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3806
timestamp 1677677812
transform 1 0 3884 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3807
timestamp 1677677812
transform 1 0 3908 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3832
timestamp 1677677812
transform 1 0 3892 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4322
timestamp 1677677812
transform 1 0 3932 0 1 2685
box -2 -2 2 2
use M3_M2  M3_M2_3667
timestamp 1677677812
transform 1 0 3948 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3685
timestamp 1677677812
transform 1 0 3956 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3723
timestamp 1677677812
transform 1 0 3980 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4193
timestamp 1677677812
transform 1 0 3948 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4194
timestamp 1677677812
transform 1 0 3964 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3745
timestamp 1677677812
transform 1 0 3972 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4195
timestamp 1677677812
transform 1 0 3980 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4295
timestamp 1677677812
transform 1 0 3956 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4296
timestamp 1677677812
transform 1 0 3972 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3808
timestamp 1677677812
transform 1 0 3956 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3860
timestamp 1677677812
transform 1 0 3948 0 1 2685
box -3 -3 3 3
use M2_M1  M2_M1_4297
timestamp 1677677812
transform 1 0 3988 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3833
timestamp 1677677812
transform 1 0 4012 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3861
timestamp 1677677812
transform 1 0 4028 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3724
timestamp 1677677812
transform 1 0 4044 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3746
timestamp 1677677812
transform 1 0 4044 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3686
timestamp 1677677812
transform 1 0 4084 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3725
timestamp 1677677812
transform 1 0 4060 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3726
timestamp 1677677812
transform 1 0 4076 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4196
timestamp 1677677812
transform 1 0 4052 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4197
timestamp 1677677812
transform 1 0 4060 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4198
timestamp 1677677812
transform 1 0 4076 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4199
timestamp 1677677812
transform 1 0 4092 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3774
timestamp 1677677812
transform 1 0 4036 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4298
timestamp 1677677812
transform 1 0 4044 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3809
timestamp 1677677812
transform 1 0 4044 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3747
timestamp 1677677812
transform 1 0 4100 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3775
timestamp 1677677812
transform 1 0 4068 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4299
timestamp 1677677812
transform 1 0 4084 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3776
timestamp 1677677812
transform 1 0 4092 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3834
timestamp 1677677812
transform 1 0 4092 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3727
timestamp 1677677812
transform 1 0 4156 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4200
timestamp 1677677812
transform 1 0 4132 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4300
timestamp 1677677812
transform 1 0 4156 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3862
timestamp 1677677812
transform 1 0 4148 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3863
timestamp 1677677812
transform 1 0 4196 0 1 2685
box -3 -3 3 3
use M3_M2  M3_M2_3687
timestamp 1677677812
transform 1 0 4236 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4301
timestamp 1677677812
transform 1 0 4244 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4302
timestamp 1677677812
transform 1 0 4252 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4201
timestamp 1677677812
transform 1 0 4292 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3777
timestamp 1677677812
transform 1 0 4292 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4303
timestamp 1677677812
transform 1 0 4316 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4319
timestamp 1677677812
transform 1 0 4300 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4321
timestamp 1677677812
transform 1 0 4308 0 1 2705
box -2 -2 2 2
use M3_M2  M3_M2_3842
timestamp 1677677812
transform 1 0 4308 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4320
timestamp 1677677812
transform 1 0 4332 0 1 2715
box -2 -2 2 2
use M2_M1  M2_M1_4304
timestamp 1677677812
transform 1 0 4348 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4305
timestamp 1677677812
transform 1 0 4364 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3843
timestamp 1677677812
transform 1 0 4364 0 1 2695
box -3 -3 3 3
use M2_M1  M2_M1_4202
timestamp 1677677812
transform 1 0 4388 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3778
timestamp 1677677812
transform 1 0 4380 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3668
timestamp 1677677812
transform 1 0 4404 0 1 2765
box -3 -3 3 3
use M3_M2  M3_M2_3728
timestamp 1677677812
transform 1 0 4412 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4203
timestamp 1677677812
transform 1 0 4404 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4306
timestamp 1677677812
transform 1 0 4412 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3835
timestamp 1677677812
transform 1 0 4404 0 1 2705
box -3 -3 3 3
use M3_M2  M3_M2_3779
timestamp 1677677812
transform 1 0 4420 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4204
timestamp 1677677812
transform 1 0 4444 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4307
timestamp 1677677812
transform 1 0 4468 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3844
timestamp 1677677812
transform 1 0 4468 0 1 2695
box -3 -3 3 3
use M3_M2  M3_M2_3688
timestamp 1677677812
transform 1 0 4564 0 1 2755
box -3 -3 3 3
use M3_M2  M3_M2_3729
timestamp 1677677812
transform 1 0 4556 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3689
timestamp 1677677812
transform 1 0 4596 0 1 2755
box -3 -3 3 3
use M2_M1  M2_M1_4205
timestamp 1677677812
transform 1 0 4556 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4206
timestamp 1677677812
transform 1 0 4572 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4207
timestamp 1677677812
transform 1 0 4588 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4308
timestamp 1677677812
transform 1 0 4540 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4309
timestamp 1677677812
transform 1 0 4548 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3780
timestamp 1677677812
transform 1 0 4556 0 1 2725
box -3 -3 3 3
use M2_M1  M2_M1_4310
timestamp 1677677812
transform 1 0 4580 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3836
timestamp 1677677812
transform 1 0 4556 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4311
timestamp 1677677812
transform 1 0 4596 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3730
timestamp 1677677812
transform 1 0 4612 0 1 2745
box -3 -3 3 3
use M3_M2  M3_M2_3669
timestamp 1677677812
transform 1 0 4628 0 1 2765
box -3 -3 3 3
use M2_M1  M2_M1_4208
timestamp 1677677812
transform 1 0 4628 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3781
timestamp 1677677812
transform 1 0 4620 0 1 2725
box -3 -3 3 3
use M3_M2  M3_M2_3731
timestamp 1677677812
transform 1 0 4660 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4209
timestamp 1677677812
transform 1 0 4644 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4210
timestamp 1677677812
transform 1 0 4660 0 1 2735
box -2 -2 2 2
use M3_M2  M3_M2_3748
timestamp 1677677812
transform 1 0 4668 0 1 2735
box -3 -3 3 3
use M3_M2  M3_M2_3732
timestamp 1677677812
transform 1 0 4716 0 1 2745
box -3 -3 3 3
use M2_M1  M2_M1_4211
timestamp 1677677812
transform 1 0 4676 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4212
timestamp 1677677812
transform 1 0 4692 0 1 2735
box -2 -2 2 2
use M2_M1  M2_M1_4312
timestamp 1677677812
transform 1 0 4652 0 1 2725
box -2 -2 2 2
use M2_M1  M2_M1_4313
timestamp 1677677812
transform 1 0 4668 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3810
timestamp 1677677812
transform 1 0 4668 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3837
timestamp 1677677812
transform 1 0 4644 0 1 2705
box -3 -3 3 3
use M2_M1  M2_M1_4314
timestamp 1677677812
transform 1 0 4716 0 1 2725
box -2 -2 2 2
use M3_M2  M3_M2_3811
timestamp 1677677812
transform 1 0 4732 0 1 2715
box -3 -3 3 3
use M3_M2  M3_M2_3749
timestamp 1677677812
transform 1 0 4788 0 1 2735
box -3 -3 3 3
use M2_M1  M2_M1_4315
timestamp 1677677812
transform 1 0 4788 0 1 2725
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_40
timestamp 1677677812
transform 1 0 24 0 1 2670
box -10 -3 10 3
use FILL  FILL_4316
timestamp 1677677812
transform 1 0 72 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4317
timestamp 1677677812
transform 1 0 80 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_298
timestamp 1677677812
transform 1 0 88 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4318
timestamp 1677677812
transform 1 0 104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4319
timestamp 1677677812
transform 1 0 112 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_183
timestamp 1677677812
transform -1 0 160 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4320
timestamp 1677677812
transform 1 0 160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4321
timestamp 1677677812
transform 1 0 168 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4322
timestamp 1677677812
transform 1 0 176 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_299
timestamp 1677677812
transform 1 0 184 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4323
timestamp 1677677812
transform 1 0 200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4324
timestamp 1677677812
transform 1 0 208 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4325
timestamp 1677677812
transform 1 0 216 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_184
timestamp 1677677812
transform 1 0 224 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4326
timestamp 1677677812
transform 1 0 264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4327
timestamp 1677677812
transform 1 0 272 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_178
timestamp 1677677812
transform 1 0 280 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4328
timestamp 1677677812
transform 1 0 320 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_300
timestamp 1677677812
transform 1 0 328 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4329
timestamp 1677677812
transform 1 0 344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4330
timestamp 1677677812
transform 1 0 352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4331
timestamp 1677677812
transform 1 0 360 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_185
timestamp 1677677812
transform 1 0 368 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4332
timestamp 1677677812
transform 1 0 408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4333
timestamp 1677677812
transform 1 0 416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4335
timestamp 1677677812
transform 1 0 424 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_267
timestamp 1677677812
transform 1 0 432 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4337
timestamp 1677677812
transform 1 0 528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4340
timestamp 1677677812
transform 1 0 536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4341
timestamp 1677677812
transform 1 0 544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4342
timestamp 1677677812
transform 1 0 552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4343
timestamp 1677677812
transform 1 0 560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4345
timestamp 1677677812
transform 1 0 568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4348
timestamp 1677677812
transform 1 0 576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4349
timestamp 1677677812
transform 1 0 584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4350
timestamp 1677677812
transform 1 0 592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4351
timestamp 1677677812
transform 1 0 600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4352
timestamp 1677677812
transform 1 0 608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4353
timestamp 1677677812
transform 1 0 616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4354
timestamp 1677677812
transform 1 0 624 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3864
timestamp 1677677812
transform 1 0 660 0 1 2675
box -3 -3 3 3
use OAI22X1  OAI22X1_179
timestamp 1677677812
transform 1 0 632 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4355
timestamp 1677677812
transform 1 0 672 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3865
timestamp 1677677812
transform 1 0 692 0 1 2675
box -3 -3 3 3
use FILL  FILL_4356
timestamp 1677677812
transform 1 0 680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4361
timestamp 1677677812
transform 1 0 688 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_302
timestamp 1677677812
transform -1 0 712 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4362
timestamp 1677677812
transform 1 0 712 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4363
timestamp 1677677812
transform 1 0 720 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4364
timestamp 1677677812
transform 1 0 728 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3866
timestamp 1677677812
transform 1 0 748 0 1 2675
box -3 -3 3 3
use FILL  FILL_4365
timestamp 1677677812
transform 1 0 736 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4366
timestamp 1677677812
transform 1 0 744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4374
timestamp 1677677812
transform 1 0 752 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_186
timestamp 1677677812
transform -1 0 800 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4375
timestamp 1677677812
transform 1 0 800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4378
timestamp 1677677812
transform 1 0 808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4379
timestamp 1677677812
transform 1 0 816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4380
timestamp 1677677812
transform 1 0 824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4381
timestamp 1677677812
transform 1 0 832 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4382
timestamp 1677677812
transform 1 0 840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4383
timestamp 1677677812
transform 1 0 848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4384
timestamp 1677677812
transform 1 0 856 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_269
timestamp 1677677812
transform 1 0 864 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4396
timestamp 1677677812
transform 1 0 960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4398
timestamp 1677677812
transform 1 0 968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4400
timestamp 1677677812
transform 1 0 976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4402
timestamp 1677677812
transform 1 0 984 0 -1 2770
box -8 -3 16 105
use NOR2X1  NOR2X1_46
timestamp 1677677812
transform 1 0 992 0 -1 2770
box -8 -3 32 105
use FILL  FILL_4404
timestamp 1677677812
transform 1 0 1016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4405
timestamp 1677677812
transform 1 0 1024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4406
timestamp 1677677812
transform 1 0 1032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4408
timestamp 1677677812
transform 1 0 1040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4410
timestamp 1677677812
transform 1 0 1048 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_189
timestamp 1677677812
transform 1 0 1056 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4417
timestamp 1677677812
transform 1 0 1096 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3867
timestamp 1677677812
transform 1 0 1116 0 1 2675
box -3 -3 3 3
use FILL  FILL_4419
timestamp 1677677812
transform 1 0 1104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4421
timestamp 1677677812
transform 1 0 1112 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4423
timestamp 1677677812
transform 1 0 1120 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3868
timestamp 1677677812
transform 1 0 1140 0 1 2675
box -3 -3 3 3
use FILL  FILL_4433
timestamp 1677677812
transform 1 0 1128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4434
timestamp 1677677812
transform 1 0 1136 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_94
timestamp 1677677812
transform 1 0 1144 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4435
timestamp 1677677812
transform 1 0 1176 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4436
timestamp 1677677812
transform 1 0 1184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4437
timestamp 1677677812
transform 1 0 1192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4438
timestamp 1677677812
transform 1 0 1200 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3869
timestamp 1677677812
transform 1 0 1228 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_271
timestamp 1677677812
transform 1 0 1208 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4439
timestamp 1677677812
transform 1 0 1304 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4441
timestamp 1677677812
transform 1 0 1312 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_305
timestamp 1677677812
transform 1 0 1320 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4445
timestamp 1677677812
transform 1 0 1336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4447
timestamp 1677677812
transform 1 0 1344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4449
timestamp 1677677812
transform 1 0 1352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4451
timestamp 1677677812
transform 1 0 1360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4458
timestamp 1677677812
transform 1 0 1368 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_95
timestamp 1677677812
transform -1 0 1408 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4459
timestamp 1677677812
transform 1 0 1408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4461
timestamp 1677677812
transform 1 0 1416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4463
timestamp 1677677812
transform 1 0 1424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4465
timestamp 1677677812
transform 1 0 1432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4471
timestamp 1677677812
transform 1 0 1440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4472
timestamp 1677677812
transform 1 0 1448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4473
timestamp 1677677812
transform 1 0 1456 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4474
timestamp 1677677812
transform 1 0 1464 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_181
timestamp 1677677812
transform -1 0 1512 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4475
timestamp 1677677812
transform 1 0 1512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4477
timestamp 1677677812
transform 1 0 1520 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4479
timestamp 1677677812
transform 1 0 1528 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4481
timestamp 1677677812
transform 1 0 1536 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4483
timestamp 1677677812
transform 1 0 1544 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4485
timestamp 1677677812
transform 1 0 1552 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4501
timestamp 1677677812
transform 1 0 1560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4502
timestamp 1677677812
transform 1 0 1568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4503
timestamp 1677677812
transform 1 0 1576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4504
timestamp 1677677812
transform 1 0 1584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4505
timestamp 1677677812
transform 1 0 1592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4506
timestamp 1677677812
transform 1 0 1600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4507
timestamp 1677677812
transform 1 0 1608 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4508
timestamp 1677677812
transform 1 0 1616 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4509
timestamp 1677677812
transform 1 0 1624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4510
timestamp 1677677812
transform 1 0 1632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4511
timestamp 1677677812
transform 1 0 1640 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_276
timestamp 1677677812
transform 1 0 1648 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4512
timestamp 1677677812
transform 1 0 1744 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4513
timestamp 1677677812
transform 1 0 1752 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4514
timestamp 1677677812
transform 1 0 1760 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4515
timestamp 1677677812
transform 1 0 1768 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4516
timestamp 1677677812
transform 1 0 1776 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_308
timestamp 1677677812
transform 1 0 1784 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4517
timestamp 1677677812
transform 1 0 1800 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4518
timestamp 1677677812
transform 1 0 1808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4519
timestamp 1677677812
transform 1 0 1816 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4520
timestamp 1677677812
transform 1 0 1824 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4521
timestamp 1677677812
transform 1 0 1832 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_277
timestamp 1677677812
transform 1 0 1840 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4522
timestamp 1677677812
transform 1 0 1936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4523
timestamp 1677677812
transform 1 0 1944 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_309
timestamp 1677677812
transform -1 0 1968 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4524
timestamp 1677677812
transform 1 0 1968 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4525
timestamp 1677677812
transform 1 0 1976 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4526
timestamp 1677677812
transform 1 0 1984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4527
timestamp 1677677812
transform 1 0 1992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4528
timestamp 1677677812
transform 1 0 2000 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3870
timestamp 1677677812
transform 1 0 2020 0 1 2675
box -3 -3 3 3
use AOI22X1  AOI22X1_190
timestamp 1677677812
transform 1 0 2008 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4529
timestamp 1677677812
transform 1 0 2048 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4530
timestamp 1677677812
transform 1 0 2056 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3871
timestamp 1677677812
transform 1 0 2076 0 1 2675
box -3 -3 3 3
use FILL  FILL_4531
timestamp 1677677812
transform 1 0 2064 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4532
timestamp 1677677812
transform 1 0 2072 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4533
timestamp 1677677812
transform 1 0 2080 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_183
timestamp 1677677812
transform -1 0 2128 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4534
timestamp 1677677812
transform 1 0 2128 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4536
timestamp 1677677812
transform 1 0 2136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4539
timestamp 1677677812
transform 1 0 2144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4540
timestamp 1677677812
transform 1 0 2152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4541
timestamp 1677677812
transform 1 0 2160 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_310
timestamp 1677677812
transform 1 0 2168 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4542
timestamp 1677677812
transform 1 0 2184 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4543
timestamp 1677677812
transform 1 0 2192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4545
timestamp 1677677812
transform 1 0 2200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4547
timestamp 1677677812
transform 1 0 2208 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3872
timestamp 1677677812
transform 1 0 2228 0 1 2675
box -3 -3 3 3
use FILL  FILL_4549
timestamp 1677677812
transform 1 0 2216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4551
timestamp 1677677812
transform 1 0 2224 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_311
timestamp 1677677812
transform 1 0 2232 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4555
timestamp 1677677812
transform 1 0 2248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4557
timestamp 1677677812
transform 1 0 2256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4559
timestamp 1677677812
transform 1 0 2264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4561
timestamp 1677677812
transform 1 0 2272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4563
timestamp 1677677812
transform 1 0 2280 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_192
timestamp 1677677812
transform 1 0 2288 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4570
timestamp 1677677812
transform 1 0 2328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4572
timestamp 1677677812
transform 1 0 2336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4574
timestamp 1677677812
transform 1 0 2344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4576
timestamp 1677677812
transform 1 0 2352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4581
timestamp 1677677812
transform 1 0 2360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4582
timestamp 1677677812
transform 1 0 2368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4583
timestamp 1677677812
transform 1 0 2376 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_194
timestamp 1677677812
transform -1 0 2424 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4584
timestamp 1677677812
transform 1 0 2424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4586
timestamp 1677677812
transform 1 0 2432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4588
timestamp 1677677812
transform 1 0 2440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4591
timestamp 1677677812
transform 1 0 2448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4592
timestamp 1677677812
transform 1 0 2456 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_312
timestamp 1677677812
transform 1 0 2464 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4593
timestamp 1677677812
transform 1 0 2480 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4594
timestamp 1677677812
transform 1 0 2488 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4595
timestamp 1677677812
transform 1 0 2496 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4597
timestamp 1677677812
transform 1 0 2504 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4599
timestamp 1677677812
transform 1 0 2512 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4601
timestamp 1677677812
transform 1 0 2520 0 -1 2770
box -8 -3 16 105
use AOI22X1  AOI22X1_196
timestamp 1677677812
transform 1 0 2528 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4605
timestamp 1677677812
transform 1 0 2568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4606
timestamp 1677677812
transform 1 0 2576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4607
timestamp 1677677812
transform 1 0 2584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4609
timestamp 1677677812
transform 1 0 2592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4611
timestamp 1677677812
transform 1 0 2600 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_314
timestamp 1677677812
transform 1 0 2608 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4613
timestamp 1677677812
transform 1 0 2624 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4615
timestamp 1677677812
transform 1 0 2632 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4617
timestamp 1677677812
transform 1 0 2640 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_279
timestamp 1677677812
transform 1 0 2648 0 -1 2770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_280
timestamp 1677677812
transform 1 0 2744 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4625
timestamp 1677677812
transform 1 0 2840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4626
timestamp 1677677812
transform 1 0 2848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4628
timestamp 1677677812
transform 1 0 2856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4635
timestamp 1677677812
transform 1 0 2864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4636
timestamp 1677677812
transform 1 0 2872 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4637
timestamp 1677677812
transform 1 0 2880 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_98
timestamp 1677677812
transform 1 0 2888 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4638
timestamp 1677677812
transform 1 0 2920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4639
timestamp 1677677812
transform 1 0 2928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4640
timestamp 1677677812
transform 1 0 2936 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4641
timestamp 1677677812
transform 1 0 2944 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4642
timestamp 1677677812
transform 1 0 2952 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4643
timestamp 1677677812
transform 1 0 2960 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4648
timestamp 1677677812
transform 1 0 2968 0 -1 2770
box -8 -3 16 105
use OAI21X1  OAI21X1_99
timestamp 1677677812
transform -1 0 3008 0 -1 2770
box -8 -3 34 105
use FILL  FILL_4649
timestamp 1677677812
transform 1 0 3008 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4651
timestamp 1677677812
transform 1 0 3016 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4661
timestamp 1677677812
transform 1 0 3024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4662
timestamp 1677677812
transform 1 0 3032 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_283
timestamp 1677677812
transform -1 0 3136 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4663
timestamp 1677677812
transform 1 0 3136 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4664
timestamp 1677677812
transform 1 0 3144 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4665
timestamp 1677677812
transform 1 0 3152 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4666
timestamp 1677677812
transform 1 0 3160 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4667
timestamp 1677677812
transform 1 0 3168 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_317
timestamp 1677677812
transform 1 0 3176 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4668
timestamp 1677677812
transform 1 0 3192 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4669
timestamp 1677677812
transform 1 0 3200 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4670
timestamp 1677677812
transform 1 0 3208 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_187
timestamp 1677677812
transform -1 0 3256 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4671
timestamp 1677677812
transform 1 0 3256 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4672
timestamp 1677677812
transform 1 0 3264 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4673
timestamp 1677677812
transform 1 0 3272 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4674
timestamp 1677677812
transform 1 0 3280 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3873
timestamp 1677677812
transform 1 0 3300 0 1 2675
box -3 -3 3 3
use FILL  FILL_4675
timestamp 1677677812
transform 1 0 3288 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4676
timestamp 1677677812
transform 1 0 3296 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4677
timestamp 1677677812
transform 1 0 3304 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_318
timestamp 1677677812
transform 1 0 3312 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4678
timestamp 1677677812
transform 1 0 3328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4679
timestamp 1677677812
transform 1 0 3336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4680
timestamp 1677677812
transform 1 0 3344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4681
timestamp 1677677812
transform 1 0 3352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4682
timestamp 1677677812
transform 1 0 3360 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4683
timestamp 1677677812
transform 1 0 3368 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4684
timestamp 1677677812
transform 1 0 3376 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4686
timestamp 1677677812
transform 1 0 3384 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4687
timestamp 1677677812
transform 1 0 3392 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4688
timestamp 1677677812
transform 1 0 3400 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4690
timestamp 1677677812
transform 1 0 3408 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4692
timestamp 1677677812
transform 1 0 3416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4694
timestamp 1677677812
transform 1 0 3424 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4696
timestamp 1677677812
transform 1 0 3432 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4698
timestamp 1677677812
transform 1 0 3440 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4700
timestamp 1677677812
transform 1 0 3448 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4702
timestamp 1677677812
transform 1 0 3456 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3874
timestamp 1677677812
transform 1 0 3476 0 1 2675
box -3 -3 3 3
use M3_M2  M3_M2_3875
timestamp 1677677812
transform 1 0 3516 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_284
timestamp 1677677812
transform 1 0 3464 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4722
timestamp 1677677812
transform 1 0 3560 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4723
timestamp 1677677812
transform 1 0 3568 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4724
timestamp 1677677812
transform 1 0 3576 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4725
timestamp 1677677812
transform 1 0 3584 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4726
timestamp 1677677812
transform 1 0 3592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4727
timestamp 1677677812
transform 1 0 3600 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_188
timestamp 1677677812
transform -1 0 3648 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4728
timestamp 1677677812
transform 1 0 3648 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4729
timestamp 1677677812
transform 1 0 3656 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4730
timestamp 1677677812
transform 1 0 3664 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4732
timestamp 1677677812
transform 1 0 3672 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4734
timestamp 1677677812
transform 1 0 3680 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4736
timestamp 1677677812
transform 1 0 3688 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4745
timestamp 1677677812
transform 1 0 3696 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4746
timestamp 1677677812
transform 1 0 3704 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_285
timestamp 1677677812
transform 1 0 3712 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4747
timestamp 1677677812
transform 1 0 3808 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4748
timestamp 1677677812
transform 1 0 3816 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_321
timestamp 1677677812
transform 1 0 3824 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4752
timestamp 1677677812
transform 1 0 3840 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4754
timestamp 1677677812
transform 1 0 3848 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4756
timestamp 1677677812
transform 1 0 3856 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4758
timestamp 1677677812
transform 1 0 3864 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4760
timestamp 1677677812
transform 1 0 3872 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_189
timestamp 1677677812
transform 1 0 3880 0 -1 2770
box -8 -3 46 105
use M3_M2  M3_M2_3876
timestamp 1677677812
transform 1 0 3932 0 1 2675
box -3 -3 3 3
use FILL  FILL_4767
timestamp 1677677812
transform 1 0 3920 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4769
timestamp 1677677812
transform 1 0 3928 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4771
timestamp 1677677812
transform 1 0 3936 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_190
timestamp 1677677812
transform 1 0 3944 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4779
timestamp 1677677812
transform 1 0 3984 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4780
timestamp 1677677812
transform 1 0 3992 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4781
timestamp 1677677812
transform 1 0 4000 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3877
timestamp 1677677812
transform 1 0 4020 0 1 2675
box -3 -3 3 3
use INVX2  INVX2_323
timestamp 1677677812
transform -1 0 4024 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4782
timestamp 1677677812
transform 1 0 4024 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4783
timestamp 1677677812
transform 1 0 4032 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4784
timestamp 1677677812
transform 1 0 4040 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4785
timestamp 1677677812
transform 1 0 4048 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3878
timestamp 1677677812
transform 1 0 4084 0 1 2675
box -3 -3 3 3
use OAI22X1  OAI22X1_191
timestamp 1677677812
transform 1 0 4056 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4786
timestamp 1677677812
transform 1 0 4096 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4787
timestamp 1677677812
transform 1 0 4104 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4789
timestamp 1677677812
transform 1 0 4112 0 -1 2770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_288
timestamp 1677677812
transform 1 0 4120 0 -1 2770
box -8 -3 104 105
use FILL  FILL_4795
timestamp 1677677812
transform 1 0 4216 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4796
timestamp 1677677812
transform 1 0 4224 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3879
timestamp 1677677812
transform 1 0 4252 0 1 2675
box -3 -3 3 3
use INVX2  INVX2_324
timestamp 1677677812
transform 1 0 4232 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4797
timestamp 1677677812
transform 1 0 4248 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4799
timestamp 1677677812
transform 1 0 4256 0 -1 2770
box -8 -3 16 105
use BUFX2  BUFX2_33
timestamp 1677677812
transform 1 0 4264 0 -1 2770
box -5 -3 28 105
use FILL  FILL_4805
timestamp 1677677812
transform 1 0 4288 0 -1 2770
box -8 -3 16 105
use NAND3X1  NAND3X1_27
timestamp 1677677812
transform -1 0 4328 0 -1 2770
box -8 -3 40 105
use FILL  FILL_4806
timestamp 1677677812
transform 1 0 4328 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4812
timestamp 1677677812
transform 1 0 4336 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4813
timestamp 1677677812
transform 1 0 4344 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4814
timestamp 1677677812
transform 1 0 4352 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4815
timestamp 1677677812
transform 1 0 4360 0 -1 2770
box -8 -3 16 105
use BUFX2  BUFX2_34
timestamp 1677677812
transform 1 0 4368 0 -1 2770
box -5 -3 28 105
use FILL  FILL_4816
timestamp 1677677812
transform 1 0 4392 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_325
timestamp 1677677812
transform 1 0 4400 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4817
timestamp 1677677812
transform 1 0 4416 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4818
timestamp 1677677812
transform 1 0 4424 0 -1 2770
box -8 -3 16 105
use M3_M2  M3_M2_3880
timestamp 1677677812
transform 1 0 4508 0 1 2675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_290
timestamp 1677677812
transform 1 0 4432 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_326
timestamp 1677677812
transform 1 0 4528 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4819
timestamp 1677677812
transform 1 0 4544 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_193
timestamp 1677677812
transform 1 0 4552 0 -1 2770
box -8 -3 46 105
use FILL  FILL_4821
timestamp 1677677812
transform 1 0 4592 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4823
timestamp 1677677812
transform 1 0 4600 0 -1 2770
box -8 -3 16 105
use FILL  FILL_4828
timestamp 1677677812
transform 1 0 4608 0 -1 2770
box -8 -3 16 105
use INVX2  INVX2_327
timestamp 1677677812
transform -1 0 4632 0 -1 2770
box -9 -3 26 105
use FILL  FILL_4829
timestamp 1677677812
transform 1 0 4632 0 -1 2770
box -8 -3 16 105
use OAI22X1  OAI22X1_194
timestamp 1677677812
transform 1 0 4640 0 -1 2770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_292
timestamp 1677677812
transform 1 0 4680 0 -1 2770
box -8 -3 104 105
use INVX2  INVX2_328
timestamp 1677677812
transform 1 0 4776 0 -1 2770
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_41
timestamp 1677677812
transform 1 0 4843 0 1 2670
box -10 -3 10 3
use M3_M2  M3_M2_3917
timestamp 1677677812
transform 1 0 84 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4442
timestamp 1677677812
transform 1 0 84 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4339
timestamp 1677677812
transform 1 0 108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4340
timestamp 1677677812
transform 1 0 124 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4034
timestamp 1677677812
transform 1 0 116 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4443
timestamp 1677677812
transform 1 0 148 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3918
timestamp 1677677812
transform 1 0 180 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4341
timestamp 1677677812
transform 1 0 164 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4342
timestamp 1677677812
transform 1 0 180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4444
timestamp 1677677812
transform 1 0 156 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4445
timestamp 1677677812
transform 1 0 164 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4446
timestamp 1677677812
transform 1 0 188 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4447
timestamp 1677677812
transform 1 0 196 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3999
timestamp 1677677812
transform 1 0 156 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4000
timestamp 1677677812
transform 1 0 188 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4035
timestamp 1677677812
transform 1 0 196 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3890
timestamp 1677677812
transform 1 0 324 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3912
timestamp 1677677812
transform 1 0 300 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3919
timestamp 1677677812
transform 1 0 300 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3920
timestamp 1677677812
transform 1 0 340 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4343
timestamp 1677677812
transform 1 0 300 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4344
timestamp 1677677812
transform 1 0 332 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4345
timestamp 1677677812
transform 1 0 340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4448
timestamp 1677677812
transform 1 0 252 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4036
timestamp 1677677812
transform 1 0 316 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3959
timestamp 1677677812
transform 1 0 348 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3921
timestamp 1677677812
transform 1 0 364 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4449
timestamp 1677677812
transform 1 0 372 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3922
timestamp 1677677812
transform 1 0 396 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4346
timestamp 1677677812
transform 1 0 468 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4347
timestamp 1677677812
transform 1 0 476 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3923
timestamp 1677677812
transform 1 0 492 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4348
timestamp 1677677812
transform 1 0 500 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3960
timestamp 1677677812
transform 1 0 508 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4349
timestamp 1677677812
transform 1 0 516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4450
timestamp 1677677812
transform 1 0 484 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4451
timestamp 1677677812
transform 1 0 492 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4452
timestamp 1677677812
transform 1 0 540 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4350
timestamp 1677677812
transform 1 0 572 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3961
timestamp 1677677812
transform 1 0 580 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3913
timestamp 1677677812
transform 1 0 596 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4351
timestamp 1677677812
transform 1 0 588 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4453
timestamp 1677677812
transform 1 0 564 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4001
timestamp 1677677812
transform 1 0 580 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4538
timestamp 1677677812
transform 1 0 596 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3924
timestamp 1677677812
transform 1 0 612 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4454
timestamp 1677677812
transform 1 0 612 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4002
timestamp 1677677812
transform 1 0 644 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4352
timestamp 1677677812
transform 1 0 740 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3881
timestamp 1677677812
transform 1 0 756 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4353
timestamp 1677677812
transform 1 0 756 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3925
timestamp 1677677812
transform 1 0 788 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4455
timestamp 1677677812
transform 1 0 788 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4456
timestamp 1677677812
transform 1 0 796 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4354
timestamp 1677677812
transform 1 0 828 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3914
timestamp 1677677812
transform 1 0 868 0 1 2635
box -3 -3 3 3
use M3_M2  M3_M2_3926
timestamp 1677677812
transform 1 0 892 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4355
timestamp 1677677812
transform 1 0 868 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4356
timestamp 1677677812
transform 1 0 884 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4357
timestamp 1677677812
transform 1 0 892 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4457
timestamp 1677677812
transform 1 0 852 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4458
timestamp 1677677812
transform 1 0 876 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4459
timestamp 1677677812
transform 1 0 884 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4003
timestamp 1677677812
transform 1 0 884 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3927
timestamp 1677677812
transform 1 0 932 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3928
timestamp 1677677812
transform 1 0 948 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4358
timestamp 1677677812
transform 1 0 940 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3962
timestamp 1677677812
transform 1 0 948 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4460
timestamp 1677677812
transform 1 0 948 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3963
timestamp 1677677812
transform 1 0 964 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3899
timestamp 1677677812
transform 1 0 996 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4359
timestamp 1677677812
transform 1 0 996 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3882
timestamp 1677677812
transform 1 0 1092 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3900
timestamp 1677677812
transform 1 0 1020 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3901
timestamp 1677677812
transform 1 0 1108 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3929
timestamp 1677677812
transform 1 0 1076 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3930
timestamp 1677677812
transform 1 0 1116 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3964
timestamp 1677677812
transform 1 0 1028 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4360
timestamp 1677677812
transform 1 0 1076 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4361
timestamp 1677677812
transform 1 0 1108 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4362
timestamp 1677677812
transform 1 0 1116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4461
timestamp 1677677812
transform 1 0 1028 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3987
timestamp 1677677812
transform 1 0 1076 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4462
timestamp 1677677812
transform 1 0 1116 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4004
timestamp 1677677812
transform 1 0 1044 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4005
timestamp 1677677812
transform 1 0 1108 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3902
timestamp 1677677812
transform 1 0 1140 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4539
timestamp 1677677812
transform 1 0 1132 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_3931
timestamp 1677677812
transform 1 0 1172 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4363
timestamp 1677677812
transform 1 0 1172 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4463
timestamp 1677677812
transform 1 0 1172 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4464
timestamp 1677677812
transform 1 0 1180 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4006
timestamp 1677677812
transform 1 0 1180 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4364
timestamp 1677677812
transform 1 0 1228 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3932
timestamp 1677677812
transform 1 0 1260 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4326
timestamp 1677677812
transform 1 0 1268 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4465
timestamp 1677677812
transform 1 0 1260 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4007
timestamp 1677677812
transform 1 0 1268 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4327
timestamp 1677677812
transform 1 0 1284 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3965
timestamp 1677677812
transform 1 0 1284 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4466
timestamp 1677677812
transform 1 0 1284 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3903
timestamp 1677677812
transform 1 0 1324 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4328
timestamp 1677677812
transform 1 0 1332 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3966
timestamp 1677677812
transform 1 0 1332 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4467
timestamp 1677677812
transform 1 0 1324 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4468
timestamp 1677677812
transform 1 0 1332 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4008
timestamp 1677677812
transform 1 0 1332 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3933
timestamp 1677677812
transform 1 0 1348 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4365
timestamp 1677677812
transform 1 0 1348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4329
timestamp 1677677812
transform 1 0 1380 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3934
timestamp 1677677812
transform 1 0 1396 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4366
timestamp 1677677812
transform 1 0 1396 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4367
timestamp 1677677812
transform 1 0 1420 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3935
timestamp 1677677812
transform 1 0 1492 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3936
timestamp 1677677812
transform 1 0 1516 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4368
timestamp 1677677812
transform 1 0 1516 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4469
timestamp 1677677812
transform 1 0 1564 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4470
timestamp 1677677812
transform 1 0 1580 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3904
timestamp 1677677812
transform 1 0 1612 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3905
timestamp 1677677812
transform 1 0 1636 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4369
timestamp 1677677812
transform 1 0 1612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4370
timestamp 1677677812
transform 1 0 1628 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4371
timestamp 1677677812
transform 1 0 1636 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4471
timestamp 1677677812
transform 1 0 1604 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4472
timestamp 1677677812
transform 1 0 1620 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4473
timestamp 1677677812
transform 1 0 1636 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4009
timestamp 1677677812
transform 1 0 1636 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4474
timestamp 1677677812
transform 1 0 1676 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4475
timestamp 1677677812
transform 1 0 1684 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3988
timestamp 1677677812
transform 1 0 1708 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4476
timestamp 1677677812
transform 1 0 1724 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4372
timestamp 1677677812
transform 1 0 1764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4373
timestamp 1677677812
transform 1 0 1788 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3891
timestamp 1677677812
transform 1 0 1828 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4374
timestamp 1677677812
transform 1 0 1812 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4477
timestamp 1677677812
transform 1 0 1804 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4037
timestamp 1677677812
transform 1 0 1804 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4478
timestamp 1677677812
transform 1 0 1828 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4479
timestamp 1677677812
transform 1 0 1868 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3937
timestamp 1677677812
transform 1 0 1892 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3906
timestamp 1677677812
transform 1 0 1948 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3938
timestamp 1677677812
transform 1 0 1932 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4375
timestamp 1677677812
transform 1 0 1892 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4376
timestamp 1677677812
transform 1 0 1900 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4377
timestamp 1677677812
transform 1 0 1932 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3967
timestamp 1677677812
transform 1 0 1980 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4480
timestamp 1677677812
transform 1 0 1980 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4038
timestamp 1677677812
transform 1 0 1988 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3892
timestamp 1677677812
transform 1 0 2116 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3939
timestamp 1677677812
transform 1 0 2020 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3940
timestamp 1677677812
transform 1 0 2060 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4378
timestamp 1677677812
transform 1 0 2020 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3968
timestamp 1677677812
transform 1 0 2036 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4379
timestamp 1677677812
transform 1 0 2060 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4380
timestamp 1677677812
transform 1 0 2116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4381
timestamp 1677677812
transform 1 0 2124 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4382
timestamp 1677677812
transform 1 0 2180 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4481
timestamp 1677677812
transform 1 0 2012 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4482
timestamp 1677677812
transform 1 0 2036 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4010
timestamp 1677677812
transform 1 0 2036 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4039
timestamp 1677677812
transform 1 0 2012 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3969
timestamp 1677677812
transform 1 0 2204 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4483
timestamp 1677677812
transform 1 0 2204 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3941
timestamp 1677677812
transform 1 0 2276 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3942
timestamp 1677677812
transform 1 0 2324 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4383
timestamp 1677677812
transform 1 0 2276 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4384
timestamp 1677677812
transform 1 0 2308 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4385
timestamp 1677677812
transform 1 0 2324 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4484
timestamp 1677677812
transform 1 0 2228 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4011
timestamp 1677677812
transform 1 0 2228 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4012
timestamp 1677677812
transform 1 0 2244 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4013
timestamp 1677677812
transform 1 0 2268 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4040
timestamp 1677677812
transform 1 0 2220 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4041
timestamp 1677677812
transform 1 0 2252 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4485
timestamp 1677677812
transform 1 0 2324 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4486
timestamp 1677677812
transform 1 0 2332 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4386
timestamp 1677677812
transform 1 0 2420 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4387
timestamp 1677677812
transform 1 0 2436 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4388
timestamp 1677677812
transform 1 0 2444 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4487
timestamp 1677677812
transform 1 0 2428 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4488
timestamp 1677677812
transform 1 0 2444 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4014
timestamp 1677677812
transform 1 0 2420 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4015
timestamp 1677677812
transform 1 0 2444 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4042
timestamp 1677677812
transform 1 0 2428 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4016
timestamp 1677677812
transform 1 0 2460 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4389
timestamp 1677677812
transform 1 0 2532 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3970
timestamp 1677677812
transform 1 0 2580 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4489
timestamp 1677677812
transform 1 0 2580 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4017
timestamp 1677677812
transform 1 0 2548 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4390
timestamp 1677677812
transform 1 0 2596 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4490
timestamp 1677677812
transform 1 0 2596 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4018
timestamp 1677677812
transform 1 0 2596 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3907
timestamp 1677677812
transform 1 0 2604 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4391
timestamp 1677677812
transform 1 0 2620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4392
timestamp 1677677812
transform 1 0 2628 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3989
timestamp 1677677812
transform 1 0 2620 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4393
timestamp 1677677812
transform 1 0 2684 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4394
timestamp 1677677812
transform 1 0 2700 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4491
timestamp 1677677812
transform 1 0 2668 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3990
timestamp 1677677812
transform 1 0 2700 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4019
timestamp 1677677812
transform 1 0 2668 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4020
timestamp 1677677812
transform 1 0 2684 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4540
timestamp 1677677812
transform 1 0 2708 0 1 2595
box -2 -2 2 2
use M3_M2  M3_M2_4043
timestamp 1677677812
transform 1 0 2708 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4492
timestamp 1677677812
transform 1 0 2748 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4044
timestamp 1677677812
transform 1 0 2748 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3893
timestamp 1677677812
transform 1 0 2764 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4493
timestamp 1677677812
transform 1 0 2764 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4494
timestamp 1677677812
transform 1 0 2772 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4021
timestamp 1677677812
transform 1 0 2764 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4045
timestamp 1677677812
transform 1 0 2796 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4395
timestamp 1677677812
transform 1 0 2820 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4396
timestamp 1677677812
transform 1 0 2828 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3991
timestamp 1677677812
transform 1 0 2820 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_4046
timestamp 1677677812
transform 1 0 2844 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3992
timestamp 1677677812
transform 1 0 2860 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4330
timestamp 1677677812
transform 1 0 2884 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3908
timestamp 1677677812
transform 1 0 2892 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4397
timestamp 1677677812
transform 1 0 2892 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4495
timestamp 1677677812
transform 1 0 2892 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4047
timestamp 1677677812
transform 1 0 2892 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4048
timestamp 1677677812
transform 1 0 2916 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4331
timestamp 1677677812
transform 1 0 2932 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4496
timestamp 1677677812
transform 1 0 2924 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4332
timestamp 1677677812
transform 1 0 2956 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3943
timestamp 1677677812
transform 1 0 2964 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3883
timestamp 1677677812
transform 1 0 2996 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4398
timestamp 1677677812
transform 1 0 2964 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3971
timestamp 1677677812
transform 1 0 2980 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4399
timestamp 1677677812
transform 1 0 2988 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3993
timestamp 1677677812
transform 1 0 2964 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3994
timestamp 1677677812
transform 1 0 2980 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4497
timestamp 1677677812
transform 1 0 2988 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3909
timestamp 1677677812
transform 1 0 3036 0 1 2645
box -3 -3 3 3
use M3_M2  M3_M2_3944
timestamp 1677677812
transform 1 0 3020 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4400
timestamp 1677677812
transform 1 0 3012 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4401
timestamp 1677677812
transform 1 0 3028 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4402
timestamp 1677677812
transform 1 0 3036 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4498
timestamp 1677677812
transform 1 0 3004 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3995
timestamp 1677677812
transform 1 0 3012 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4499
timestamp 1677677812
transform 1 0 3020 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4500
timestamp 1677677812
transform 1 0 3060 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4022
timestamp 1677677812
transform 1 0 3060 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3945
timestamp 1677677812
transform 1 0 3116 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4403
timestamp 1677677812
transform 1 0 3116 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4501
timestamp 1677677812
transform 1 0 3156 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3884
timestamp 1677677812
transform 1 0 3228 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3946
timestamp 1677677812
transform 1 0 3292 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3972
timestamp 1677677812
transform 1 0 3252 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4404
timestamp 1677677812
transform 1 0 3260 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4405
timestamp 1677677812
transform 1 0 3292 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4502
timestamp 1677677812
transform 1 0 3212 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4503
timestamp 1677677812
transform 1 0 3300 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4023
timestamp 1677677812
transform 1 0 3212 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3947
timestamp 1677677812
transform 1 0 3324 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4504
timestamp 1677677812
transform 1 0 3324 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3885
timestamp 1677677812
transform 1 0 3348 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4406
timestamp 1677677812
transform 1 0 3340 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4407
timestamp 1677677812
transform 1 0 3348 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4505
timestamp 1677677812
transform 1 0 3364 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4024
timestamp 1677677812
transform 1 0 3364 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4408
timestamp 1677677812
transform 1 0 3380 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3973
timestamp 1677677812
transform 1 0 3388 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4409
timestamp 1677677812
transform 1 0 3396 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4506
timestamp 1677677812
transform 1 0 3380 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4507
timestamp 1677677812
transform 1 0 3388 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4508
timestamp 1677677812
transform 1 0 3404 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4049
timestamp 1677677812
transform 1 0 3404 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4025
timestamp 1677677812
transform 1 0 3420 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4509
timestamp 1677677812
transform 1 0 3452 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3894
timestamp 1677677812
transform 1 0 3484 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3895
timestamp 1677677812
transform 1 0 3500 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4323
timestamp 1677677812
transform 1 0 3484 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4333
timestamp 1677677812
transform 1 0 3476 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3974
timestamp 1677677812
transform 1 0 3476 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4410
timestamp 1677677812
transform 1 0 3492 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3975
timestamp 1677677812
transform 1 0 3500 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3910
timestamp 1677677812
transform 1 0 3524 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4334
timestamp 1677677812
transform 1 0 3524 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3948
timestamp 1677677812
transform 1 0 3540 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3949
timestamp 1677677812
transform 1 0 3564 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4411
timestamp 1677677812
transform 1 0 3540 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4412
timestamp 1677677812
transform 1 0 3556 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4413
timestamp 1677677812
transform 1 0 3564 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4510
timestamp 1677677812
transform 1 0 3532 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4511
timestamp 1677677812
transform 1 0 3548 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4026
timestamp 1677677812
transform 1 0 3532 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4512
timestamp 1677677812
transform 1 0 3572 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4513
timestamp 1677677812
transform 1 0 3580 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4027
timestamp 1677677812
transform 1 0 3572 0 1 2595
box -3 -3 3 3
use M2_M1  M2_M1_4541
timestamp 1677677812
transform 1 0 3692 0 1 2585
box -2 -2 2 2
use M3_M2  M3_M2_3976
timestamp 1677677812
transform 1 0 3732 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3886
timestamp 1677677812
transform 1 0 3764 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3950
timestamp 1677677812
transform 1 0 3748 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4414
timestamp 1677677812
transform 1 0 3748 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3977
timestamp 1677677812
transform 1 0 3756 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4415
timestamp 1677677812
transform 1 0 3764 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4416
timestamp 1677677812
transform 1 0 3772 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4417
timestamp 1677677812
transform 1 0 3780 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4514
timestamp 1677677812
transform 1 0 3740 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4515
timestamp 1677677812
transform 1 0 3756 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4542
timestamp 1677677812
transform 1 0 3732 0 1 2585
box -2 -2 2 2
use M3_M2  M3_M2_3951
timestamp 1677677812
transform 1 0 3836 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4516
timestamp 1677677812
transform 1 0 3836 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3911
timestamp 1677677812
transform 1 0 3868 0 1 2645
box -3 -3 3 3
use M2_M1  M2_M1_4418
timestamp 1677677812
transform 1 0 3852 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3978
timestamp 1677677812
transform 1 0 3860 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4419
timestamp 1677677812
transform 1 0 3868 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4517
timestamp 1677677812
transform 1 0 3860 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4518
timestamp 1677677812
transform 1 0 3884 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3979
timestamp 1677677812
transform 1 0 3924 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4420
timestamp 1677677812
transform 1 0 3940 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3887
timestamp 1677677812
transform 1 0 3956 0 1 2665
box -3 -3 3 3
use M3_M2  M3_M2_3952
timestamp 1677677812
transform 1 0 3964 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4421
timestamp 1677677812
transform 1 0 3972 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3980
timestamp 1677677812
transform 1 0 3980 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4422
timestamp 1677677812
transform 1 0 3988 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4519
timestamp 1677677812
transform 1 0 3964 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4520
timestamp 1677677812
transform 1 0 3996 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4028
timestamp 1677677812
transform 1 0 3988 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4050
timestamp 1677677812
transform 1 0 3972 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4423
timestamp 1677677812
transform 1 0 4012 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4521
timestamp 1677677812
transform 1 0 4028 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4029
timestamp 1677677812
transform 1 0 4036 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3953
timestamp 1677677812
transform 1 0 4076 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4424
timestamp 1677677812
transform 1 0 4060 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4425
timestamp 1677677812
transform 1 0 4076 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4522
timestamp 1677677812
transform 1 0 4068 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3996
timestamp 1677677812
transform 1 0 4076 0 1 2605
box -3 -3 3 3
use M3_M2  M3_M2_3954
timestamp 1677677812
transform 1 0 4092 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4426
timestamp 1677677812
transform 1 0 4092 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4523
timestamp 1677677812
transform 1 0 4084 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4051
timestamp 1677677812
transform 1 0 4060 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_4030
timestamp 1677677812
transform 1 0 4116 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_4052
timestamp 1677677812
transform 1 0 4140 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3888
timestamp 1677677812
transform 1 0 4180 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4427
timestamp 1677677812
transform 1 0 4180 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3981
timestamp 1677677812
transform 1 0 4228 0 1 2615
box -3 -3 3 3
use M3_M2  M3_M2_3997
timestamp 1677677812
transform 1 0 4180 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4524
timestamp 1677677812
transform 1 0 4228 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4031
timestamp 1677677812
transform 1 0 4180 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3889
timestamp 1677677812
transform 1 0 4244 0 1 2665
box -3 -3 3 3
use M2_M1  M2_M1_4324
timestamp 1677677812
transform 1 0 4252 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4335
timestamp 1677677812
transform 1 0 4244 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3955
timestamp 1677677812
transform 1 0 4252 0 1 2625
box -3 -3 3 3
use M3_M2  M3_M2_3915
timestamp 1677677812
transform 1 0 4276 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4428
timestamp 1677677812
transform 1 0 4276 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_4053
timestamp 1677677812
transform 1 0 4276 0 1 2585
box -3 -3 3 3
use M2_M1  M2_M1_4336
timestamp 1677677812
transform 1 0 4308 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4525
timestamp 1677677812
transform 1 0 4308 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4054
timestamp 1677677812
transform 1 0 4308 0 1 2585
box -3 -3 3 3
use M3_M2  M3_M2_3896
timestamp 1677677812
transform 1 0 4348 0 1 2655
box -3 -3 3 3
use M3_M2  M3_M2_3916
timestamp 1677677812
transform 1 0 4340 0 1 2635
box -3 -3 3 3
use M2_M1  M2_M1_4325
timestamp 1677677812
transform 1 0 4348 0 1 2635
box -2 -2 2 2
use M2_M1  M2_M1_4337
timestamp 1677677812
transform 1 0 4340 0 1 2625
box -2 -2 2 2
use M2_M1  M2_M1_4429
timestamp 1677677812
transform 1 0 4332 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3956
timestamp 1677677812
transform 1 0 4356 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4430
timestamp 1677677812
transform 1 0 4356 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4526
timestamp 1677677812
transform 1 0 4372 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3897
timestamp 1677677812
transform 1 0 4404 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4338
timestamp 1677677812
transform 1 0 4404 0 1 2625
box -2 -2 2 2
use M3_M2  M3_M2_3898
timestamp 1677677812
transform 1 0 4452 0 1 2655
box -3 -3 3 3
use M2_M1  M2_M1_4431
timestamp 1677677812
transform 1 0 4412 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4432
timestamp 1677677812
transform 1 0 4436 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3982
timestamp 1677677812
transform 1 0 4444 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4527
timestamp 1677677812
transform 1 0 4428 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4528
timestamp 1677677812
transform 1 0 4452 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4433
timestamp 1677677812
transform 1 0 4468 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3983
timestamp 1677677812
transform 1 0 4492 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4529
timestamp 1677677812
transform 1 0 4492 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3984
timestamp 1677677812
transform 1 0 4564 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4434
timestamp 1677677812
transform 1 0 4572 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3985
timestamp 1677677812
transform 1 0 4596 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4530
timestamp 1677677812
transform 1 0 4524 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_3957
timestamp 1677677812
transform 1 0 4636 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4435
timestamp 1677677812
transform 1 0 4612 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4436
timestamp 1677677812
transform 1 0 4620 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4437
timestamp 1677677812
transform 1 0 4636 0 1 2615
box -2 -2 2 2
use M3_M2  M3_M2_3986
timestamp 1677677812
transform 1 0 4644 0 1 2615
box -3 -3 3 3
use M2_M1  M2_M1_4438
timestamp 1677677812
transform 1 0 4652 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4439
timestamp 1677677812
transform 1 0 4660 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4531
timestamp 1677677812
transform 1 0 4628 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4532
timestamp 1677677812
transform 1 0 4644 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4533
timestamp 1677677812
transform 1 0 4652 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4032
timestamp 1677677812
transform 1 0 4628 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3958
timestamp 1677677812
transform 1 0 4692 0 1 2625
box -3 -3 3 3
use M2_M1  M2_M1_4440
timestamp 1677677812
transform 1 0 4692 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4441
timestamp 1677677812
transform 1 0 4708 0 1 2615
box -2 -2 2 2
use M2_M1  M2_M1_4534
timestamp 1677677812
transform 1 0 4668 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4535
timestamp 1677677812
transform 1 0 4684 0 1 2605
box -2 -2 2 2
use M2_M1  M2_M1_4536
timestamp 1677677812
transform 1 0 4700 0 1 2605
box -2 -2 2 2
use M3_M2  M3_M2_4033
timestamp 1677677812
transform 1 0 4692 0 1 2595
box -3 -3 3 3
use M3_M2  M3_M2_3998
timestamp 1677677812
transform 1 0 4708 0 1 2605
box -3 -3 3 3
use M2_M1  M2_M1_4537
timestamp 1677677812
transform 1 0 4788 0 1 2605
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_42
timestamp 1677677812
transform 1 0 48 0 1 2570
box -10 -3 10 3
use FILL  FILL_4837
timestamp 1677677812
transform 1 0 72 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_329
timestamp 1677677812
transform 1 0 80 0 1 2570
box -9 -3 26 105
use FILL  FILL_4838
timestamp 1677677812
transform 1 0 96 0 1 2570
box -8 -3 16 105
use FILL  FILL_4839
timestamp 1677677812
transform 1 0 104 0 1 2570
box -8 -3 16 105
use FILL  FILL_4840
timestamp 1677677812
transform 1 0 112 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_330
timestamp 1677677812
transform -1 0 136 0 1 2570
box -9 -3 26 105
use FILL  FILL_4841
timestamp 1677677812
transform 1 0 136 0 1 2570
box -8 -3 16 105
use FILL  FILL_4842
timestamp 1677677812
transform 1 0 144 0 1 2570
box -8 -3 16 105
use FILL  FILL_4843
timestamp 1677677812
transform 1 0 152 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_200
timestamp 1677677812
transform -1 0 200 0 1 2570
box -8 -3 46 105
use FILL  FILL_4844
timestamp 1677677812
transform 1 0 200 0 1 2570
box -8 -3 16 105
use FILL  FILL_4845
timestamp 1677677812
transform 1 0 208 0 1 2570
box -8 -3 16 105
use FILL  FILL_4846
timestamp 1677677812
transform 1 0 216 0 1 2570
box -8 -3 16 105
use FILL  FILL_4847
timestamp 1677677812
transform 1 0 224 0 1 2570
box -8 -3 16 105
use FILL  FILL_4848
timestamp 1677677812
transform 1 0 232 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_293
timestamp 1677677812
transform 1 0 240 0 1 2570
box -8 -3 104 105
use FILL  FILL_4849
timestamp 1677677812
transform 1 0 336 0 1 2570
box -8 -3 16 105
use FILL  FILL_4858
timestamp 1677677812
transform 1 0 344 0 1 2570
box -8 -3 16 105
use FILL  FILL_4859
timestamp 1677677812
transform 1 0 352 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_332
timestamp 1677677812
transform -1 0 376 0 1 2570
box -9 -3 26 105
use FILL  FILL_4860
timestamp 1677677812
transform 1 0 376 0 1 2570
box -8 -3 16 105
use FILL  FILL_4861
timestamp 1677677812
transform 1 0 384 0 1 2570
box -8 -3 16 105
use FILL  FILL_4862
timestamp 1677677812
transform 1 0 392 0 1 2570
box -8 -3 16 105
use FILL  FILL_4865
timestamp 1677677812
transform 1 0 400 0 1 2570
box -8 -3 16 105
use FILL  FILL_4867
timestamp 1677677812
transform 1 0 408 0 1 2570
box -8 -3 16 105
use FILL  FILL_4869
timestamp 1677677812
transform 1 0 416 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4055
timestamp 1677677812
transform 1 0 444 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_333
timestamp 1677677812
transform -1 0 440 0 1 2570
box -9 -3 26 105
use FILL  FILL_4870
timestamp 1677677812
transform 1 0 440 0 1 2570
box -8 -3 16 105
use FILL  FILL_4875
timestamp 1677677812
transform 1 0 448 0 1 2570
box -8 -3 16 105
use FILL  FILL_4877
timestamp 1677677812
transform 1 0 456 0 1 2570
box -8 -3 16 105
use FILL  FILL_4879
timestamp 1677677812
transform 1 0 464 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4056
timestamp 1677677812
transform 1 0 484 0 1 2575
box -3 -3 3 3
use FILL  FILL_4881
timestamp 1677677812
transform 1 0 472 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_202
timestamp 1677677812
transform 1 0 480 0 1 2570
box -8 -3 46 105
use FILL  FILL_4882
timestamp 1677677812
transform 1 0 520 0 1 2570
box -8 -3 16 105
use FILL  FILL_4883
timestamp 1677677812
transform 1 0 528 0 1 2570
box -8 -3 16 105
use FILL  FILL_4884
timestamp 1677677812
transform 1 0 536 0 1 2570
box -8 -3 16 105
use FILL  FILL_4885
timestamp 1677677812
transform 1 0 544 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_203
timestamp 1677677812
transform -1 0 592 0 1 2570
box -8 -3 46 105
use FILL  FILL_4886
timestamp 1677677812
transform 1 0 592 0 1 2570
box -8 -3 16 105
use FILL  FILL_4887
timestamp 1677677812
transform 1 0 600 0 1 2570
box -8 -3 16 105
use FILL  FILL_4888
timestamp 1677677812
transform 1 0 608 0 1 2570
box -8 -3 16 105
use FILL  FILL_4893
timestamp 1677677812
transform 1 0 616 0 1 2570
box -8 -3 16 105
use FILL  FILL_4895
timestamp 1677677812
transform 1 0 624 0 1 2570
box -8 -3 16 105
use FILL  FILL_4897
timestamp 1677677812
transform 1 0 632 0 1 2570
box -8 -3 16 105
use FILL  FILL_4899
timestamp 1677677812
transform 1 0 640 0 1 2570
box -8 -3 16 105
use FILL  FILL_4900
timestamp 1677677812
transform 1 0 648 0 1 2570
box -8 -3 16 105
use FILL  FILL_4901
timestamp 1677677812
transform 1 0 656 0 1 2570
box -8 -3 16 105
use FILL  FILL_4902
timestamp 1677677812
transform 1 0 664 0 1 2570
box -8 -3 16 105
use FILL  FILL_4903
timestamp 1677677812
transform 1 0 672 0 1 2570
box -8 -3 16 105
use FILL  FILL_4904
timestamp 1677677812
transform 1 0 680 0 1 2570
box -8 -3 16 105
use FILL  FILL_4906
timestamp 1677677812
transform 1 0 688 0 1 2570
box -8 -3 16 105
use FILL  FILL_4908
timestamp 1677677812
transform 1 0 696 0 1 2570
box -8 -3 16 105
use FILL  FILL_4910
timestamp 1677677812
transform 1 0 704 0 1 2570
box -8 -3 16 105
use FILL  FILL_4912
timestamp 1677677812
transform 1 0 712 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_49
timestamp 1677677812
transform 1 0 720 0 1 2570
box -8 -3 32 105
use FILL  FILL_4914
timestamp 1677677812
transform 1 0 744 0 1 2570
box -8 -3 16 105
use FILL  FILL_4917
timestamp 1677677812
transform 1 0 752 0 1 2570
box -8 -3 16 105
use FILL  FILL_4919
timestamp 1677677812
transform 1 0 760 0 1 2570
box -8 -3 16 105
use FILL  FILL_4921
timestamp 1677677812
transform 1 0 768 0 1 2570
box -8 -3 16 105
use FILL  FILL_4923
timestamp 1677677812
transform 1 0 776 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4057
timestamp 1677677812
transform 1 0 796 0 1 2575
box -3 -3 3 3
use FILL  FILL_4925
timestamp 1677677812
transform 1 0 784 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_336
timestamp 1677677812
transform 1 0 792 0 1 2570
box -9 -3 26 105
use FILL  FILL_4927
timestamp 1677677812
transform 1 0 808 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4058
timestamp 1677677812
transform 1 0 828 0 1 2575
box -3 -3 3 3
use FILL  FILL_4928
timestamp 1677677812
transform 1 0 816 0 1 2570
box -8 -3 16 105
use FILL  FILL_4929
timestamp 1677677812
transform 1 0 824 0 1 2570
box -8 -3 16 105
use FILL  FILL_4930
timestamp 1677677812
transform 1 0 832 0 1 2570
box -8 -3 16 105
use FILL  FILL_4931
timestamp 1677677812
transform 1 0 840 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4059
timestamp 1677677812
transform 1 0 884 0 1 2575
box -3 -3 3 3
use AOI22X1  AOI22X1_205
timestamp 1677677812
transform 1 0 848 0 1 2570
box -8 -3 46 105
use FILL  FILL_4934
timestamp 1677677812
transform 1 0 888 0 1 2570
box -8 -3 16 105
use FILL  FILL_4941
timestamp 1677677812
transform 1 0 896 0 1 2570
box -8 -3 16 105
use FILL  FILL_4942
timestamp 1677677812
transform 1 0 904 0 1 2570
box -8 -3 16 105
use FILL  FILL_4943
timestamp 1677677812
transform 1 0 912 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4060
timestamp 1677677812
transform 1 0 948 0 1 2575
box -3 -3 3 3
use AOI22X1  AOI22X1_206
timestamp 1677677812
transform 1 0 920 0 1 2570
box -8 -3 46 105
use FILL  FILL_4944
timestamp 1677677812
transform 1 0 960 0 1 2570
box -8 -3 16 105
use FILL  FILL_4949
timestamp 1677677812
transform 1 0 968 0 1 2570
box -8 -3 16 105
use FILL  FILL_4951
timestamp 1677677812
transform 1 0 976 0 1 2570
box -8 -3 16 105
use FILL  FILL_4953
timestamp 1677677812
transform 1 0 984 0 1 2570
box -8 -3 16 105
use FILL  FILL_4955
timestamp 1677677812
transform 1 0 992 0 1 2570
box -8 -3 16 105
use FILL  FILL_4957
timestamp 1677677812
transform 1 0 1000 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4061
timestamp 1677677812
transform 1 0 1020 0 1 2575
box -3 -3 3 3
use FILL  FILL_4958
timestamp 1677677812
transform 1 0 1008 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_297
timestamp 1677677812
transform 1 0 1016 0 1 2570
box -8 -3 104 105
use INVX2  INVX2_337
timestamp 1677677812
transform 1 0 1112 0 1 2570
box -9 -3 26 105
use FILL  FILL_4959
timestamp 1677677812
transform 1 0 1128 0 1 2570
box -8 -3 16 105
use FILL  FILL_4969
timestamp 1677677812
transform 1 0 1136 0 1 2570
box -8 -3 16 105
use FILL  FILL_4971
timestamp 1677677812
transform 1 0 1144 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_51
timestamp 1677677812
transform 1 0 1152 0 1 2570
box -8 -3 32 105
use FILL  FILL_4973
timestamp 1677677812
transform 1 0 1176 0 1 2570
box -8 -3 16 105
use FILL  FILL_4974
timestamp 1677677812
transform 1 0 1184 0 1 2570
box -8 -3 16 105
use FILL  FILL_4975
timestamp 1677677812
transform 1 0 1192 0 1 2570
box -8 -3 16 105
use FILL  FILL_4976
timestamp 1677677812
transform 1 0 1200 0 1 2570
box -8 -3 16 105
use FILL  FILL_4977
timestamp 1677677812
transform 1 0 1208 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_100
timestamp 1677677812
transform 1 0 1216 0 1 2570
box -8 -3 34 105
use FILL  FILL_4978
timestamp 1677677812
transform 1 0 1248 0 1 2570
box -8 -3 16 105
use FILL  FILL_4987
timestamp 1677677812
transform 1 0 1256 0 1 2570
box -8 -3 16 105
use FILL  FILL_4989
timestamp 1677677812
transform 1 0 1264 0 1 2570
box -8 -3 16 105
use FILL  FILL_4991
timestamp 1677677812
transform 1 0 1272 0 1 2570
box -8 -3 16 105
use FILL  FILL_4992
timestamp 1677677812
transform 1 0 1280 0 1 2570
box -8 -3 16 105
use FILL  FILL_4993
timestamp 1677677812
transform 1 0 1288 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_101
timestamp 1677677812
transform -1 0 1328 0 1 2570
box -8 -3 34 105
use FILL  FILL_4994
timestamp 1677677812
transform 1 0 1328 0 1 2570
box -8 -3 16 105
use FILL  FILL_4999
timestamp 1677677812
transform 1 0 1336 0 1 2570
box -8 -3 16 105
use FILL  FILL_5001
timestamp 1677677812
transform 1 0 1344 0 1 2570
box -8 -3 16 105
use FILL  FILL_5002
timestamp 1677677812
transform 1 0 1352 0 1 2570
box -8 -3 16 105
use FILL  FILL_5003
timestamp 1677677812
transform 1 0 1360 0 1 2570
box -8 -3 16 105
use FILL  FILL_5004
timestamp 1677677812
transform 1 0 1368 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_103
timestamp 1677677812
transform -1 0 1408 0 1 2570
box -8 -3 34 105
use FILL  FILL_5005
timestamp 1677677812
transform 1 0 1408 0 1 2570
box -8 -3 16 105
use FILL  FILL_5010
timestamp 1677677812
transform 1 0 1416 0 1 2570
box -8 -3 16 105
use FILL  FILL_5012
timestamp 1677677812
transform 1 0 1424 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_339
timestamp 1677677812
transform -1 0 1448 0 1 2570
box -9 -3 26 105
use FILL  FILL_5013
timestamp 1677677812
transform 1 0 1448 0 1 2570
box -8 -3 16 105
use FILL  FILL_5014
timestamp 1677677812
transform 1 0 1456 0 1 2570
box -8 -3 16 105
use FILL  FILL_5018
timestamp 1677677812
transform 1 0 1464 0 1 2570
box -8 -3 16 105
use FILL  FILL_5020
timestamp 1677677812
transform 1 0 1472 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_298
timestamp 1677677812
transform -1 0 1576 0 1 2570
box -8 -3 104 105
use FILL  FILL_5021
timestamp 1677677812
transform 1 0 1576 0 1 2570
box -8 -3 16 105
use FILL  FILL_5022
timestamp 1677677812
transform 1 0 1584 0 1 2570
box -8 -3 16 105
use FILL  FILL_5026
timestamp 1677677812
transform 1 0 1592 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4062
timestamp 1677677812
transform 1 0 1612 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_196
timestamp 1677677812
transform -1 0 1640 0 1 2570
box -8 -3 46 105
use FILL  FILL_5027
timestamp 1677677812
transform 1 0 1640 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_341
timestamp 1677677812
transform -1 0 1664 0 1 2570
box -9 -3 26 105
use FILL  FILL_5028
timestamp 1677677812
transform 1 0 1664 0 1 2570
box -8 -3 16 105
use FILL  FILL_5037
timestamp 1677677812
transform 1 0 1672 0 1 2570
box -8 -3 16 105
use FILL  FILL_5038
timestamp 1677677812
transform 1 0 1680 0 1 2570
box -8 -3 16 105
use FILL  FILL_5039
timestamp 1677677812
transform 1 0 1688 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4063
timestamp 1677677812
transform 1 0 1708 0 1 2575
box -3 -3 3 3
use FILL  FILL_5040
timestamp 1677677812
transform 1 0 1696 0 1 2570
box -8 -3 16 105
use FILL  FILL_5041
timestamp 1677677812
transform 1 0 1704 0 1 2570
box -8 -3 16 105
use FILL  FILL_5042
timestamp 1677677812
transform 1 0 1712 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_35
timestamp 1677677812
transform -1 0 1744 0 1 2570
box -5 -3 28 105
use FILL  FILL_5043
timestamp 1677677812
transform 1 0 1744 0 1 2570
box -8 -3 16 105
use FILL  FILL_5044
timestamp 1677677812
transform 1 0 1752 0 1 2570
box -8 -3 16 105
use FILL  FILL_5045
timestamp 1677677812
transform 1 0 1760 0 1 2570
box -8 -3 16 105
use FILL  FILL_5046
timestamp 1677677812
transform 1 0 1768 0 1 2570
box -8 -3 16 105
use FILL  FILL_5047
timestamp 1677677812
transform 1 0 1776 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_36
timestamp 1677677812
transform 1 0 1784 0 1 2570
box -5 -3 28 105
use BUFX2  BUFX2_37
timestamp 1677677812
transform 1 0 1808 0 1 2570
box -5 -3 28 105
use FILL  FILL_5050
timestamp 1677677812
transform 1 0 1832 0 1 2570
box -8 -3 16 105
use FILL  FILL_5055
timestamp 1677677812
transform 1 0 1840 0 1 2570
box -8 -3 16 105
use FILL  FILL_5057
timestamp 1677677812
transform 1 0 1848 0 1 2570
box -8 -3 16 105
use FILL  FILL_5059
timestamp 1677677812
transform 1 0 1856 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_343
timestamp 1677677812
transform 1 0 1864 0 1 2570
box -9 -3 26 105
use FILL  FILL_5061
timestamp 1677677812
transform 1 0 1880 0 1 2570
box -8 -3 16 105
use FILL  FILL_5062
timestamp 1677677812
transform 1 0 1888 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_301
timestamp 1677677812
transform -1 0 1992 0 1 2570
box -8 -3 104 105
use FILL  FILL_5063
timestamp 1677677812
transform 1 0 1992 0 1 2570
box -8 -3 16 105
use FILL  FILL_5064
timestamp 1677677812
transform 1 0 2000 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_344
timestamp 1677677812
transform 1 0 2008 0 1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_302
timestamp 1677677812
transform 1 0 2024 0 1 2570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_303
timestamp 1677677812
transform -1 0 2216 0 1 2570
box -8 -3 104 105
use M3_M2  M3_M2_4064
timestamp 1677677812
transform 1 0 2308 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_304
timestamp 1677677812
transform 1 0 2216 0 1 2570
box -8 -3 104 105
use M3_M2  M3_M2_4065
timestamp 1677677812
transform 1 0 2332 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_345
timestamp 1677677812
transform -1 0 2328 0 1 2570
box -9 -3 26 105
use FILL  FILL_5065
timestamp 1677677812
transform 1 0 2328 0 1 2570
box -8 -3 16 105
use FILL  FILL_5066
timestamp 1677677812
transform 1 0 2336 0 1 2570
box -8 -3 16 105
use FILL  FILL_5067
timestamp 1677677812
transform 1 0 2344 0 1 2570
box -8 -3 16 105
use FILL  FILL_5107
timestamp 1677677812
transform 1 0 2352 0 1 2570
box -8 -3 16 105
use FILL  FILL_5109
timestamp 1677677812
transform 1 0 2360 0 1 2570
box -8 -3 16 105
use FILL  FILL_5111
timestamp 1677677812
transform 1 0 2368 0 1 2570
box -8 -3 16 105
use FILL  FILL_5113
timestamp 1677677812
transform 1 0 2376 0 1 2570
box -8 -3 16 105
use FILL  FILL_5115
timestamp 1677677812
transform 1 0 2384 0 1 2570
box -8 -3 16 105
use FILL  FILL_5117
timestamp 1677677812
transform 1 0 2392 0 1 2570
box -8 -3 16 105
use FILL  FILL_5119
timestamp 1677677812
transform 1 0 2400 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_197
timestamp 1677677812
transform -1 0 2448 0 1 2570
box -8 -3 46 105
use FILL  FILL_5120
timestamp 1677677812
transform 1 0 2448 0 1 2570
box -8 -3 16 105
use FILL  FILL_5121
timestamp 1677677812
transform 1 0 2456 0 1 2570
box -8 -3 16 105
use FILL  FILL_5125
timestamp 1677677812
transform 1 0 2464 0 1 2570
box -8 -3 16 105
use FILL  FILL_5127
timestamp 1677677812
transform 1 0 2472 0 1 2570
box -8 -3 16 105
use FILL  FILL_5129
timestamp 1677677812
transform 1 0 2480 0 1 2570
box -8 -3 16 105
use FILL  FILL_5131
timestamp 1677677812
transform 1 0 2488 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4066
timestamp 1677677812
transform 1 0 2580 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_305
timestamp 1677677812
transform -1 0 2592 0 1 2570
box -8 -3 104 105
use FILL  FILL_5132
timestamp 1677677812
transform 1 0 2592 0 1 2570
box -8 -3 16 105
use FILL  FILL_5142
timestamp 1677677812
transform 1 0 2600 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_348
timestamp 1677677812
transform 1 0 2608 0 1 2570
box -9 -3 26 105
use FILL  FILL_5144
timestamp 1677677812
transform 1 0 2624 0 1 2570
box -8 -3 16 105
use FILL  FILL_5145
timestamp 1677677812
transform 1 0 2632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5148
timestamp 1677677812
transform 1 0 2640 0 1 2570
box -8 -3 16 105
use FILL  FILL_5150
timestamp 1677677812
transform 1 0 2648 0 1 2570
box -8 -3 16 105
use FILL  FILL_5152
timestamp 1677677812
transform 1 0 2656 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_214
timestamp 1677677812
transform 1 0 2664 0 1 2570
box -8 -3 46 105
use FILL  FILL_5154
timestamp 1677677812
transform 1 0 2704 0 1 2570
box -8 -3 16 105
use FILL  FILL_5155
timestamp 1677677812
transform 1 0 2712 0 1 2570
box -8 -3 16 105
use FILL  FILL_5156
timestamp 1677677812
transform 1 0 2720 0 1 2570
box -8 -3 16 105
use FILL  FILL_5157
timestamp 1677677812
transform 1 0 2728 0 1 2570
box -8 -3 16 105
use FILL  FILL_5158
timestamp 1677677812
transform 1 0 2736 0 1 2570
box -8 -3 16 105
use FILL  FILL_5159
timestamp 1677677812
transform 1 0 2744 0 1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_52
timestamp 1677677812
transform 1 0 2752 0 1 2570
box -8 -3 32 105
use FILL  FILL_5160
timestamp 1677677812
transform 1 0 2776 0 1 2570
box -8 -3 16 105
use FILL  FILL_5162
timestamp 1677677812
transform 1 0 2784 0 1 2570
box -8 -3 16 105
use FILL  FILL_5164
timestamp 1677677812
transform 1 0 2792 0 1 2570
box -8 -3 16 105
use FILL  FILL_5166
timestamp 1677677812
transform 1 0 2800 0 1 2570
box -8 -3 16 105
use FILL  FILL_5168
timestamp 1677677812
transform 1 0 2808 0 1 2570
box -8 -3 16 105
use FILL  FILL_5170
timestamp 1677677812
transform 1 0 2816 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_104
timestamp 1677677812
transform 1 0 2824 0 1 2570
box -8 -3 34 105
use FILL  FILL_5172
timestamp 1677677812
transform 1 0 2856 0 1 2570
box -8 -3 16 105
use FILL  FILL_5173
timestamp 1677677812
transform 1 0 2864 0 1 2570
box -8 -3 16 105
use FILL  FILL_5176
timestamp 1677677812
transform 1 0 2872 0 1 2570
box -8 -3 16 105
use FILL  FILL_5178
timestamp 1677677812
transform 1 0 2880 0 1 2570
box -8 -3 16 105
use FILL  FILL_5180
timestamp 1677677812
transform 1 0 2888 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_351
timestamp 1677677812
transform 1 0 2896 0 1 2570
box -9 -3 26 105
use FILL  FILL_5182
timestamp 1677677812
transform 1 0 2912 0 1 2570
box -8 -3 16 105
use FILL  FILL_5183
timestamp 1677677812
transform 1 0 2920 0 1 2570
box -8 -3 16 105
use FILL  FILL_5185
timestamp 1677677812
transform 1 0 2928 0 1 2570
box -8 -3 16 105
use FILL  FILL_5187
timestamp 1677677812
transform 1 0 2936 0 1 2570
box -8 -3 16 105
use FILL  FILL_5189
timestamp 1677677812
transform 1 0 2944 0 1 2570
box -8 -3 16 105
use FILL  FILL_5190
timestamp 1677677812
transform 1 0 2952 0 1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_106
timestamp 1677677812
transform -1 0 2992 0 1 2570
box -8 -3 34 105
use FILL  FILL_5191
timestamp 1677677812
transform 1 0 2992 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_199
timestamp 1677677812
transform -1 0 3040 0 1 2570
box -8 -3 46 105
use FILL  FILL_5192
timestamp 1677677812
transform 1 0 3040 0 1 2570
box -8 -3 16 105
use FILL  FILL_5199
timestamp 1677677812
transform 1 0 3048 0 1 2570
box -8 -3 16 105
use FILL  FILL_5200
timestamp 1677677812
transform 1 0 3056 0 1 2570
box -8 -3 16 105
use FILL  FILL_5201
timestamp 1677677812
transform 1 0 3064 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_307
timestamp 1677677812
transform -1 0 3168 0 1 2570
box -8 -3 104 105
use FILL  FILL_5202
timestamp 1677677812
transform 1 0 3168 0 1 2570
box -8 -3 16 105
use FILL  FILL_5203
timestamp 1677677812
transform 1 0 3176 0 1 2570
box -8 -3 16 105
use FILL  FILL_5204
timestamp 1677677812
transform 1 0 3184 0 1 2570
box -8 -3 16 105
use FILL  FILL_5208
timestamp 1677677812
transform 1 0 3192 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4067
timestamp 1677677812
transform 1 0 3228 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_309
timestamp 1677677812
transform 1 0 3200 0 1 2570
box -8 -3 104 105
use BUFX2  BUFX2_42
timestamp 1677677812
transform -1 0 3320 0 1 2570
box -5 -3 28 105
use FILL  FILL_5209
timestamp 1677677812
transform 1 0 3320 0 1 2570
box -8 -3 16 105
use FILL  FILL_5210
timestamp 1677677812
transform 1 0 3328 0 1 2570
box -8 -3 16 105
use FILL  FILL_5211
timestamp 1677677812
transform 1 0 3336 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_352
timestamp 1677677812
transform 1 0 3344 0 1 2570
box -9 -3 26 105
use FILL  FILL_5212
timestamp 1677677812
transform 1 0 3360 0 1 2570
box -8 -3 16 105
use FILL  FILL_5225
timestamp 1677677812
transform 1 0 3368 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_215
timestamp 1677677812
transform -1 0 3416 0 1 2570
box -8 -3 46 105
use FILL  FILL_5226
timestamp 1677677812
transform 1 0 3416 0 1 2570
box -8 -3 16 105
use FILL  FILL_5230
timestamp 1677677812
transform 1 0 3424 0 1 2570
box -8 -3 16 105
use FILL  FILL_5232
timestamp 1677677812
transform 1 0 3432 0 1 2570
box -8 -3 16 105
use FILL  FILL_5233
timestamp 1677677812
transform 1 0 3440 0 1 2570
box -8 -3 16 105
use FILL  FILL_5234
timestamp 1677677812
transform 1 0 3448 0 1 2570
box -8 -3 16 105
use FILL  FILL_5235
timestamp 1677677812
transform 1 0 3456 0 1 2570
box -8 -3 16 105
use FILL  FILL_5237
timestamp 1677677812
transform 1 0 3464 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_30
timestamp 1677677812
transform -1 0 3504 0 1 2570
box -8 -3 40 105
use FILL  FILL_5238
timestamp 1677677812
transform 1 0 3504 0 1 2570
box -8 -3 16 105
use FILL  FILL_5239
timestamp 1677677812
transform 1 0 3512 0 1 2570
box -8 -3 16 105
use FILL  FILL_5243
timestamp 1677677812
transform 1 0 3520 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_200
timestamp 1677677812
transform -1 0 3568 0 1 2570
box -8 -3 46 105
use FILL  FILL_5244
timestamp 1677677812
transform 1 0 3568 0 1 2570
box -8 -3 16 105
use FILL  FILL_5245
timestamp 1677677812
transform 1 0 3576 0 1 2570
box -8 -3 16 105
use FILL  FILL_5249
timestamp 1677677812
transform 1 0 3584 0 1 2570
box -8 -3 16 105
use FILL  FILL_5251
timestamp 1677677812
transform 1 0 3592 0 1 2570
box -8 -3 16 105
use FILL  FILL_5253
timestamp 1677677812
transform 1 0 3600 0 1 2570
box -8 -3 16 105
use FILL  FILL_5254
timestamp 1677677812
transform 1 0 3608 0 1 2570
box -8 -3 16 105
use FILL  FILL_5255
timestamp 1677677812
transform 1 0 3616 0 1 2570
box -8 -3 16 105
use FILL  FILL_5257
timestamp 1677677812
transform 1 0 3624 0 1 2570
box -8 -3 16 105
use FILL  FILL_5259
timestamp 1677677812
transform 1 0 3632 0 1 2570
box -8 -3 16 105
use FILL  FILL_5261
timestamp 1677677812
transform 1 0 3640 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_354
timestamp 1677677812
transform 1 0 3648 0 1 2570
box -9 -3 26 105
use FILL  FILL_5263
timestamp 1677677812
transform 1 0 3664 0 1 2570
box -8 -3 16 105
use FILL  FILL_5264
timestamp 1677677812
transform 1 0 3672 0 1 2570
box -8 -3 16 105
use FILL  FILL_5267
timestamp 1677677812
transform 1 0 3680 0 1 2570
box -8 -3 16 105
use FILL  FILL_5269
timestamp 1677677812
transform 1 0 3688 0 1 2570
box -8 -3 16 105
use FILL  FILL_5271
timestamp 1677677812
transform 1 0 3696 0 1 2570
box -8 -3 16 105
use FILL  FILL_5272
timestamp 1677677812
transform 1 0 3704 0 1 2570
box -8 -3 16 105
use FILL  FILL_5273
timestamp 1677677812
transform 1 0 3712 0 1 2570
box -8 -3 16 105
use FILL  FILL_5274
timestamp 1677677812
transform 1 0 3720 0 1 2570
box -8 -3 16 105
use FILL  FILL_5275
timestamp 1677677812
transform 1 0 3728 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_202
timestamp 1677677812
transform -1 0 3776 0 1 2570
box -8 -3 46 105
use FILL  FILL_5276
timestamp 1677677812
transform 1 0 3776 0 1 2570
box -8 -3 16 105
use FILL  FILL_5277
timestamp 1677677812
transform 1 0 3784 0 1 2570
box -8 -3 16 105
use FILL  FILL_5278
timestamp 1677677812
transform 1 0 3792 0 1 2570
box -8 -3 16 105
use FILL  FILL_5279
timestamp 1677677812
transform 1 0 3800 0 1 2570
box -8 -3 16 105
use FILL  FILL_5280
timestamp 1677677812
transform 1 0 3808 0 1 2570
box -8 -3 16 105
use FILL  FILL_5281
timestamp 1677677812
transform 1 0 3816 0 1 2570
box -8 -3 16 105
use FILL  FILL_5282
timestamp 1677677812
transform 1 0 3824 0 1 2570
box -8 -3 16 105
use FILL  FILL_5283
timestamp 1677677812
transform 1 0 3832 0 1 2570
box -8 -3 16 105
use FILL  FILL_5284
timestamp 1677677812
transform 1 0 3840 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_216
timestamp 1677677812
transform -1 0 3888 0 1 2570
box -8 -3 46 105
use FILL  FILL_5285
timestamp 1677677812
transform 1 0 3888 0 1 2570
box -8 -3 16 105
use FILL  FILL_5286
timestamp 1677677812
transform 1 0 3896 0 1 2570
box -8 -3 16 105
use FILL  FILL_5287
timestamp 1677677812
transform 1 0 3904 0 1 2570
box -8 -3 16 105
use FILL  FILL_5288
timestamp 1677677812
transform 1 0 3912 0 1 2570
box -8 -3 16 105
use FILL  FILL_5289
timestamp 1677677812
transform 1 0 3920 0 1 2570
box -8 -3 16 105
use FILL  FILL_5294
timestamp 1677677812
transform 1 0 3928 0 1 2570
box -8 -3 16 105
use FILL  FILL_5296
timestamp 1677677812
transform 1 0 3936 0 1 2570
box -8 -3 16 105
use FILL  FILL_5298
timestamp 1677677812
transform 1 0 3944 0 1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_218
timestamp 1677677812
transform 1 0 3952 0 1 2570
box -8 -3 46 105
use FILL  FILL_5300
timestamp 1677677812
transform 1 0 3992 0 1 2570
box -8 -3 16 105
use FILL  FILL_5305
timestamp 1677677812
transform 1 0 4000 0 1 2570
box -8 -3 16 105
use FILL  FILL_5307
timestamp 1677677812
transform 1 0 4008 0 1 2570
box -8 -3 16 105
use FILL  FILL_5309
timestamp 1677677812
transform 1 0 4016 0 1 2570
box -8 -3 16 105
use FILL  FILL_5311
timestamp 1677677812
transform 1 0 4024 0 1 2570
box -8 -3 16 105
use FILL  FILL_5313
timestamp 1677677812
transform 1 0 4032 0 1 2570
box -8 -3 16 105
use FILL  FILL_5315
timestamp 1677677812
transform 1 0 4040 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4068
timestamp 1677677812
transform 1 0 4068 0 1 2575
box -3 -3 3 3
use OAI22X1  OAI22X1_203
timestamp 1677677812
transform 1 0 4048 0 1 2570
box -8 -3 46 105
use FILL  FILL_5317
timestamp 1677677812
transform 1 0 4088 0 1 2570
box -8 -3 16 105
use FILL  FILL_5324
timestamp 1677677812
transform 1 0 4096 0 1 2570
box -8 -3 16 105
use FILL  FILL_5326
timestamp 1677677812
transform 1 0 4104 0 1 2570
box -8 -3 16 105
use FILL  FILL_5327
timestamp 1677677812
transform 1 0 4112 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4069
timestamp 1677677812
transform 1 0 4132 0 1 2575
box -3 -3 3 3
use INVX2  INVX2_358
timestamp 1677677812
transform -1 0 4136 0 1 2570
box -9 -3 26 105
use FILL  FILL_5328
timestamp 1677677812
transform 1 0 4136 0 1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_311
timestamp 1677677812
transform -1 0 4240 0 1 2570
box -8 -3 104 105
use FILL  FILL_5329
timestamp 1677677812
transform 1 0 4240 0 1 2570
box -8 -3 16 105
use FILL  FILL_5330
timestamp 1677677812
transform 1 0 4248 0 1 2570
box -8 -3 16 105
use FILL  FILL_5331
timestamp 1677677812
transform 1 0 4256 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_32
timestamp 1677677812
transform 1 0 4264 0 1 2570
box -8 -3 40 105
use FILL  FILL_5332
timestamp 1677677812
transform 1 0 4296 0 1 2570
box -8 -3 16 105
use FILL  FILL_5339
timestamp 1677677812
transform 1 0 4304 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_360
timestamp 1677677812
transform 1 0 4312 0 1 2570
box -9 -3 26 105
use FILL  FILL_5341
timestamp 1677677812
transform 1 0 4328 0 1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_33
timestamp 1677677812
transform -1 0 4368 0 1 2570
box -8 -3 40 105
use FILL  FILL_5342
timestamp 1677677812
transform 1 0 4368 0 1 2570
box -8 -3 16 105
use FILL  FILL_5346
timestamp 1677677812
transform 1 0 4376 0 1 2570
box -8 -3 16 105
use FILL  FILL_5348
timestamp 1677677812
transform 1 0 4384 0 1 2570
box -8 -3 16 105
use FILL  FILL_5349
timestamp 1677677812
transform 1 0 4392 0 1 2570
box -8 -3 16 105
use FILL  FILL_5350
timestamp 1677677812
transform 1 0 4400 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_206
timestamp 1677677812
transform 1 0 4408 0 1 2570
box -8 -3 46 105
use FILL  FILL_5351
timestamp 1677677812
transform 1 0 4448 0 1 2570
box -8 -3 16 105
use FILL  FILL_5352
timestamp 1677677812
transform 1 0 4456 0 1 2570
box -8 -3 16 105
use BUFX2  BUFX2_48
timestamp 1677677812
transform 1 0 4464 0 1 2570
box -5 -3 28 105
use FILL  FILL_5353
timestamp 1677677812
transform 1 0 4488 0 1 2570
box -8 -3 16 105
use FILL  FILL_5361
timestamp 1677677812
transform 1 0 4496 0 1 2570
box -8 -3 16 105
use FILL  FILL_5363
timestamp 1677677812
transform 1 0 4504 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4070
timestamp 1677677812
transform 1 0 4580 0 1 2575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_313
timestamp 1677677812
transform 1 0 4512 0 1 2570
box -8 -3 104 105
use FILL  FILL_5365
timestamp 1677677812
transform 1 0 4608 0 1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4071
timestamp 1677677812
transform 1 0 4644 0 1 2575
box -3 -3 3 3
use AOI22X1  AOI22X1_220
timestamp 1677677812
transform -1 0 4656 0 1 2570
box -8 -3 46 105
use FILL  FILL_5366
timestamp 1677677812
transform 1 0 4656 0 1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_207
timestamp 1677677812
transform 1 0 4664 0 1 2570
box -8 -3 46 105
use FILL  FILL_5367
timestamp 1677677812
transform 1 0 4704 0 1 2570
box -8 -3 16 105
use FILL  FILL_5368
timestamp 1677677812
transform 1 0 4712 0 1 2570
box -8 -3 16 105
use FILL  FILL_5369
timestamp 1677677812
transform 1 0 4720 0 1 2570
box -8 -3 16 105
use INVX2  INVX2_362
timestamp 1677677812
transform -1 0 4744 0 1 2570
box -9 -3 26 105
use FILL  FILL_5370
timestamp 1677677812
transform 1 0 4744 0 1 2570
box -8 -3 16 105
use FILL  FILL_5371
timestamp 1677677812
transform 1 0 4752 0 1 2570
box -8 -3 16 105
use FILL  FILL_5372
timestamp 1677677812
transform 1 0 4760 0 1 2570
box -8 -3 16 105
use FILL  FILL_5373
timestamp 1677677812
transform 1 0 4768 0 1 2570
box -8 -3 16 105
use FILL  FILL_5374
timestamp 1677677812
transform 1 0 4776 0 1 2570
box -8 -3 16 105
use FILL  FILL_5375
timestamp 1677677812
transform 1 0 4784 0 1 2570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_43
timestamp 1677677812
transform 1 0 4819 0 1 2570
box -10 -3 10 3
use M3_M2  M3_M2_4096
timestamp 1677677812
transform 1 0 164 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4547
timestamp 1677677812
transform 1 0 84 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4640
timestamp 1677677812
transform 1 0 108 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4641
timestamp 1677677812
transform 1 0 164 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4548
timestamp 1677677812
transform 1 0 204 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4549
timestamp 1677677812
transform 1 0 228 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4642
timestamp 1677677812
transform 1 0 212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4643
timestamp 1677677812
transform 1 0 252 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4164
timestamp 1677677812
transform 1 0 212 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4165
timestamp 1677677812
transform 1 0 252 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4201
timestamp 1677677812
transform 1 0 204 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4202
timestamp 1677677812
transform 1 0 244 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4211
timestamp 1677677812
transform 1 0 228 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4212
timestamp 1677677812
transform 1 0 292 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4543
timestamp 1677677812
transform 1 0 332 0 1 2545
box -2 -2 2 2
use M2_M1  M2_M1_4644
timestamp 1677677812
transform 1 0 332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4645
timestamp 1677677812
transform 1 0 348 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4550
timestamp 1677677812
transform 1 0 364 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4646
timestamp 1677677812
transform 1 0 372 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4551
timestamp 1677677812
transform 1 0 396 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4647
timestamp 1677677812
transform 1 0 404 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4213
timestamp 1677677812
transform 1 0 404 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4110
timestamp 1677677812
transform 1 0 564 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4552
timestamp 1677677812
transform 1 0 484 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4553
timestamp 1677677812
transform 1 0 572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4648
timestamp 1677677812
transform 1 0 508 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4649
timestamp 1677677812
transform 1 0 564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4650
timestamp 1677677812
transform 1 0 572 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4166
timestamp 1677677812
transform 1 0 508 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4214
timestamp 1677677812
transform 1 0 540 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4167
timestamp 1677677812
transform 1 0 572 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4072
timestamp 1677677812
transform 1 0 588 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4153
timestamp 1677677812
transform 1 0 588 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4111
timestamp 1677677812
transform 1 0 612 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4554
timestamp 1677677812
transform 1 0 612 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4651
timestamp 1677677812
transform 1 0 620 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4097
timestamp 1677677812
transform 1 0 676 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4112
timestamp 1677677812
transform 1 0 668 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4555
timestamp 1677677812
transform 1 0 660 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4556
timestamp 1677677812
transform 1 0 676 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4652
timestamp 1677677812
transform 1 0 668 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4168
timestamp 1677677812
transform 1 0 668 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4169
timestamp 1677677812
transform 1 0 692 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4653
timestamp 1677677812
transform 1 0 716 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4654
timestamp 1677677812
transform 1 0 756 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4098
timestamp 1677677812
transform 1 0 828 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4557
timestamp 1677677812
transform 1 0 804 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4558
timestamp 1677677812
transform 1 0 812 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4559
timestamp 1677677812
transform 1 0 828 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4655
timestamp 1677677812
transform 1 0 820 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4656
timestamp 1677677812
transform 1 0 836 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4560
timestamp 1677677812
transform 1 0 892 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4073
timestamp 1677677812
transform 1 0 924 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4561
timestamp 1677677812
transform 1 0 932 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4657
timestamp 1677677812
transform 1 0 908 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4658
timestamp 1677677812
transform 1 0 924 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4198
timestamp 1677677812
transform 1 0 924 0 1 2505
box -3 -3 3 3
use M2_M1  M2_M1_4544
timestamp 1677677812
transform 1 0 948 0 1 2545
box -2 -2 2 2
use M3_M2  M3_M2_4074
timestamp 1677677812
transform 1 0 1020 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4203
timestamp 1677677812
transform 1 0 1012 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4562
timestamp 1677677812
transform 1 0 1036 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4154
timestamp 1677677812
transform 1 0 1036 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4170
timestamp 1677677812
transform 1 0 1052 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4075
timestamp 1677677812
transform 1 0 1068 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4099
timestamp 1677677812
transform 1 0 1084 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4100
timestamp 1677677812
transform 1 0 1100 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4563
timestamp 1677677812
transform 1 0 1076 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4564
timestamp 1677677812
transform 1 0 1084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4659
timestamp 1677677812
transform 1 0 1068 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4140
timestamp 1677677812
transform 1 0 1092 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4101
timestamp 1677677812
transform 1 0 1116 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4565
timestamp 1677677812
transform 1 0 1108 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4660
timestamp 1677677812
transform 1 0 1092 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4155
timestamp 1677677812
transform 1 0 1100 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4171
timestamp 1677677812
transform 1 0 1076 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4172
timestamp 1677677812
transform 1 0 1092 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4113
timestamp 1677677812
transform 1 0 1132 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4141
timestamp 1677677812
transform 1 0 1132 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4156
timestamp 1677677812
transform 1 0 1124 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4661
timestamp 1677677812
transform 1 0 1132 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4173
timestamp 1677677812
transform 1 0 1140 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4662
timestamp 1677677812
transform 1 0 1172 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4102
timestamp 1677677812
transform 1 0 1196 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4566
timestamp 1677677812
transform 1 0 1188 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4663
timestamp 1677677812
transform 1 0 1196 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4664
timestamp 1677677812
transform 1 0 1212 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4665
timestamp 1677677812
transform 1 0 1228 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4567
timestamp 1677677812
transform 1 0 1260 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4752
timestamp 1677677812
transform 1 0 1268 0 1 2505
box -2 -2 2 2
use M3_M2  M3_M2_4114
timestamp 1677677812
transform 1 0 1284 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4666
timestamp 1677677812
transform 1 0 1284 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4174
timestamp 1677677812
transform 1 0 1284 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4215
timestamp 1677677812
transform 1 0 1292 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4076
timestamp 1677677812
transform 1 0 1316 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4115
timestamp 1677677812
transform 1 0 1308 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4568
timestamp 1677677812
transform 1 0 1316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4742
timestamp 1677677812
transform 1 0 1308 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4216
timestamp 1677677812
transform 1 0 1308 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4667
timestamp 1677677812
transform 1 0 1324 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4116
timestamp 1677677812
transform 1 0 1364 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4569
timestamp 1677677812
transform 1 0 1364 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4668
timestamp 1677677812
transform 1 0 1388 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4669
timestamp 1677677812
transform 1 0 1404 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4743
timestamp 1677677812
transform 1 0 1436 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4117
timestamp 1677677812
transform 1 0 1452 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4570
timestamp 1677677812
transform 1 0 1452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4670
timestamp 1677677812
transform 1 0 1484 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4217
timestamp 1677677812
transform 1 0 1476 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4571
timestamp 1677677812
transform 1 0 1572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4671
timestamp 1677677812
transform 1 0 1548 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4218
timestamp 1677677812
transform 1 0 1516 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4572
timestamp 1677677812
transform 1 0 1588 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4573
timestamp 1677677812
transform 1 0 1604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4672
timestamp 1677677812
transform 1 0 1604 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4118
timestamp 1677677812
transform 1 0 1620 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4574
timestamp 1677677812
transform 1 0 1628 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4673
timestamp 1677677812
transform 1 0 1676 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4077
timestamp 1677677812
transform 1 0 1692 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4078
timestamp 1677677812
transform 1 0 1724 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4079
timestamp 1677677812
transform 1 0 1764 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4119
timestamp 1677677812
transform 1 0 1716 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4575
timestamp 1677677812
transform 1 0 1764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4674
timestamp 1677677812
transform 1 0 1716 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4204
timestamp 1677677812
transform 1 0 1684 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4576
timestamp 1677677812
transform 1 0 1780 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4219
timestamp 1677677812
transform 1 0 1780 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4675
timestamp 1677677812
transform 1 0 1812 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4080
timestamp 1677677812
transform 1 0 1828 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4676
timestamp 1677677812
transform 1 0 1836 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4081
timestamp 1677677812
transform 1 0 1908 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4120
timestamp 1677677812
transform 1 0 1876 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4121
timestamp 1677677812
transform 1 0 1900 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4577
timestamp 1677677812
transform 1 0 1876 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4578
timestamp 1677677812
transform 1 0 1892 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4579
timestamp 1677677812
transform 1 0 1900 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4677
timestamp 1677677812
transform 1 0 1868 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4678
timestamp 1677677812
transform 1 0 1884 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4122
timestamp 1677677812
transform 1 0 1980 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4580
timestamp 1677677812
transform 1 0 1980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4679
timestamp 1677677812
transform 1 0 1964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4680
timestamp 1677677812
transform 1 0 1972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4681
timestamp 1677677812
transform 1 0 1988 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4175
timestamp 1677677812
transform 1 0 1964 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4682
timestamp 1677677812
transform 1 0 2012 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4176
timestamp 1677677812
transform 1 0 2012 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4123
timestamp 1677677812
transform 1 0 2076 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4683
timestamp 1677677812
transform 1 0 2068 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4581
timestamp 1677677812
transform 1 0 2100 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4082
timestamp 1677677812
transform 1 0 2132 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4124
timestamp 1677677812
transform 1 0 2132 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4582
timestamp 1677677812
transform 1 0 2132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4583
timestamp 1677677812
transform 1 0 2156 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4157
timestamp 1677677812
transform 1 0 2156 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4684
timestamp 1677677812
transform 1 0 2220 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4584
timestamp 1677677812
transform 1 0 2244 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4083
timestamp 1677677812
transform 1 0 2260 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4585
timestamp 1677677812
transform 1 0 2260 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4142
timestamp 1677677812
transform 1 0 2292 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4685
timestamp 1677677812
transform 1 0 2292 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4084
timestamp 1677677812
transform 1 0 2308 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4586
timestamp 1677677812
transform 1 0 2316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4587
timestamp 1677677812
transform 1 0 2332 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4588
timestamp 1677677812
transform 1 0 2340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4686
timestamp 1677677812
transform 1 0 2308 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4687
timestamp 1677677812
transform 1 0 2324 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4205
timestamp 1677677812
transform 1 0 2316 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4143
timestamp 1677677812
transform 1 0 2364 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4688
timestamp 1677677812
transform 1 0 2356 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4206
timestamp 1677677812
transform 1 0 2348 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4689
timestamp 1677677812
transform 1 0 2388 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4085
timestamp 1677677812
transform 1 0 2436 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4589
timestamp 1677677812
transform 1 0 2436 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4690
timestamp 1677677812
transform 1 0 2420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4691
timestamp 1677677812
transform 1 0 2428 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4692
timestamp 1677677812
transform 1 0 2444 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4220
timestamp 1677677812
transform 1 0 2428 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4590
timestamp 1677677812
transform 1 0 2460 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4144
timestamp 1677677812
transform 1 0 2492 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4693
timestamp 1677677812
transform 1 0 2532 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4591
timestamp 1677677812
transform 1 0 2548 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4592
timestamp 1677677812
transform 1 0 2564 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4593
timestamp 1677677812
transform 1 0 2572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4694
timestamp 1677677812
transform 1 0 2556 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4207
timestamp 1677677812
transform 1 0 2564 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4695
timestamp 1677677812
transform 1 0 2588 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4696
timestamp 1677677812
transform 1 0 2620 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4697
timestamp 1677677812
transform 1 0 2660 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4177
timestamp 1677677812
transform 1 0 2660 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4594
timestamp 1677677812
transform 1 0 2676 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4595
timestamp 1677677812
transform 1 0 2764 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4698
timestamp 1677677812
transform 1 0 2700 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4699
timestamp 1677677812
transform 1 0 2756 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4178
timestamp 1677677812
transform 1 0 2700 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4208
timestamp 1677677812
transform 1 0 2756 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4596
timestamp 1677677812
transform 1 0 2796 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4700
timestamp 1677677812
transform 1 0 2788 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4158
timestamp 1677677812
transform 1 0 2820 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4701
timestamp 1677677812
transform 1 0 2828 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4086
timestamp 1677677812
transform 1 0 2868 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4597
timestamp 1677677812
transform 1 0 2860 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4545
timestamp 1677677812
transform 1 0 2868 0 1 2545
box -2 -2 2 2
use M3_M2  M3_M2_4087
timestamp 1677677812
transform 1 0 2892 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4125
timestamp 1677677812
transform 1 0 2884 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4744
timestamp 1677677812
transform 1 0 2892 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4598
timestamp 1677677812
transform 1 0 2908 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4159
timestamp 1677677812
transform 1 0 2908 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4088
timestamp 1677677812
transform 1 0 2924 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4126
timestamp 1677677812
transform 1 0 2924 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4599
timestamp 1677677812
transform 1 0 2924 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4702
timestamp 1677677812
transform 1 0 2916 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4703
timestamp 1677677812
transform 1 0 2972 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4745
timestamp 1677677812
transform 1 0 2956 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4179
timestamp 1677677812
transform 1 0 2972 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4600
timestamp 1677677812
transform 1 0 2996 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4704
timestamp 1677677812
transform 1 0 2996 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4180
timestamp 1677677812
transform 1 0 3004 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4127
timestamp 1677677812
transform 1 0 3020 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4601
timestamp 1677677812
transform 1 0 3020 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4221
timestamp 1677677812
transform 1 0 3028 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4128
timestamp 1677677812
transform 1 0 3124 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4602
timestamp 1677677812
transform 1 0 3060 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4129
timestamp 1677677812
transform 1 0 3156 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4705
timestamp 1677677812
transform 1 0 3044 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4706
timestamp 1677677812
transform 1 0 3084 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4707
timestamp 1677677812
transform 1 0 3140 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4708
timestamp 1677677812
transform 1 0 3148 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4181
timestamp 1677677812
transform 1 0 3044 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4182
timestamp 1677677812
transform 1 0 3148 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4603
timestamp 1677677812
transform 1 0 3180 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4604
timestamp 1677677812
transform 1 0 3196 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4183
timestamp 1677677812
transform 1 0 3196 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4089
timestamp 1677677812
transform 1 0 3220 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4709
timestamp 1677677812
transform 1 0 3260 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4130
timestamp 1677677812
transform 1 0 3316 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4605
timestamp 1677677812
transform 1 0 3316 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4746
timestamp 1677677812
transform 1 0 3308 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4131
timestamp 1677677812
transform 1 0 3340 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4184
timestamp 1677677812
transform 1 0 3340 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4747
timestamp 1677677812
transform 1 0 3356 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4753
timestamp 1677677812
transform 1 0 3340 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4606
timestamp 1677677812
transform 1 0 3396 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4160
timestamp 1677677812
transform 1 0 3388 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4748
timestamp 1677677812
transform 1 0 3404 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4754
timestamp 1677677812
transform 1 0 3388 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4710
timestamp 1677677812
transform 1 0 3420 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4222
timestamp 1677677812
transform 1 0 3420 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4711
timestamp 1677677812
transform 1 0 3436 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4223
timestamp 1677677812
transform 1 0 3436 0 1 2485
box -3 -3 3 3
use M2_M1  M2_M1_4607
timestamp 1677677812
transform 1 0 3452 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4608
timestamp 1677677812
transform 1 0 3468 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4749
timestamp 1677677812
transform 1 0 3460 0 1 2515
box -2 -2 2 2
use M3_M2  M3_M2_4224
timestamp 1677677812
transform 1 0 3460 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4103
timestamp 1677677812
transform 1 0 3492 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4712
timestamp 1677677812
transform 1 0 3500 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4609
timestamp 1677677812
transform 1 0 3516 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4750
timestamp 1677677812
transform 1 0 3508 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4755
timestamp 1677677812
transform 1 0 3492 0 1 2505
box -2 -2 2 2
use M2_M1  M2_M1_4610
timestamp 1677677812
transform 1 0 3556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4611
timestamp 1677677812
transform 1 0 3572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4713
timestamp 1677677812
transform 1 0 3548 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4714
timestamp 1677677812
transform 1 0 3564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4751
timestamp 1677677812
transform 1 0 3580 0 1 2515
box -2 -2 2 2
use M2_M1  M2_M1_4715
timestamp 1677677812
transform 1 0 3588 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4612
timestamp 1677677812
transform 1 0 3604 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4613
timestamp 1677677812
transform 1 0 3620 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4716
timestamp 1677677812
transform 1 0 3676 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4185
timestamp 1677677812
transform 1 0 3676 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4145
timestamp 1677677812
transform 1 0 3692 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4717
timestamp 1677677812
transform 1 0 3692 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4090
timestamp 1677677812
transform 1 0 3724 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4091
timestamp 1677677812
transform 1 0 3740 0 1 2565
box -3 -3 3 3
use M2_M1  M2_M1_4614
timestamp 1677677812
transform 1 0 3716 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4146
timestamp 1677677812
transform 1 0 3724 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4104
timestamp 1677677812
transform 1 0 3756 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4105
timestamp 1677677812
transform 1 0 3788 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4106
timestamp 1677677812
transform 1 0 3836 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4615
timestamp 1677677812
transform 1 0 3740 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4616
timestamp 1677677812
transform 1 0 3756 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4718
timestamp 1677677812
transform 1 0 3724 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4719
timestamp 1677677812
transform 1 0 3788 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4186
timestamp 1677677812
transform 1 0 3780 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4187
timestamp 1677677812
transform 1 0 3820 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4107
timestamp 1677677812
transform 1 0 3876 0 1 2555
box -3 -3 3 3
use M2_M1  M2_M1_4617
timestamp 1677677812
transform 1 0 3892 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4147
timestamp 1677677812
transform 1 0 3900 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4720
timestamp 1677677812
transform 1 0 3876 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4721
timestamp 1677677812
transform 1 0 3884 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4722
timestamp 1677677812
transform 1 0 3900 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4723
timestamp 1677677812
transform 1 0 3916 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4188
timestamp 1677677812
transform 1 0 3884 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4189
timestamp 1677677812
transform 1 0 3908 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4209
timestamp 1677677812
transform 1 0 3876 0 1 2495
box -3 -3 3 3
use M3_M2  M3_M2_4210
timestamp 1677677812
transform 1 0 3916 0 1 2495
box -3 -3 3 3
use M2_M1  M2_M1_4724
timestamp 1677677812
transform 1 0 3964 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4618
timestamp 1677677812
transform 1 0 3980 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4619
timestamp 1677677812
transform 1 0 4044 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4620
timestamp 1677677812
transform 1 0 4084 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4621
timestamp 1677677812
transform 1 0 4116 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4148
timestamp 1677677812
transform 1 0 4124 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4622
timestamp 1677677812
transform 1 0 4132 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4623
timestamp 1677677812
transform 1 0 4148 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4161
timestamp 1677677812
transform 1 0 4116 0 1 2525
box -3 -3 3 3
use M2_M1  M2_M1_4725
timestamp 1677677812
transform 1 0 4124 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4726
timestamp 1677677812
transform 1 0 4140 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4190
timestamp 1677677812
transform 1 0 4140 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4092
timestamp 1677677812
transform 1 0 4196 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4093
timestamp 1677677812
transform 1 0 4228 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4132
timestamp 1677677812
transform 1 0 4244 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4624
timestamp 1677677812
transform 1 0 4196 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4625
timestamp 1677677812
transform 1 0 4284 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4727
timestamp 1677677812
transform 1 0 4244 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4728
timestamp 1677677812
transform 1 0 4276 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4729
timestamp 1677677812
transform 1 0 4284 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4162
timestamp 1677677812
transform 1 0 4292 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4191
timestamp 1677677812
transform 1 0 4244 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4192
timestamp 1677677812
transform 1 0 4284 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4626
timestamp 1677677812
transform 1 0 4308 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4163
timestamp 1677677812
transform 1 0 4308 0 1 2525
box -3 -3 3 3
use M3_M2  M3_M2_4108
timestamp 1677677812
transform 1 0 4332 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4109
timestamp 1677677812
transform 1 0 4364 0 1 2555
box -3 -3 3 3
use M3_M2  M3_M2_4133
timestamp 1677677812
transform 1 0 4340 0 1 2545
box -3 -3 3 3
use M3_M2  M3_M2_4134
timestamp 1677677812
transform 1 0 4356 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4627
timestamp 1677677812
transform 1 0 4340 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4628
timestamp 1677677812
transform 1 0 4356 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4629
timestamp 1677677812
transform 1 0 4364 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4730
timestamp 1677677812
transform 1 0 4332 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4731
timestamp 1677677812
transform 1 0 4348 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4193
timestamp 1677677812
transform 1 0 4348 0 1 2515
box -3 -3 3 3
use M2_M1  M2_M1_4732
timestamp 1677677812
transform 1 0 4380 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4149
timestamp 1677677812
transform 1 0 4412 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4733
timestamp 1677677812
transform 1 0 4404 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4734
timestamp 1677677812
transform 1 0 4420 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4546
timestamp 1677677812
transform 1 0 4436 0 1 2545
box -2 -2 2 2
use M3_M2  M3_M2_4150
timestamp 1677677812
transform 1 0 4444 0 1 2535
box -3 -3 3 3
use M3_M2  M3_M2_4135
timestamp 1677677812
transform 1 0 4468 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4630
timestamp 1677677812
transform 1 0 4460 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4631
timestamp 1677677812
transform 1 0 4468 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4136
timestamp 1677677812
transform 1 0 4556 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4632
timestamp 1677677812
transform 1 0 4556 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4633
timestamp 1677677812
transform 1 0 4572 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4735
timestamp 1677677812
transform 1 0 4548 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4736
timestamp 1677677812
transform 1 0 4564 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4737
timestamp 1677677812
transform 1 0 4580 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4634
timestamp 1677677812
transform 1 0 4604 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4194
timestamp 1677677812
transform 1 0 4604 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4094
timestamp 1677677812
transform 1 0 4644 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4137
timestamp 1677677812
transform 1 0 4652 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4635
timestamp 1677677812
transform 1 0 4628 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4151
timestamp 1677677812
transform 1 0 4636 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4636
timestamp 1677677812
transform 1 0 4644 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4138
timestamp 1677677812
transform 1 0 4684 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4637
timestamp 1677677812
transform 1 0 4668 0 1 2535
box -2 -2 2 2
use M3_M2  M3_M2_4152
timestamp 1677677812
transform 1 0 4676 0 1 2535
box -3 -3 3 3
use M2_M1  M2_M1_4638
timestamp 1677677812
transform 1 0 4684 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4738
timestamp 1677677812
transform 1 0 4660 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4739
timestamp 1677677812
transform 1 0 4676 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4195
timestamp 1677677812
transform 1 0 4636 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4196
timestamp 1677677812
transform 1 0 4652 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4199
timestamp 1677677812
transform 1 0 4660 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4095
timestamp 1677677812
transform 1 0 4740 0 1 2565
box -3 -3 3 3
use M3_M2  M3_M2_4139
timestamp 1677677812
transform 1 0 4732 0 1 2545
box -3 -3 3 3
use M2_M1  M2_M1_4639
timestamp 1677677812
transform 1 0 4708 0 1 2535
box -2 -2 2 2
use M2_M1  M2_M1_4740
timestamp 1677677812
transform 1 0 4732 0 1 2525
box -2 -2 2 2
use M2_M1  M2_M1_4741
timestamp 1677677812
transform 1 0 4788 0 1 2525
box -2 -2 2 2
use M3_M2  M3_M2_4197
timestamp 1677677812
transform 1 0 4796 0 1 2515
box -3 -3 3 3
use M3_M2  M3_M2_4200
timestamp 1677677812
transform 1 0 4732 0 1 2505
box -3 -3 3 3
use M3_M2  M3_M2_4225
timestamp 1677677812
transform 1 0 4692 0 1 2485
box -3 -3 3 3
use M3_M2  M3_M2_4226
timestamp 1677677812
transform 1 0 4724 0 1 2485
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_44
timestamp 1677677812
transform 1 0 24 0 1 2470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_294
timestamp 1677677812
transform 1 0 72 0 -1 2570
box -8 -3 104 105
use FILL  FILL_4850
timestamp 1677677812
transform 1 0 168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4851
timestamp 1677677812
transform 1 0 176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4852
timestamp 1677677812
transform 1 0 184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4853
timestamp 1677677812
transform 1 0 192 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_331
timestamp 1677677812
transform 1 0 200 0 -1 2570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_295
timestamp 1677677812
transform 1 0 216 0 -1 2570
box -8 -3 104 105
use FILL  FILL_4854
timestamp 1677677812
transform 1 0 312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4855
timestamp 1677677812
transform 1 0 320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4856
timestamp 1677677812
transform 1 0 328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4857
timestamp 1677677812
transform 1 0 336 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4863
timestamp 1677677812
transform 1 0 344 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_201
timestamp 1677677812
transform -1 0 392 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4864
timestamp 1677677812
transform 1 0 392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4866
timestamp 1677677812
transform 1 0 400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4868
timestamp 1677677812
transform 1 0 408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4871
timestamp 1677677812
transform 1 0 416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4872
timestamp 1677677812
transform 1 0 424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4873
timestamp 1677677812
transform 1 0 432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4874
timestamp 1677677812
transform 1 0 440 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4876
timestamp 1677677812
transform 1 0 448 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4878
timestamp 1677677812
transform 1 0 456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4880
timestamp 1677677812
transform 1 0 464 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_296
timestamp 1677677812
transform 1 0 472 0 -1 2570
box -8 -3 104 105
use FILL  FILL_4889
timestamp 1677677812
transform 1 0 568 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4890
timestamp 1677677812
transform 1 0 576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4891
timestamp 1677677812
transform 1 0 584 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_334
timestamp 1677677812
transform 1 0 592 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4892
timestamp 1677677812
transform 1 0 608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4894
timestamp 1677677812
transform 1 0 616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4896
timestamp 1677677812
transform 1 0 624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4898
timestamp 1677677812
transform 1 0 632 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4227
timestamp 1677677812
transform 1 0 668 0 1 2475
box -3 -3 3 3
use OAI22X1  OAI22X1_195
timestamp 1677677812
transform 1 0 640 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4905
timestamp 1677677812
transform 1 0 680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4907
timestamp 1677677812
transform 1 0 688 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4909
timestamp 1677677812
transform 1 0 696 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4911
timestamp 1677677812
transform 1 0 704 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4913
timestamp 1677677812
transform 1 0 712 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4915
timestamp 1677677812
transform 1 0 720 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_335
timestamp 1677677812
transform -1 0 744 0 -1 2570
box -9 -3 26 105
use FILL  FILL_4916
timestamp 1677677812
transform 1 0 744 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4918
timestamp 1677677812
transform 1 0 752 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4920
timestamp 1677677812
transform 1 0 760 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4922
timestamp 1677677812
transform 1 0 768 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4924
timestamp 1677677812
transform 1 0 776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4926
timestamp 1677677812
transform 1 0 784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4932
timestamp 1677677812
transform 1 0 792 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_204
timestamp 1677677812
transform -1 0 840 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4933
timestamp 1677677812
transform 1 0 840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4935
timestamp 1677677812
transform 1 0 848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4936
timestamp 1677677812
transform 1 0 856 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4937
timestamp 1677677812
transform 1 0 864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4938
timestamp 1677677812
transform 1 0 872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4939
timestamp 1677677812
transform 1 0 880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4940
timestamp 1677677812
transform 1 0 888 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4945
timestamp 1677677812
transform 1 0 896 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_207
timestamp 1677677812
transform -1 0 944 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4946
timestamp 1677677812
transform 1 0 944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4947
timestamp 1677677812
transform 1 0 952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4948
timestamp 1677677812
transform 1 0 960 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4950
timestamp 1677677812
transform 1 0 968 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4952
timestamp 1677677812
transform 1 0 976 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4954
timestamp 1677677812
transform 1 0 984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4956
timestamp 1677677812
transform 1 0 992 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_50
timestamp 1677677812
transform 1 0 1000 0 -1 2570
box -8 -3 32 105
use FILL  FILL_4960
timestamp 1677677812
transform 1 0 1024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4961
timestamp 1677677812
transform 1 0 1032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4962
timestamp 1677677812
transform 1 0 1040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4963
timestamp 1677677812
transform 1 0 1048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4964
timestamp 1677677812
transform 1 0 1056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4965
timestamp 1677677812
transform 1 0 1064 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_208
timestamp 1677677812
transform 1 0 1072 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4966
timestamp 1677677812
transform 1 0 1112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4967
timestamp 1677677812
transform 1 0 1120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4968
timestamp 1677677812
transform 1 0 1128 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4970
timestamp 1677677812
transform 1 0 1136 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4972
timestamp 1677677812
transform 1 0 1144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4979
timestamp 1677677812
transform 1 0 1152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4980
timestamp 1677677812
transform 1 0 1160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4981
timestamp 1677677812
transform 1 0 1168 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_209
timestamp 1677677812
transform 1 0 1176 0 -1 2570
box -8 -3 46 105
use FILL  FILL_4982
timestamp 1677677812
transform 1 0 1216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4983
timestamp 1677677812
transform 1 0 1224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4984
timestamp 1677677812
transform 1 0 1232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4985
timestamp 1677677812
transform 1 0 1240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4986
timestamp 1677677812
transform 1 0 1248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4988
timestamp 1677677812
transform 1 0 1256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4990
timestamp 1677677812
transform 1 0 1264 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_102
timestamp 1677677812
transform 1 0 1272 0 -1 2570
box -8 -3 34 105
use FILL  FILL_4995
timestamp 1677677812
transform 1 0 1304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4996
timestamp 1677677812
transform 1 0 1312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4997
timestamp 1677677812
transform 1 0 1320 0 -1 2570
box -8 -3 16 105
use FILL  FILL_4998
timestamp 1677677812
transform 1 0 1328 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5000
timestamp 1677677812
transform 1 0 1336 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_338
timestamp 1677677812
transform 1 0 1344 0 -1 2570
box -9 -3 26 105
use NAND2X1  NAND2X1_2
timestamp 1677677812
transform 1 0 1360 0 -1 2570
box -8 -3 32 105
use FILL  FILL_5006
timestamp 1677677812
transform 1 0 1384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5007
timestamp 1677677812
transform 1 0 1392 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5008
timestamp 1677677812
transform 1 0 1400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5009
timestamp 1677677812
transform 1 0 1408 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5011
timestamp 1677677812
transform 1 0 1416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5015
timestamp 1677677812
transform 1 0 1424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5016
timestamp 1677677812
transform 1 0 1432 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_340
timestamp 1677677812
transform -1 0 1456 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5017
timestamp 1677677812
transform 1 0 1456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5019
timestamp 1677677812
transform 1 0 1464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5023
timestamp 1677677812
transform 1 0 1472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5024
timestamp 1677677812
transform 1 0 1480 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_299
timestamp 1677677812
transform -1 0 1584 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5025
timestamp 1677677812
transform 1 0 1584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5029
timestamp 1677677812
transform 1 0 1592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5030
timestamp 1677677812
transform 1 0 1600 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_342
timestamp 1677677812
transform 1 0 1608 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5031
timestamp 1677677812
transform 1 0 1624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5032
timestamp 1677677812
transform 1 0 1632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5033
timestamp 1677677812
transform 1 0 1640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5034
timestamp 1677677812
transform 1 0 1648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5035
timestamp 1677677812
transform 1 0 1656 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5036
timestamp 1677677812
transform 1 0 1664 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5048
timestamp 1677677812
transform 1 0 1672 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_300
timestamp 1677677812
transform -1 0 1776 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5049
timestamp 1677677812
transform 1 0 1776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5051
timestamp 1677677812
transform 1 0 1784 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4228
timestamp 1677677812
transform 1 0 1820 0 1 2475
box -3 -3 3 3
use BUFX2  BUFX2_38
timestamp 1677677812
transform -1 0 1816 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5052
timestamp 1677677812
transform 1 0 1816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5053
timestamp 1677677812
transform 1 0 1824 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5054
timestamp 1677677812
transform 1 0 1832 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5056
timestamp 1677677812
transform 1 0 1840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5058
timestamp 1677677812
transform 1 0 1848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5060
timestamp 1677677812
transform 1 0 1856 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_210
timestamp 1677677812
transform 1 0 1864 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5068
timestamp 1677677812
transform 1 0 1904 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5069
timestamp 1677677812
transform 1 0 1912 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5070
timestamp 1677677812
transform 1 0 1920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5071
timestamp 1677677812
transform 1 0 1928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5072
timestamp 1677677812
transform 1 0 1936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5073
timestamp 1677677812
transform 1 0 1944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5074
timestamp 1677677812
transform 1 0 1952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5075
timestamp 1677677812
transform 1 0 1960 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_211
timestamp 1677677812
transform 1 0 1968 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5076
timestamp 1677677812
transform 1 0 2008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5077
timestamp 1677677812
transform 1 0 2016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5078
timestamp 1677677812
transform 1 0 2024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5079
timestamp 1677677812
transform 1 0 2032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5080
timestamp 1677677812
transform 1 0 2040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5081
timestamp 1677677812
transform 1 0 2048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5082
timestamp 1677677812
transform 1 0 2056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5083
timestamp 1677677812
transform 1 0 2064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5084
timestamp 1677677812
transform 1 0 2072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5085
timestamp 1677677812
transform 1 0 2080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5086
timestamp 1677677812
transform 1 0 2088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5087
timestamp 1677677812
transform 1 0 2096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5088
timestamp 1677677812
transform 1 0 2104 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5089
timestamp 1677677812
transform 1 0 2112 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5090
timestamp 1677677812
transform 1 0 2120 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5091
timestamp 1677677812
transform 1 0 2128 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_346
timestamp 1677677812
transform 1 0 2136 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5092
timestamp 1677677812
transform 1 0 2152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5093
timestamp 1677677812
transform 1 0 2160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5094
timestamp 1677677812
transform 1 0 2168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5095
timestamp 1677677812
transform 1 0 2176 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5096
timestamp 1677677812
transform 1 0 2184 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_39
timestamp 1677677812
transform -1 0 2216 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5097
timestamp 1677677812
transform 1 0 2216 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5098
timestamp 1677677812
transform 1 0 2224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5099
timestamp 1677677812
transform 1 0 2232 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_347
timestamp 1677677812
transform 1 0 2240 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5100
timestamp 1677677812
transform 1 0 2256 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5101
timestamp 1677677812
transform 1 0 2264 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5102
timestamp 1677677812
transform 1 0 2272 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5103
timestamp 1677677812
transform 1 0 2280 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5104
timestamp 1677677812
transform 1 0 2288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5105
timestamp 1677677812
transform 1 0 2296 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_212
timestamp 1677677812
transform 1 0 2304 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5106
timestamp 1677677812
transform 1 0 2344 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5108
timestamp 1677677812
transform 1 0 2352 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5110
timestamp 1677677812
transform 1 0 2360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5112
timestamp 1677677812
transform 1 0 2368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5114
timestamp 1677677812
transform 1 0 2376 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5116
timestamp 1677677812
transform 1 0 2384 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5118
timestamp 1677677812
transform 1 0 2392 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4229
timestamp 1677677812
transform 1 0 2412 0 1 2475
box -3 -3 3 3
use FILL  FILL_5122
timestamp 1677677812
transform 1 0 2400 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5123
timestamp 1677677812
transform 1 0 2408 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4230
timestamp 1677677812
transform 1 0 2428 0 1 2475
box -3 -3 3 3
use OAI22X1  OAI22X1_198
timestamp 1677677812
transform 1 0 2416 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5124
timestamp 1677677812
transform 1 0 2456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5126
timestamp 1677677812
transform 1 0 2464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5128
timestamp 1677677812
transform 1 0 2472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5130
timestamp 1677677812
transform 1 0 2480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5133
timestamp 1677677812
transform 1 0 2488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5134
timestamp 1677677812
transform 1 0 2496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5135
timestamp 1677677812
transform 1 0 2504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5136
timestamp 1677677812
transform 1 0 2512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5137
timestamp 1677677812
transform 1 0 2520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5138
timestamp 1677677812
transform 1 0 2528 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_213
timestamp 1677677812
transform 1 0 2536 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5139
timestamp 1677677812
transform 1 0 2576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5140
timestamp 1677677812
transform 1 0 2584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5141
timestamp 1677677812
transform 1 0 2592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5143
timestamp 1677677812
transform 1 0 2600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5146
timestamp 1677677812
transform 1 0 2608 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_349
timestamp 1677677812
transform 1 0 2616 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5147
timestamp 1677677812
transform 1 0 2632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5149
timestamp 1677677812
transform 1 0 2640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5151
timestamp 1677677812
transform 1 0 2648 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5153
timestamp 1677677812
transform 1 0 2656 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_306
timestamp 1677677812
transform 1 0 2664 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_350
timestamp 1677677812
transform 1 0 2760 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5161
timestamp 1677677812
transform 1 0 2776 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5163
timestamp 1677677812
transform 1 0 2784 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5165
timestamp 1677677812
transform 1 0 2792 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5167
timestamp 1677677812
transform 1 0 2800 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5169
timestamp 1677677812
transform 1 0 2808 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5171
timestamp 1677677812
transform 1 0 2816 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5174
timestamp 1677677812
transform 1 0 2824 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_105
timestamp 1677677812
transform 1 0 2832 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5175
timestamp 1677677812
transform 1 0 2864 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5177
timestamp 1677677812
transform 1 0 2872 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5179
timestamp 1677677812
transform 1 0 2880 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5181
timestamp 1677677812
transform 1 0 2888 0 -1 2570
box -8 -3 16 105
use NOR2X1  NOR2X1_53
timestamp 1677677812
transform 1 0 2896 0 -1 2570
box -8 -3 32 105
use FILL  FILL_5184
timestamp 1677677812
transform 1 0 2920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5186
timestamp 1677677812
transform 1 0 2928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5188
timestamp 1677677812
transform 1 0 2936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5193
timestamp 1677677812
transform 1 0 2944 0 -1 2570
box -8 -3 16 105
use OAI21X1  OAI21X1_107
timestamp 1677677812
transform -1 0 2984 0 -1 2570
box -8 -3 34 105
use FILL  FILL_5194
timestamp 1677677812
transform 1 0 2984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5195
timestamp 1677677812
transform 1 0 2992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5196
timestamp 1677677812
transform 1 0 3000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5197
timestamp 1677677812
transform 1 0 3008 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_40
timestamp 1677677812
transform -1 0 3040 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5198
timestamp 1677677812
transform 1 0 3040 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_308
timestamp 1677677812
transform 1 0 3048 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5205
timestamp 1677677812
transform 1 0 3144 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5206
timestamp 1677677812
transform 1 0 3152 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_41
timestamp 1677677812
transform 1 0 3160 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5207
timestamp 1677677812
transform 1 0 3184 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5213
timestamp 1677677812
transform 1 0 3192 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_43
timestamp 1677677812
transform -1 0 3224 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5214
timestamp 1677677812
transform 1 0 3224 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5215
timestamp 1677677812
transform 1 0 3232 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5216
timestamp 1677677812
transform 1 0 3240 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5217
timestamp 1677677812
transform 1 0 3248 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5218
timestamp 1677677812
transform 1 0 3256 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_44
timestamp 1677677812
transform 1 0 3264 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5219
timestamp 1677677812
transform 1 0 3288 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5220
timestamp 1677677812
transform 1 0 3296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5221
timestamp 1677677812
transform 1 0 3304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5222
timestamp 1677677812
transform 1 0 3312 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5223
timestamp 1677677812
transform 1 0 3320 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_28
timestamp 1677677812
transform -1 0 3360 0 -1 2570
box -8 -3 40 105
use FILL  FILL_5224
timestamp 1677677812
transform 1 0 3360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5227
timestamp 1677677812
transform 1 0 3368 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_29
timestamp 1677677812
transform -1 0 3408 0 -1 2570
box -8 -3 40 105
use FILL  FILL_5228
timestamp 1677677812
transform 1 0 3408 0 -1 2570
box -8 -3 16 105
use M3_M2  M3_M2_4231
timestamp 1677677812
transform 1 0 3428 0 1 2475
box -3 -3 3 3
use FILL  FILL_5229
timestamp 1677677812
transform 1 0 3416 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5231
timestamp 1677677812
transform 1 0 3424 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_45
timestamp 1677677812
transform 1 0 3432 0 -1 2570
box -5 -3 28 105
use FILL  FILL_5236
timestamp 1677677812
transform 1 0 3456 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5240
timestamp 1677677812
transform 1 0 3464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5241
timestamp 1677677812
transform 1 0 3472 0 -1 2570
box -8 -3 16 105
use NAND3X1  NAND3X1_31
timestamp 1677677812
transform -1 0 3512 0 -1 2570
box -8 -3 40 105
use FILL  FILL_5242
timestamp 1677677812
transform 1 0 3512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5246
timestamp 1677677812
transform 1 0 3520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5247
timestamp 1677677812
transform 1 0 3528 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_201
timestamp 1677677812
transform 1 0 3536 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5248
timestamp 1677677812
transform 1 0 3576 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5250
timestamp 1677677812
transform 1 0 3584 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5252
timestamp 1677677812
transform 1 0 3592 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_353
timestamp 1677677812
transform 1 0 3600 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5256
timestamp 1677677812
transform 1 0 3616 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5258
timestamp 1677677812
transform 1 0 3624 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5260
timestamp 1677677812
transform 1 0 3632 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5262
timestamp 1677677812
transform 1 0 3640 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5265
timestamp 1677677812
transform 1 0 3648 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_355
timestamp 1677677812
transform 1 0 3656 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5266
timestamp 1677677812
transform 1 0 3672 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5268
timestamp 1677677812
transform 1 0 3680 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5270
timestamp 1677677812
transform 1 0 3688 0 -1 2570
box -8 -3 16 105
use BUFX2  BUFX2_46
timestamp 1677677812
transform 1 0 3696 0 -1 2570
box -5 -3 28 105
use BUFX2  BUFX2_47
timestamp 1677677812
transform 1 0 3720 0 -1 2570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_310
timestamp 1677677812
transform 1 0 3744 0 -1 2570
box -8 -3 104 105
use FILL  FILL_5290
timestamp 1677677812
transform 1 0 3840 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5291
timestamp 1677677812
transform 1 0 3848 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5292
timestamp 1677677812
transform 1 0 3856 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_356
timestamp 1677677812
transform 1 0 3864 0 -1 2570
box -9 -3 26 105
use M3_M2  M3_M2_4232
timestamp 1677677812
transform 1 0 3900 0 1 2475
box -3 -3 3 3
use AOI22X1  AOI22X1_217
timestamp 1677677812
transform 1 0 3880 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5293
timestamp 1677677812
transform 1 0 3920 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5295
timestamp 1677677812
transform 1 0 3928 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5297
timestamp 1677677812
transform 1 0 3936 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5299
timestamp 1677677812
transform 1 0 3944 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5301
timestamp 1677677812
transform 1 0 3952 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5302
timestamp 1677677812
transform 1 0 3960 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_357
timestamp 1677677812
transform -1 0 3984 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5303
timestamp 1677677812
transform 1 0 3984 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5304
timestamp 1677677812
transform 1 0 3992 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5306
timestamp 1677677812
transform 1 0 4000 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5308
timestamp 1677677812
transform 1 0 4008 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5310
timestamp 1677677812
transform 1 0 4016 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5312
timestamp 1677677812
transform 1 0 4024 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5314
timestamp 1677677812
transform 1 0 4032 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5316
timestamp 1677677812
transform 1 0 4040 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5318
timestamp 1677677812
transform 1 0 4048 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5319
timestamp 1677677812
transform 1 0 4056 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5320
timestamp 1677677812
transform 1 0 4064 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5321
timestamp 1677677812
transform 1 0 4072 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5322
timestamp 1677677812
transform 1 0 4080 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5323
timestamp 1677677812
transform 1 0 4088 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5325
timestamp 1677677812
transform 1 0 4096 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5333
timestamp 1677677812
transform 1 0 4104 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_204
timestamp 1677677812
transform -1 0 4152 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5334
timestamp 1677677812
transform 1 0 4152 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5335
timestamp 1677677812
transform 1 0 4160 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5336
timestamp 1677677812
transform 1 0 4168 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5337
timestamp 1677677812
transform 1 0 4176 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_312
timestamp 1677677812
transform 1 0 4184 0 -1 2570
box -8 -3 104 105
use INVX2  INVX2_359
timestamp 1677677812
transform 1 0 4280 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5338
timestamp 1677677812
transform 1 0 4296 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5340
timestamp 1677677812
transform 1 0 4304 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5343
timestamp 1677677812
transform 1 0 4312 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_205
timestamp 1677677812
transform -1 0 4360 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5344
timestamp 1677677812
transform 1 0 4360 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5345
timestamp 1677677812
transform 1 0 4368 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5347
timestamp 1677677812
transform 1 0 4376 0 -1 2570
box -8 -3 16 105
use AOI22X1  AOI22X1_219
timestamp 1677677812
transform 1 0 4384 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5354
timestamp 1677677812
transform 1 0 4424 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5355
timestamp 1677677812
transform 1 0 4432 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5356
timestamp 1677677812
transform 1 0 4440 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_361
timestamp 1677677812
transform -1 0 4464 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5357
timestamp 1677677812
transform 1 0 4464 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5358
timestamp 1677677812
transform 1 0 4472 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5359
timestamp 1677677812
transform 1 0 4480 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5360
timestamp 1677677812
transform 1 0 4488 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5362
timestamp 1677677812
transform 1 0 4496 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5364
timestamp 1677677812
transform 1 0 4504 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5376
timestamp 1677677812
transform 1 0 4512 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5377
timestamp 1677677812
transform 1 0 4520 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5378
timestamp 1677677812
transform 1 0 4528 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5379
timestamp 1677677812
transform 1 0 4536 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5380
timestamp 1677677812
transform 1 0 4544 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_208
timestamp 1677677812
transform 1 0 4552 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5381
timestamp 1677677812
transform 1 0 4592 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5382
timestamp 1677677812
transform 1 0 4600 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5383
timestamp 1677677812
transform 1 0 4608 0 -1 2570
box -8 -3 16 105
use FILL  FILL_5384
timestamp 1677677812
transform 1 0 4616 0 -1 2570
box -8 -3 16 105
use INVX2  INVX2_363
timestamp 1677677812
transform 1 0 4624 0 -1 2570
box -9 -3 26 105
use FILL  FILL_5385
timestamp 1677677812
transform 1 0 4640 0 -1 2570
box -8 -3 16 105
use OAI22X1  OAI22X1_209
timestamp 1677677812
transform 1 0 4648 0 -1 2570
box -8 -3 46 105
use FILL  FILL_5386
timestamp 1677677812
transform 1 0 4688 0 -1 2570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_314
timestamp 1677677812
transform 1 0 4696 0 -1 2570
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_45
timestamp 1677677812
transform 1 0 4843 0 1 2470
box -10 -3 10 3
use M2_M1  M2_M1_4769
timestamp 1677677812
transform 1 0 124 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4291
timestamp 1677677812
transform 1 0 140 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4860
timestamp 1677677812
transform 1 0 140 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4292
timestamp 1677677812
transform 1 0 180 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4770
timestamp 1677677812
transform 1 0 164 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4771
timestamp 1677677812
transform 1 0 180 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4861
timestamp 1677677812
transform 1 0 164 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4352
timestamp 1677677812
transform 1 0 180 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4862
timestamp 1677677812
transform 1 0 188 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4372
timestamp 1677677812
transform 1 0 164 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4863
timestamp 1677677812
transform 1 0 212 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4262
timestamp 1677677812
transform 1 0 228 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4772
timestamp 1677677812
transform 1 0 228 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4773
timestamp 1677677812
transform 1 0 244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4774
timestamp 1677677812
transform 1 0 260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4864
timestamp 1677677812
transform 1 0 236 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4336
timestamp 1677677812
transform 1 0 284 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4865
timestamp 1677677812
transform 1 0 284 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4775
timestamp 1677677812
transform 1 0 308 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4776
timestamp 1677677812
transform 1 0 324 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4337
timestamp 1677677812
transform 1 0 332 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4866
timestamp 1677677812
transform 1 0 300 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4867
timestamp 1677677812
transform 1 0 316 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4868
timestamp 1677677812
transform 1 0 332 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4373
timestamp 1677677812
transform 1 0 300 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4374
timestamp 1677677812
transform 1 0 316 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4395
timestamp 1677677812
transform 1 0 308 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4396
timestamp 1677677812
transform 1 0 340 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4293
timestamp 1677677812
transform 1 0 412 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4338
timestamp 1677677812
transform 1 0 364 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4294
timestamp 1677677812
transform 1 0 452 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4777
timestamp 1677677812
transform 1 0 412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4778
timestamp 1677677812
transform 1 0 444 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4779
timestamp 1677677812
transform 1 0 452 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4869
timestamp 1677677812
transform 1 0 364 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4397
timestamp 1677677812
transform 1 0 444 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4295
timestamp 1677677812
transform 1 0 484 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4780
timestamp 1677677812
transform 1 0 476 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4353
timestamp 1677677812
transform 1 0 476 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4870
timestamp 1677677812
transform 1 0 484 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4296
timestamp 1677677812
transform 1 0 516 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4781
timestamp 1677677812
transform 1 0 516 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4871
timestamp 1677677812
transform 1 0 500 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4398
timestamp 1677677812
transform 1 0 500 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4782
timestamp 1677677812
transform 1 0 540 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4375
timestamp 1677677812
transform 1 0 532 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4872
timestamp 1677677812
transform 1 0 548 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4942
timestamp 1677677812
transform 1 0 540 0 1 2395
box -2 -2 2 2
use M2_M1  M2_M1_4783
timestamp 1677677812
transform 1 0 564 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4297
timestamp 1677677812
transform 1 0 612 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4784
timestamp 1677677812
transform 1 0 612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4785
timestamp 1677677812
transform 1 0 620 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4873
timestamp 1677677812
transform 1 0 612 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4339
timestamp 1677677812
transform 1 0 628 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4874
timestamp 1677677812
transform 1 0 628 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4249
timestamp 1677677812
transform 1 0 652 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4786
timestamp 1677677812
transform 1 0 660 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4787
timestamp 1677677812
transform 1 0 716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4788
timestamp 1677677812
transform 1 0 764 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4789
timestamp 1677677812
transform 1 0 772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4875
timestamp 1677677812
transform 1 0 652 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4876
timestamp 1677677812
transform 1 0 668 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4877
timestamp 1677677812
transform 1 0 684 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4376
timestamp 1677677812
transform 1 0 668 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4878
timestamp 1677677812
transform 1 0 772 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4263
timestamp 1677677812
transform 1 0 836 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4790
timestamp 1677677812
transform 1 0 820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4879
timestamp 1677677812
transform 1 0 812 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4399
timestamp 1677677812
transform 1 0 804 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4354
timestamp 1677677812
transform 1 0 828 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4298
timestamp 1677677812
transform 1 0 844 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4880
timestamp 1677677812
transform 1 0 844 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4400
timestamp 1677677812
transform 1 0 876 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4264
timestamp 1677677812
transform 1 0 900 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4401
timestamp 1677677812
transform 1 0 908 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4250
timestamp 1677677812
transform 1 0 948 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4265
timestamp 1677677812
transform 1 0 1060 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4759
timestamp 1677677812
transform 1 0 1124 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4881
timestamp 1677677812
transform 1 0 1140 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4299
timestamp 1677677812
transform 1 0 1164 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4791
timestamp 1677677812
transform 1 0 1164 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4233
timestamp 1677677812
transform 1 0 1188 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4234
timestamp 1677677812
transform 1 0 1220 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4266
timestamp 1677677812
transform 1 0 1180 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4300
timestamp 1677677812
transform 1 0 1212 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4792
timestamp 1677677812
transform 1 0 1212 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4793
timestamp 1677677812
transform 1 0 1260 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4882
timestamp 1677677812
transform 1 0 1180 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4760
timestamp 1677677812
transform 1 0 1284 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4340
timestamp 1677677812
transform 1 0 1284 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4883
timestamp 1677677812
transform 1 0 1276 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4402
timestamp 1677677812
transform 1 0 1276 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4267
timestamp 1677677812
transform 1 0 1324 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4794
timestamp 1677677812
transform 1 0 1324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4884
timestamp 1677677812
transform 1 0 1380 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4268
timestamp 1677677812
transform 1 0 1404 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4761
timestamp 1677677812
transform 1 0 1388 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4341
timestamp 1677677812
transform 1 0 1388 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4795
timestamp 1677677812
transform 1 0 1404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4885
timestamp 1677677812
transform 1 0 1388 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4403
timestamp 1677677812
transform 1 0 1380 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4235
timestamp 1677677812
transform 1 0 1436 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4269
timestamp 1677677812
transform 1 0 1452 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4886
timestamp 1677677812
transform 1 0 1484 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4796
timestamp 1677677812
transform 1 0 1524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4797
timestamp 1677677812
transform 1 0 1540 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4798
timestamp 1677677812
transform 1 0 1556 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4887
timestamp 1677677812
transform 1 0 1532 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4888
timestamp 1677677812
transform 1 0 1548 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4404
timestamp 1677677812
transform 1 0 1540 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4270
timestamp 1677677812
transform 1 0 1572 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4241
timestamp 1677677812
transform 1 0 1588 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4889
timestamp 1677677812
transform 1 0 1588 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4799
timestamp 1677677812
transform 1 0 1604 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4405
timestamp 1677677812
transform 1 0 1612 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4271
timestamp 1677677812
transform 1 0 1628 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4800
timestamp 1677677812
transform 1 0 1668 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4890
timestamp 1677677812
transform 1 0 1628 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4406
timestamp 1677677812
transform 1 0 1644 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4801
timestamp 1677677812
transform 1 0 1740 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4407
timestamp 1677677812
transform 1 0 1764 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4272
timestamp 1677677812
transform 1 0 1780 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4802
timestamp 1677677812
transform 1 0 1788 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4251
timestamp 1677677812
transform 1 0 1820 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4273
timestamp 1677677812
transform 1 0 1812 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4301
timestamp 1677677812
transform 1 0 1804 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4274
timestamp 1677677812
transform 1 0 1828 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4891
timestamp 1677677812
transform 1 0 1820 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4408
timestamp 1677677812
transform 1 0 1812 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4302
timestamp 1677677812
transform 1 0 1892 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4803
timestamp 1677677812
transform 1 0 1892 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4804
timestamp 1677677812
transform 1 0 1908 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4892
timestamp 1677677812
transform 1 0 1884 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4893
timestamp 1677677812
transform 1 0 1900 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4894
timestamp 1677677812
transform 1 0 1932 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4275
timestamp 1677677812
transform 1 0 1972 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4377
timestamp 1677677812
transform 1 0 1964 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4355
timestamp 1677677812
transform 1 0 2020 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4303
timestamp 1677677812
transform 1 0 2092 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4342
timestamp 1677677812
transform 1 0 2068 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4805
timestamp 1677677812
transform 1 0 2092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4895
timestamp 1677677812
transform 1 0 2060 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4896
timestamp 1677677812
transform 1 0 2084 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4897
timestamp 1677677812
transform 1 0 2100 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4409
timestamp 1677677812
transform 1 0 2068 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4410
timestamp 1677677812
transform 1 0 2084 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4276
timestamp 1677677812
transform 1 0 2196 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4236
timestamp 1677677812
transform 1 0 2236 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4237
timestamp 1677677812
transform 1 0 2252 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4277
timestamp 1677677812
transform 1 0 2252 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4806
timestamp 1677677812
transform 1 0 2252 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4898
timestamp 1677677812
transform 1 0 2244 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4356
timestamp 1677677812
transform 1 0 2252 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4304
timestamp 1677677812
transform 1 0 2276 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4807
timestamp 1677677812
transform 1 0 2276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4808
timestamp 1677677812
transform 1 0 2292 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4411
timestamp 1677677812
transform 1 0 2284 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4357
timestamp 1677677812
transform 1 0 2300 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4412
timestamp 1677677812
transform 1 0 2300 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4305
timestamp 1677677812
transform 1 0 2332 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4809
timestamp 1677677812
transform 1 0 2324 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4899
timestamp 1677677812
transform 1 0 2332 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4943
timestamp 1677677812
transform 1 0 2340 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4278
timestamp 1677677812
transform 1 0 2396 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4306
timestamp 1677677812
transform 1 0 2404 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4252
timestamp 1677677812
transform 1 0 2444 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4279
timestamp 1677677812
transform 1 0 2492 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4307
timestamp 1677677812
transform 1 0 2444 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4810
timestamp 1677677812
transform 1 0 2404 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4811
timestamp 1677677812
transform 1 0 2412 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4812
timestamp 1677677812
transform 1 0 2444 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4358
timestamp 1677677812
transform 1 0 2404 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4359
timestamp 1677677812
transform 1 0 2460 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4900
timestamp 1677677812
transform 1 0 2492 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4378
timestamp 1677677812
transform 1 0 2492 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4238
timestamp 1677677812
transform 1 0 2508 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4813
timestamp 1677677812
transform 1 0 2508 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4901
timestamp 1677677812
transform 1 0 2548 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4308
timestamp 1677677812
transform 1 0 2572 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4814
timestamp 1677677812
transform 1 0 2572 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4815
timestamp 1677677812
transform 1 0 2588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4902
timestamp 1677677812
transform 1 0 2564 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4280
timestamp 1677677812
transform 1 0 2628 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4903
timestamp 1677677812
transform 1 0 2628 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4309
timestamp 1677677812
transform 1 0 2644 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4904
timestamp 1677677812
transform 1 0 2644 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4310
timestamp 1677677812
transform 1 0 2684 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4816
timestamp 1677677812
transform 1 0 2684 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4311
timestamp 1677677812
transform 1 0 2724 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4817
timestamp 1677677812
transform 1 0 2724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4905
timestamp 1677677812
transform 1 0 2700 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4281
timestamp 1677677812
transform 1 0 2788 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4312
timestamp 1677677812
transform 1 0 2788 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4818
timestamp 1677677812
transform 1 0 2788 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4944
timestamp 1677677812
transform 1 0 2788 0 1 2395
box -2 -2 2 2
use M3_M2  M3_M2_4253
timestamp 1677677812
transform 1 0 2804 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4282
timestamp 1677677812
transform 1 0 2820 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4313
timestamp 1677677812
transform 1 0 2828 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4906
timestamp 1677677812
transform 1 0 2820 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4907
timestamp 1677677812
transform 1 0 2828 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4762
timestamp 1677677812
transform 1 0 2844 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4413
timestamp 1677677812
transform 1 0 2844 0 1 2385
box -3 -3 3 3
use M2_M1  M2_M1_4819
timestamp 1677677812
transform 1 0 2868 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4379
timestamp 1677677812
transform 1 0 2868 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4239
timestamp 1677677812
transform 1 0 2900 0 1 2465
box -3 -3 3 3
use M3_M2  M3_M2_4360
timestamp 1677677812
transform 1 0 2900 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4908
timestamp 1677677812
transform 1 0 2916 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4380
timestamp 1677677812
transform 1 0 2916 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4361
timestamp 1677677812
transform 1 0 2940 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4763
timestamp 1677677812
transform 1 0 2956 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4820
timestamp 1677677812
transform 1 0 2996 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4314
timestamp 1677677812
transform 1 0 3012 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4909
timestamp 1677677812
transform 1 0 3012 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4242
timestamp 1677677812
transform 1 0 3052 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4821
timestamp 1677677812
transform 1 0 3044 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4315
timestamp 1677677812
transform 1 0 3076 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4822
timestamp 1677677812
transform 1 0 3076 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4910
timestamp 1677677812
transform 1 0 3052 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4911
timestamp 1677677812
transform 1 0 3068 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4316
timestamp 1677677812
transform 1 0 3108 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4823
timestamp 1677677812
transform 1 0 3108 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4317
timestamp 1677677812
transform 1 0 3124 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4912
timestamp 1677677812
transform 1 0 3124 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4913
timestamp 1677677812
transform 1 0 3140 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4318
timestamp 1677677812
transform 1 0 3172 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4824
timestamp 1677677812
transform 1 0 3196 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4914
timestamp 1677677812
transform 1 0 3228 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4825
timestamp 1677677812
transform 1 0 3244 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4362
timestamp 1677677812
transform 1 0 3244 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4254
timestamp 1677677812
transform 1 0 3268 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4319
timestamp 1677677812
transform 1 0 3292 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4756
timestamp 1677677812
transform 1 0 3316 0 1 2435
box -2 -2 2 2
use M2_M1  M2_M1_4764
timestamp 1677677812
transform 1 0 3300 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4826
timestamp 1677677812
transform 1 0 3276 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4343
timestamp 1677677812
transform 1 0 3292 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4915
timestamp 1677677812
transform 1 0 3268 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4381
timestamp 1677677812
transform 1 0 3252 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4363
timestamp 1677677812
transform 1 0 3276 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4916
timestamp 1677677812
transform 1 0 3292 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4320
timestamp 1677677812
transform 1 0 3316 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4765
timestamp 1677677812
transform 1 0 3332 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4382
timestamp 1677677812
transform 1 0 3300 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4383
timestamp 1677677812
transform 1 0 3348 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4283
timestamp 1677677812
transform 1 0 3372 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4757
timestamp 1677677812
transform 1 0 3380 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_4321
timestamp 1677677812
transform 1 0 3388 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4827
timestamp 1677677812
transform 1 0 3388 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4766
timestamp 1677677812
transform 1 0 3428 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4284
timestamp 1677677812
transform 1 0 3452 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4322
timestamp 1677677812
transform 1 0 3460 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4828
timestamp 1677677812
transform 1 0 3460 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4829
timestamp 1677677812
transform 1 0 3476 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4917
timestamp 1677677812
transform 1 0 3444 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4918
timestamp 1677677812
transform 1 0 3452 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4364
timestamp 1677677812
transform 1 0 3460 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4243
timestamp 1677677812
transform 1 0 3516 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4830
timestamp 1677677812
transform 1 0 3500 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4344
timestamp 1677677812
transform 1 0 3508 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4919
timestamp 1677677812
transform 1 0 3508 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4831
timestamp 1677677812
transform 1 0 3556 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4345
timestamp 1677677812
transform 1 0 3588 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4832
timestamp 1677677812
transform 1 0 3604 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4920
timestamp 1677677812
transform 1 0 3524 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4365
timestamp 1677677812
transform 1 0 3548 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4384
timestamp 1677677812
transform 1 0 3524 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4244
timestamp 1677677812
transform 1 0 3628 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4285
timestamp 1677677812
transform 1 0 3652 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4833
timestamp 1677677812
transform 1 0 3636 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4834
timestamp 1677677812
transform 1 0 3652 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4921
timestamp 1677677812
transform 1 0 3620 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4922
timestamp 1677677812
transform 1 0 3628 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4414
timestamp 1677677812
transform 1 0 3620 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4366
timestamp 1677677812
transform 1 0 3636 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4245
timestamp 1677677812
transform 1 0 3668 0 1 2455
box -3 -3 3 3
use M2_M1  M2_M1_4923
timestamp 1677677812
transform 1 0 3644 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4924
timestamp 1677677812
transform 1 0 3660 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4385
timestamp 1677677812
transform 1 0 3644 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4415
timestamp 1677677812
transform 1 0 3644 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4367
timestamp 1677677812
transform 1 0 3668 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4925
timestamp 1677677812
transform 1 0 3676 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4246
timestamp 1677677812
transform 1 0 3700 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4323
timestamp 1677677812
transform 1 0 3756 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4346
timestamp 1677677812
transform 1 0 3692 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4347
timestamp 1677677812
transform 1 0 3716 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4835
timestamp 1677677812
transform 1 0 3724 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4926
timestamp 1677677812
transform 1 0 3692 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4386
timestamp 1677677812
transform 1 0 3724 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4416
timestamp 1677677812
transform 1 0 3692 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4417
timestamp 1677677812
transform 1 0 3732 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4286
timestamp 1677677812
transform 1 0 3820 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4836
timestamp 1677677812
transform 1 0 3820 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4837
timestamp 1677677812
transform 1 0 3852 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4927
timestamp 1677677812
transform 1 0 3924 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4255
timestamp 1677677812
transform 1 0 3940 0 1 2445
box -3 -3 3 3
use M2_M1  M2_M1_4838
timestamp 1677677812
transform 1 0 3948 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4839
timestamp 1677677812
transform 1 0 3964 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4928
timestamp 1677677812
transform 1 0 3940 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4929
timestamp 1677677812
transform 1 0 3956 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4387
timestamp 1677677812
transform 1 0 3956 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4840
timestamp 1677677812
transform 1 0 3980 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4930
timestamp 1677677812
transform 1 0 3980 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4324
timestamp 1677677812
transform 1 0 4068 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4841
timestamp 1677677812
transform 1 0 4036 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4368
timestamp 1677677812
transform 1 0 4028 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4842
timestamp 1677677812
transform 1 0 4092 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4931
timestamp 1677677812
transform 1 0 4068 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4932
timestamp 1677677812
transform 1 0 4084 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4388
timestamp 1677677812
transform 1 0 4036 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4389
timestamp 1677677812
transform 1 0 4068 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4369
timestamp 1677677812
transform 1 0 4092 0 1 2405
box -3 -3 3 3
use M2_M1  M2_M1_4843
timestamp 1677677812
transform 1 0 4116 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4325
timestamp 1677677812
transform 1 0 4132 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4256
timestamp 1677677812
transform 1 0 4148 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4326
timestamp 1677677812
transform 1 0 4172 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4844
timestamp 1677677812
transform 1 0 4172 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4327
timestamp 1677677812
transform 1 0 4260 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4328
timestamp 1677677812
transform 1 0 4276 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4845
timestamp 1677677812
transform 1 0 4244 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4846
timestamp 1677677812
transform 1 0 4260 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4348
timestamp 1677677812
transform 1 0 4268 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4847
timestamp 1677677812
transform 1 0 4276 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4933
timestamp 1677677812
transform 1 0 4220 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4934
timestamp 1677677812
transform 1 0 4236 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4935
timestamp 1677677812
transform 1 0 4252 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4936
timestamp 1677677812
transform 1 0 4268 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4937
timestamp 1677677812
transform 1 0 4276 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4349
timestamp 1677677812
transform 1 0 4292 0 1 2415
box -3 -3 3 3
use M2_M1  M2_M1_4767
timestamp 1677677812
transform 1 0 4324 0 1 2425
box -2 -2 2 2
use M3_M2  M3_M2_4370
timestamp 1677677812
transform 1 0 4316 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4240
timestamp 1677677812
transform 1 0 4340 0 1 2465
box -3 -3 3 3
use M2_M1  M2_M1_4758
timestamp 1677677812
transform 1 0 4340 0 1 2435
box -2 -2 2 2
use M3_M2  M3_M2_4287
timestamp 1677677812
transform 1 0 4348 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4329
timestamp 1677677812
transform 1 0 4340 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4768
timestamp 1677677812
transform 1 0 4364 0 1 2425
box -2 -2 2 2
use M2_M1  M2_M1_4848
timestamp 1677677812
transform 1 0 4348 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4350
timestamp 1677677812
transform 1 0 4356 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4351
timestamp 1677677812
transform 1 0 4380 0 1 2415
box -3 -3 3 3
use M3_M2  M3_M2_4257
timestamp 1677677812
transform 1 0 4476 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4258
timestamp 1677677812
transform 1 0 4524 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4330
timestamp 1677677812
transform 1 0 4524 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4849
timestamp 1677677812
transform 1 0 4428 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4850
timestamp 1677677812
transform 1 0 4460 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4851
timestamp 1677677812
transform 1 0 4524 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4938
timestamp 1677677812
transform 1 0 4380 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4390
timestamp 1677677812
transform 1 0 4380 0 1 2395
box -3 -3 3 3
use M2_M1  M2_M1_4939
timestamp 1677677812
transform 1 0 4476 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4418
timestamp 1677677812
transform 1 0 4468 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4331
timestamp 1677677812
transform 1 0 4572 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4332
timestamp 1677677812
transform 1 0 4588 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4247
timestamp 1677677812
transform 1 0 4604 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4288
timestamp 1677677812
transform 1 0 4612 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4333
timestamp 1677677812
transform 1 0 4620 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4852
timestamp 1677677812
transform 1 0 4580 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4853
timestamp 1677677812
transform 1 0 4588 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4854
timestamp 1677677812
transform 1 0 4596 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4855
timestamp 1677677812
transform 1 0 4612 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4856
timestamp 1677677812
transform 1 0 4628 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4391
timestamp 1677677812
transform 1 0 4580 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4392
timestamp 1677677812
transform 1 0 4596 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4419
timestamp 1677677812
transform 1 0 4588 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4420
timestamp 1677677812
transform 1 0 4628 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4248
timestamp 1677677812
transform 1 0 4644 0 1 2455
box -3 -3 3 3
use M3_M2  M3_M2_4259
timestamp 1677677812
transform 1 0 4644 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4260
timestamp 1677677812
transform 1 0 4660 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4261
timestamp 1677677812
transform 1 0 4676 0 1 2445
box -3 -3 3 3
use M3_M2  M3_M2_4289
timestamp 1677677812
transform 1 0 4668 0 1 2435
box -3 -3 3 3
use M2_M1  M2_M1_4857
timestamp 1677677812
transform 1 0 4660 0 1 2415
box -2 -2 2 2
use M3_M2  M3_M2_4290
timestamp 1677677812
transform 1 0 4716 0 1 2435
box -3 -3 3 3
use M3_M2  M3_M2_4334
timestamp 1677677812
transform 1 0 4676 0 1 2425
box -3 -3 3 3
use M3_M2  M3_M2_4335
timestamp 1677677812
transform 1 0 4772 0 1 2425
box -3 -3 3 3
use M2_M1  M2_M1_4858
timestamp 1677677812
transform 1 0 4716 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4859
timestamp 1677677812
transform 1 0 4772 0 1 2415
box -2 -2 2 2
use M2_M1  M2_M1_4940
timestamp 1677677812
transform 1 0 4676 0 1 2405
box -2 -2 2 2
use M2_M1  M2_M1_4941
timestamp 1677677812
transform 1 0 4692 0 1 2405
box -2 -2 2 2
use M3_M2  M3_M2_4371
timestamp 1677677812
transform 1 0 4716 0 1 2405
box -3 -3 3 3
use M3_M2  M3_M2_4393
timestamp 1677677812
transform 1 0 4708 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4394
timestamp 1677677812
transform 1 0 4724 0 1 2395
box -3 -3 3 3
use M3_M2  M3_M2_4421
timestamp 1677677812
transform 1 0 4692 0 1 2385
box -3 -3 3 3
use M3_M2  M3_M2_4422
timestamp 1677677812
transform 1 0 4756 0 1 2385
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_46
timestamp 1677677812
transform 1 0 48 0 1 2370
box -10 -3 10 3
use M3_M2  M3_M2_4423
timestamp 1677677812
transform 1 0 84 0 1 2375
box -3 -3 3 3
use FILL  FILL_5387
timestamp 1677677812
transform 1 0 72 0 1 2370
box -8 -3 16 105
use FILL  FILL_5388
timestamp 1677677812
transform 1 0 80 0 1 2370
box -8 -3 16 105
use FILL  FILL_5389
timestamp 1677677812
transform 1 0 88 0 1 2370
box -8 -3 16 105
use FILL  FILL_5390
timestamp 1677677812
transform 1 0 96 0 1 2370
box -8 -3 16 105
use FILL  FILL_5391
timestamp 1677677812
transform 1 0 104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5392
timestamp 1677677812
transform 1 0 112 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_364
timestamp 1677677812
transform -1 0 136 0 1 2370
box -9 -3 26 105
use FILL  FILL_5393
timestamp 1677677812
transform 1 0 136 0 1 2370
box -8 -3 16 105
use FILL  FILL_5394
timestamp 1677677812
transform 1 0 144 0 1 2370
box -8 -3 16 105
use FILL  FILL_5395
timestamp 1677677812
transform 1 0 152 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_221
timestamp 1677677812
transform -1 0 200 0 1 2370
box -8 -3 46 105
use FILL  FILL_5396
timestamp 1677677812
transform 1 0 200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5397
timestamp 1677677812
transform 1 0 208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5398
timestamp 1677677812
transform 1 0 216 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_222
timestamp 1677677812
transform 1 0 224 0 1 2370
box -8 -3 46 105
use FILL  FILL_5399
timestamp 1677677812
transform 1 0 264 0 1 2370
box -8 -3 16 105
use FILL  FILL_5401
timestamp 1677677812
transform 1 0 272 0 1 2370
box -8 -3 16 105
use FILL  FILL_5403
timestamp 1677677812
transform 1 0 280 0 1 2370
box -8 -3 16 105
use FILL  FILL_5405
timestamp 1677677812
transform 1 0 288 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_210
timestamp 1677677812
transform -1 0 336 0 1 2370
box -8 -3 46 105
use FILL  FILL_5406
timestamp 1677677812
transform 1 0 336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5407
timestamp 1677677812
transform 1 0 344 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4424
timestamp 1677677812
transform 1 0 364 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_316
timestamp 1677677812
transform 1 0 352 0 1 2370
box -8 -3 104 105
use FILL  FILL_5408
timestamp 1677677812
transform 1 0 448 0 1 2370
box -8 -3 16 105
use FILL  FILL_5409
timestamp 1677677812
transform 1 0 456 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_366
timestamp 1677677812
transform -1 0 480 0 1 2370
box -9 -3 26 105
use FILL  FILL_5410
timestamp 1677677812
transform 1 0 480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5411
timestamp 1677677812
transform 1 0 488 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4425
timestamp 1677677812
transform 1 0 508 0 1 2375
box -3 -3 3 3
use AOI22X1  AOI22X1_225
timestamp 1677677812
transform -1 0 536 0 1 2370
box -8 -3 46 105
use M3_M2  M3_M2_4426
timestamp 1677677812
transform 1 0 548 0 1 2375
box -3 -3 3 3
use FILL  FILL_5412
timestamp 1677677812
transform 1 0 536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5413
timestamp 1677677812
transform 1 0 544 0 1 2370
box -8 -3 16 105
use FILL  FILL_5414
timestamp 1677677812
transform 1 0 552 0 1 2370
box -8 -3 16 105
use FILL  FILL_5415
timestamp 1677677812
transform 1 0 560 0 1 2370
box -8 -3 16 105
use FILL  FILL_5416
timestamp 1677677812
transform 1 0 568 0 1 2370
box -8 -3 16 105
use FILL  FILL_5426
timestamp 1677677812
transform 1 0 576 0 1 2370
box -8 -3 16 105
use FILL  FILL_5428
timestamp 1677677812
transform 1 0 584 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4427
timestamp 1677677812
transform 1 0 612 0 1 2375
box -3 -3 3 3
use NOR2X1  NOR2X1_54
timestamp 1677677812
transform 1 0 592 0 1 2370
box -8 -3 32 105
use FILL  FILL_5430
timestamp 1677677812
transform 1 0 616 0 1 2370
box -8 -3 16 105
use FILL  FILL_5431
timestamp 1677677812
transform 1 0 624 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_212
timestamp 1677677812
transform 1 0 632 0 1 2370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_318
timestamp 1677677812
transform 1 0 672 0 1 2370
box -8 -3 104 105
use FILL  FILL_5432
timestamp 1677677812
transform 1 0 768 0 1 2370
box -8 -3 16 105
use FILL  FILL_5433
timestamp 1677677812
transform 1 0 776 0 1 2370
box -8 -3 16 105
use FILL  FILL_5440
timestamp 1677677812
transform 1 0 784 0 1 2370
box -8 -3 16 105
use FILL  FILL_5442
timestamp 1677677812
transform 1 0 792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5444
timestamp 1677677812
transform 1 0 800 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_108
timestamp 1677677812
transform 1 0 808 0 1 2370
box -8 -3 34 105
use FILL  FILL_5446
timestamp 1677677812
transform 1 0 840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5447
timestamp 1677677812
transform 1 0 848 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4428
timestamp 1677677812
transform 1 0 868 0 1 2375
box -3 -3 3 3
use FILL  FILL_5448
timestamp 1677677812
transform 1 0 856 0 1 2370
box -8 -3 16 105
use FILL  FILL_5452
timestamp 1677677812
transform 1 0 864 0 1 2370
box -8 -3 16 105
use FILL  FILL_5454
timestamp 1677677812
transform 1 0 872 0 1 2370
box -8 -3 16 105
use FILL  FILL_5456
timestamp 1677677812
transform 1 0 880 0 1 2370
box -8 -3 16 105
use FILL  FILL_5458
timestamp 1677677812
transform 1 0 888 0 1 2370
box -8 -3 16 105
use FILL  FILL_5460
timestamp 1677677812
transform 1 0 896 0 1 2370
box -8 -3 16 105
use FILL  FILL_5462
timestamp 1677677812
transform 1 0 904 0 1 2370
box -8 -3 16 105
use FILL  FILL_5464
timestamp 1677677812
transform 1 0 912 0 1 2370
box -8 -3 16 105
use FILL  FILL_5465
timestamp 1677677812
transform 1 0 920 0 1 2370
box -8 -3 16 105
use FILL  FILL_5466
timestamp 1677677812
transform 1 0 928 0 1 2370
box -8 -3 16 105
use FILL  FILL_5467
timestamp 1677677812
transform 1 0 936 0 1 2370
box -8 -3 16 105
use FILL  FILL_5468
timestamp 1677677812
transform 1 0 944 0 1 2370
box -8 -3 16 105
use FILL  FILL_5469
timestamp 1677677812
transform 1 0 952 0 1 2370
box -8 -3 16 105
use FILL  FILL_5471
timestamp 1677677812
transform 1 0 960 0 1 2370
box -8 -3 16 105
use FILL  FILL_5473
timestamp 1677677812
transform 1 0 968 0 1 2370
box -8 -3 16 105
use FILL  FILL_5475
timestamp 1677677812
transform 1 0 976 0 1 2370
box -8 -3 16 105
use FILL  FILL_5477
timestamp 1677677812
transform 1 0 984 0 1 2370
box -8 -3 16 105
use FILL  FILL_5479
timestamp 1677677812
transform 1 0 992 0 1 2370
box -8 -3 16 105
use FILL  FILL_5481
timestamp 1677677812
transform 1 0 1000 0 1 2370
box -8 -3 16 105
use FILL  FILL_5483
timestamp 1677677812
transform 1 0 1008 0 1 2370
box -8 -3 16 105
use FILL  FILL_5485
timestamp 1677677812
transform 1 0 1016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5487
timestamp 1677677812
transform 1 0 1024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5489
timestamp 1677677812
transform 1 0 1032 0 1 2370
box -8 -3 16 105
use FILL  FILL_5490
timestamp 1677677812
transform 1 0 1040 0 1 2370
box -8 -3 16 105
use FILL  FILL_5491
timestamp 1677677812
transform 1 0 1048 0 1 2370
box -8 -3 16 105
use FILL  FILL_5492
timestamp 1677677812
transform 1 0 1056 0 1 2370
box -8 -3 16 105
use FILL  FILL_5493
timestamp 1677677812
transform 1 0 1064 0 1 2370
box -8 -3 16 105
use FILL  FILL_5494
timestamp 1677677812
transform 1 0 1072 0 1 2370
box -8 -3 16 105
use FILL  FILL_5495
timestamp 1677677812
transform 1 0 1080 0 1 2370
box -8 -3 16 105
use FILL  FILL_5496
timestamp 1677677812
transform 1 0 1088 0 1 2370
box -8 -3 16 105
use FILL  FILL_5497
timestamp 1677677812
transform 1 0 1096 0 1 2370
box -8 -3 16 105
use FILL  FILL_5498
timestamp 1677677812
transform 1 0 1104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5499
timestamp 1677677812
transform 1 0 1112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5500
timestamp 1677677812
transform 1 0 1120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5501
timestamp 1677677812
transform 1 0 1128 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4429
timestamp 1677677812
transform 1 0 1164 0 1 2375
box -3 -3 3 3
use INVX2  INVX2_368
timestamp 1677677812
transform 1 0 1136 0 1 2370
box -9 -3 26 105
use FILL  FILL_5503
timestamp 1677677812
transform 1 0 1152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5504
timestamp 1677677812
transform 1 0 1160 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4430
timestamp 1677677812
transform 1 0 1260 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_321
timestamp 1677677812
transform 1 0 1168 0 1 2370
box -8 -3 104 105
use FILL  FILL_5505
timestamp 1677677812
transform 1 0 1264 0 1 2370
box -8 -3 16 105
use FILL  FILL_5516
timestamp 1677677812
transform 1 0 1272 0 1 2370
box -8 -3 16 105
use FILL  FILL_5518
timestamp 1677677812
transform 1 0 1280 0 1 2370
box -8 -3 16 105
use FILL  FILL_5520
timestamp 1677677812
transform 1 0 1288 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_110
timestamp 1677677812
transform -1 0 1328 0 1 2370
box -8 -3 34 105
use FILL  FILL_5522
timestamp 1677677812
transform 1 0 1328 0 1 2370
box -8 -3 16 105
use FILL  FILL_5524
timestamp 1677677812
transform 1 0 1336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5526
timestamp 1677677812
transform 1 0 1344 0 1 2370
box -8 -3 16 105
use FILL  FILL_5528
timestamp 1677677812
transform 1 0 1352 0 1 2370
box -8 -3 16 105
use FILL  FILL_5530
timestamp 1677677812
transform 1 0 1360 0 1 2370
box -8 -3 16 105
use FILL  FILL_5532
timestamp 1677677812
transform 1 0 1368 0 1 2370
box -8 -3 16 105
use FILL  FILL_5534
timestamp 1677677812
transform 1 0 1376 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_112
timestamp 1677677812
transform -1 0 1416 0 1 2370
box -8 -3 34 105
use FILL  FILL_5535
timestamp 1677677812
transform 1 0 1416 0 1 2370
box -8 -3 16 105
use FILL  FILL_5536
timestamp 1677677812
transform 1 0 1424 0 1 2370
box -8 -3 16 105
use FILL  FILL_5537
timestamp 1677677812
transform 1 0 1432 0 1 2370
box -8 -3 16 105
use FILL  FILL_5538
timestamp 1677677812
transform 1 0 1440 0 1 2370
box -8 -3 16 105
use FILL  FILL_5539
timestamp 1677677812
transform 1 0 1448 0 1 2370
box -8 -3 16 105
use FILL  FILL_5540
timestamp 1677677812
transform 1 0 1456 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_370
timestamp 1677677812
transform -1 0 1480 0 1 2370
box -9 -3 26 105
use FILL  FILL_5541
timestamp 1677677812
transform 1 0 1480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5544
timestamp 1677677812
transform 1 0 1488 0 1 2370
box -8 -3 16 105
use FILL  FILL_5546
timestamp 1677677812
transform 1 0 1496 0 1 2370
box -8 -3 16 105
use FILL  FILL_5548
timestamp 1677677812
transform 1 0 1504 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4431
timestamp 1677677812
transform 1 0 1532 0 1 2375
box -3 -3 3 3
use FILL  FILL_5550
timestamp 1677677812
transform 1 0 1512 0 1 2370
box -8 -3 16 105
use FILL  FILL_5552
timestamp 1677677812
transform 1 0 1520 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_213
timestamp 1677677812
transform -1 0 1568 0 1 2370
box -8 -3 46 105
use M3_M2  M3_M2_4432
timestamp 1677677812
transform 1 0 1580 0 1 2375
box -3 -3 3 3
use FILL  FILL_5554
timestamp 1677677812
transform 1 0 1568 0 1 2370
box -8 -3 16 105
use FILL  FILL_5556
timestamp 1677677812
transform 1 0 1576 0 1 2370
box -8 -3 16 105
use FILL  FILL_5558
timestamp 1677677812
transform 1 0 1584 0 1 2370
box -8 -3 16 105
use FILL  FILL_5560
timestamp 1677677812
transform 1 0 1592 0 1 2370
box -8 -3 16 105
use FILL  FILL_5562
timestamp 1677677812
transform 1 0 1600 0 1 2370
box -8 -3 16 105
use FILL  FILL_5564
timestamp 1677677812
transform 1 0 1608 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4433
timestamp 1677677812
transform 1 0 1684 0 1 2375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_323
timestamp 1677677812
transform 1 0 1616 0 1 2370
box -8 -3 104 105
use FILL  FILL_5566
timestamp 1677677812
transform 1 0 1712 0 1 2370
box -8 -3 16 105
use FILL  FILL_5575
timestamp 1677677812
transform 1 0 1720 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_371
timestamp 1677677812
transform 1 0 1728 0 1 2370
box -9 -3 26 105
use FILL  FILL_5577
timestamp 1677677812
transform 1 0 1744 0 1 2370
box -8 -3 16 105
use FILL  FILL_5578
timestamp 1677677812
transform 1 0 1752 0 1 2370
box -8 -3 16 105
use FILL  FILL_5579
timestamp 1677677812
transform 1 0 1760 0 1 2370
box -8 -3 16 105
use FILL  FILL_5580
timestamp 1677677812
transform 1 0 1768 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4434
timestamp 1677677812
transform 1 0 1788 0 1 2375
box -3 -3 3 3
use FILL  FILL_5581
timestamp 1677677812
transform 1 0 1776 0 1 2370
box -8 -3 16 105
use FILL  FILL_5582
timestamp 1677677812
transform 1 0 1784 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_51
timestamp 1677677812
transform 1 0 1792 0 1 2370
box -5 -3 28 105
use FILL  FILL_5583
timestamp 1677677812
transform 1 0 1816 0 1 2370
box -8 -3 16 105
use FILL  FILL_5584
timestamp 1677677812
transform 1 0 1824 0 1 2370
box -8 -3 16 105
use FILL  FILL_5585
timestamp 1677677812
transform 1 0 1832 0 1 2370
box -8 -3 16 105
use FILL  FILL_5588
timestamp 1677677812
transform 1 0 1840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5590
timestamp 1677677812
transform 1 0 1848 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4435
timestamp 1677677812
transform 1 0 1868 0 1 2375
box -3 -3 3 3
use FILL  FILL_5592
timestamp 1677677812
transform 1 0 1856 0 1 2370
box -8 -3 16 105
use FILL  FILL_5594
timestamp 1677677812
transform 1 0 1864 0 1 2370
box -8 -3 16 105
use FILL  FILL_5595
timestamp 1677677812
transform 1 0 1872 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4436
timestamp 1677677812
transform 1 0 1900 0 1 2375
box -3 -3 3 3
use OAI22X1  OAI22X1_216
timestamp 1677677812
transform -1 0 1920 0 1 2370
box -8 -3 46 105
use FILL  FILL_5596
timestamp 1677677812
transform 1 0 1920 0 1 2370
box -8 -3 16 105
use FILL  FILL_5597
timestamp 1677677812
transform 1 0 1928 0 1 2370
box -8 -3 16 105
use FILL  FILL_5598
timestamp 1677677812
transform 1 0 1936 0 1 2370
box -8 -3 16 105
use FILL  FILL_5599
timestamp 1677677812
transform 1 0 1944 0 1 2370
box -8 -3 16 105
use FILL  FILL_5600
timestamp 1677677812
transform 1 0 1952 0 1 2370
box -8 -3 16 105
use FILL  FILL_5601
timestamp 1677677812
transform 1 0 1960 0 1 2370
box -8 -3 16 105
use FILL  FILL_5602
timestamp 1677677812
transform 1 0 1968 0 1 2370
box -8 -3 16 105
use FILL  FILL_5603
timestamp 1677677812
transform 1 0 1976 0 1 2370
box -8 -3 16 105
use FILL  FILL_5604
timestamp 1677677812
transform 1 0 1984 0 1 2370
box -8 -3 16 105
use FILL  FILL_5605
timestamp 1677677812
transform 1 0 1992 0 1 2370
box -8 -3 16 105
use FILL  FILL_5606
timestamp 1677677812
transform 1 0 2000 0 1 2370
box -8 -3 16 105
use FILL  FILL_5607
timestamp 1677677812
transform 1 0 2008 0 1 2370
box -8 -3 16 105
use FILL  FILL_5608
timestamp 1677677812
transform 1 0 2016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5609
timestamp 1677677812
transform 1 0 2024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5610
timestamp 1677677812
transform 1 0 2032 0 1 2370
box -8 -3 16 105
use FILL  FILL_5611
timestamp 1677677812
transform 1 0 2040 0 1 2370
box -8 -3 16 105
use FILL  FILL_5612
timestamp 1677677812
transform 1 0 2048 0 1 2370
box -8 -3 16 105
use FILL  FILL_5613
timestamp 1677677812
transform 1 0 2056 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_217
timestamp 1677677812
transform 1 0 2064 0 1 2370
box -8 -3 46 105
use FILL  FILL_5614
timestamp 1677677812
transform 1 0 2104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5625
timestamp 1677677812
transform 1 0 2112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5627
timestamp 1677677812
transform 1 0 2120 0 1 2370
box -8 -3 16 105
use FILL  FILL_5629
timestamp 1677677812
transform 1 0 2128 0 1 2370
box -8 -3 16 105
use FILL  FILL_5631
timestamp 1677677812
transform 1 0 2136 0 1 2370
box -8 -3 16 105
use FILL  FILL_5633
timestamp 1677677812
transform 1 0 2144 0 1 2370
box -8 -3 16 105
use FILL  FILL_5635
timestamp 1677677812
transform 1 0 2152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5636
timestamp 1677677812
transform 1 0 2160 0 1 2370
box -8 -3 16 105
use FILL  FILL_5637
timestamp 1677677812
transform 1 0 2168 0 1 2370
box -8 -3 16 105
use FILL  FILL_5638
timestamp 1677677812
transform 1 0 2176 0 1 2370
box -8 -3 16 105
use FILL  FILL_5639
timestamp 1677677812
transform 1 0 2184 0 1 2370
box -8 -3 16 105
use FILL  FILL_5640
timestamp 1677677812
transform 1 0 2192 0 1 2370
box -8 -3 16 105
use FILL  FILL_5641
timestamp 1677677812
transform 1 0 2200 0 1 2370
box -8 -3 16 105
use FILL  FILL_5644
timestamp 1677677812
transform 1 0 2208 0 1 2370
box -8 -3 16 105
use FILL  FILL_5646
timestamp 1677677812
transform 1 0 2216 0 1 2370
box -8 -3 16 105
use FILL  FILL_5648
timestamp 1677677812
transform 1 0 2224 0 1 2370
box -8 -3 16 105
use FILL  FILL_5650
timestamp 1677677812
transform 1 0 2232 0 1 2370
box -8 -3 16 105
use FILL  FILL_5652
timestamp 1677677812
transform 1 0 2240 0 1 2370
box -8 -3 16 105
use FILL  FILL_5654
timestamp 1677677812
transform 1 0 2248 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_231
timestamp 1677677812
transform 1 0 2256 0 1 2370
box -8 -3 46 105
use FILL  FILL_5656
timestamp 1677677812
transform 1 0 2296 0 1 2370
box -8 -3 16 105
use FILL  FILL_5660
timestamp 1677677812
transform 1 0 2304 0 1 2370
box -8 -3 16 105
use FILL  FILL_5662
timestamp 1677677812
transform 1 0 2312 0 1 2370
box -8 -3 16 105
use FILL  FILL_5664
timestamp 1677677812
transform 1 0 2320 0 1 2370
box -8 -3 16 105
use FILL  FILL_5666
timestamp 1677677812
transform 1 0 2328 0 1 2370
box -8 -3 16 105
use FILL  FILL_5668
timestamp 1677677812
transform 1 0 2336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5669
timestamp 1677677812
transform 1 0 2344 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_374
timestamp 1677677812
transform 1 0 2352 0 1 2370
box -9 -3 26 105
use FILL  FILL_5670
timestamp 1677677812
transform 1 0 2368 0 1 2370
box -8 -3 16 105
use FILL  FILL_5671
timestamp 1677677812
transform 1 0 2376 0 1 2370
box -8 -3 16 105
use FILL  FILL_5673
timestamp 1677677812
transform 1 0 2384 0 1 2370
box -8 -3 16 105
use FILL  FILL_5675
timestamp 1677677812
transform 1 0 2392 0 1 2370
box -8 -3 16 105
use FILL  FILL_5677
timestamp 1677677812
transform 1 0 2400 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_326
timestamp 1677677812
transform -1 0 2504 0 1 2370
box -8 -3 104 105
use FILL  FILL_5678
timestamp 1677677812
transform 1 0 2504 0 1 2370
box -8 -3 16 105
use FILL  FILL_5679
timestamp 1677677812
transform 1 0 2512 0 1 2370
box -8 -3 16 105
use FILL  FILL_5680
timestamp 1677677812
transform 1 0 2520 0 1 2370
box -8 -3 16 105
use FILL  FILL_5681
timestamp 1677677812
transform 1 0 2528 0 1 2370
box -8 -3 16 105
use FILL  FILL_5687
timestamp 1677677812
transform 1 0 2536 0 1 2370
box -8 -3 16 105
use FILL  FILL_5689
timestamp 1677677812
transform 1 0 2544 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_233
timestamp 1677677812
transform 1 0 2552 0 1 2370
box -8 -3 46 105
use FILL  FILL_5691
timestamp 1677677812
transform 1 0 2592 0 1 2370
box -8 -3 16 105
use FILL  FILL_5698
timestamp 1677677812
transform 1 0 2600 0 1 2370
box -8 -3 16 105
use FILL  FILL_5700
timestamp 1677677812
transform 1 0 2608 0 1 2370
box -8 -3 16 105
use FILL  FILL_5702
timestamp 1677677812
transform 1 0 2616 0 1 2370
box -8 -3 16 105
use FILL  FILL_5704
timestamp 1677677812
transform 1 0 2624 0 1 2370
box -8 -3 16 105
use FILL  FILL_5706
timestamp 1677677812
transform 1 0 2632 0 1 2370
box -8 -3 16 105
use FILL  FILL_5708
timestamp 1677677812
transform 1 0 2640 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_375
timestamp 1677677812
transform 1 0 2648 0 1 2370
box -9 -3 26 105
use FILL  FILL_5710
timestamp 1677677812
transform 1 0 2664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5712
timestamp 1677677812
transform 1 0 2672 0 1 2370
box -8 -3 16 105
use FILL  FILL_5714
timestamp 1677677812
transform 1 0 2680 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_328
timestamp 1677677812
transform 1 0 2688 0 1 2370
box -8 -3 104 105
use FILL  FILL_5716
timestamp 1677677812
transform 1 0 2784 0 1 2370
box -8 -3 16 105
use FILL  FILL_5718
timestamp 1677677812
transform 1 0 2792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5720
timestamp 1677677812
transform 1 0 2800 0 1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_56
timestamp 1677677812
transform 1 0 2808 0 1 2370
box -8 -3 32 105
use FILL  FILL_5722
timestamp 1677677812
transform 1 0 2832 0 1 2370
box -8 -3 16 105
use FILL  FILL_5723
timestamp 1677677812
transform 1 0 2840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5724
timestamp 1677677812
transform 1 0 2848 0 1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4437
timestamp 1677677812
transform 1 0 2868 0 1 2375
box -3 -3 3 3
use FILL  FILL_5725
timestamp 1677677812
transform 1 0 2856 0 1 2370
box -8 -3 16 105
use FILL  FILL_5726
timestamp 1677677812
transform 1 0 2864 0 1 2370
box -8 -3 16 105
use FILL  FILL_5731
timestamp 1677677812
transform 1 0 2872 0 1 2370
box -8 -3 16 105
use FILL  FILL_5733
timestamp 1677677812
transform 1 0 2880 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_114
timestamp 1677677812
transform 1 0 2888 0 1 2370
box -8 -3 34 105
use FILL  FILL_5735
timestamp 1677677812
transform 1 0 2920 0 1 2370
box -8 -3 16 105
use FILL  FILL_5736
timestamp 1677677812
transform 1 0 2928 0 1 2370
box -8 -3 16 105
use FILL  FILL_5740
timestamp 1677677812
transform 1 0 2936 0 1 2370
box -8 -3 16 105
use FILL  FILL_5742
timestamp 1677677812
transform 1 0 2944 0 1 2370
box -8 -3 16 105
use FILL  FILL_5744
timestamp 1677677812
transform 1 0 2952 0 1 2370
box -8 -3 16 105
use FILL  FILL_5746
timestamp 1677677812
transform 1 0 2960 0 1 2370
box -8 -3 16 105
use FILL  FILL_5748
timestamp 1677677812
transform 1 0 2968 0 1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_115
timestamp 1677677812
transform -1 0 3008 0 1 2370
box -8 -3 34 105
use FILL  FILL_5750
timestamp 1677677812
transform 1 0 3008 0 1 2370
box -8 -3 16 105
use FILL  FILL_5752
timestamp 1677677812
transform 1 0 3016 0 1 2370
box -8 -3 16 105
use FILL  FILL_5754
timestamp 1677677812
transform 1 0 3024 0 1 2370
box -8 -3 16 105
use FILL  FILL_5756
timestamp 1677677812
transform 1 0 3032 0 1 2370
box -8 -3 16 105
use FILL  FILL_5758
timestamp 1677677812
transform 1 0 3040 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_218
timestamp 1677677812
transform 1 0 3048 0 1 2370
box -8 -3 46 105
use FILL  FILL_5760
timestamp 1677677812
transform 1 0 3088 0 1 2370
box -8 -3 16 105
use FILL  FILL_5761
timestamp 1677677812
transform 1 0 3096 0 1 2370
box -8 -3 16 105
use FILL  FILL_5762
timestamp 1677677812
transform 1 0 3104 0 1 2370
box -8 -3 16 105
use FILL  FILL_5763
timestamp 1677677812
transform 1 0 3112 0 1 2370
box -8 -3 16 105
use FILL  FILL_5764
timestamp 1677677812
transform 1 0 3120 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_377
timestamp 1677677812
transform -1 0 3144 0 1 2370
box -9 -3 26 105
use FILL  FILL_5765
timestamp 1677677812
transform 1 0 3144 0 1 2370
box -8 -3 16 105
use FILL  FILL_5767
timestamp 1677677812
transform 1 0 3152 0 1 2370
box -8 -3 16 105
use FILL  FILL_5769
timestamp 1677677812
transform 1 0 3160 0 1 2370
box -8 -3 16 105
use FILL  FILL_5771
timestamp 1677677812
transform 1 0 3168 0 1 2370
box -8 -3 16 105
use FILL  FILL_5772
timestamp 1677677812
transform 1 0 3176 0 1 2370
box -8 -3 16 105
use FILL  FILL_5773
timestamp 1677677812
transform 1 0 3184 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_53
timestamp 1677677812
transform 1 0 3192 0 1 2370
box -5 -3 28 105
use FILL  FILL_5775
timestamp 1677677812
transform 1 0 3216 0 1 2370
box -8 -3 16 105
use FILL  FILL_5776
timestamp 1677677812
transform 1 0 3224 0 1 2370
box -8 -3 16 105
use FILL  FILL_5779
timestamp 1677677812
transform 1 0 3232 0 1 2370
box -8 -3 16 105
use FILL  FILL_5781
timestamp 1677677812
transform 1 0 3240 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_55
timestamp 1677677812
transform 1 0 3248 0 1 2370
box -5 -3 28 105
use BUFX2  BUFX2_56
timestamp 1677677812
transform 1 0 3272 0 1 2370
box -5 -3 28 105
use FILL  FILL_5783
timestamp 1677677812
transform 1 0 3296 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_34
timestamp 1677677812
transform -1 0 3336 0 1 2370
box -8 -3 40 105
use FILL  FILL_5784
timestamp 1677677812
transform 1 0 3336 0 1 2370
box -8 -3 16 105
use FILL  FILL_5797
timestamp 1677677812
transform 1 0 3344 0 1 2370
box -8 -3 16 105
use FILL  FILL_5799
timestamp 1677677812
transform 1 0 3352 0 1 2370
box -8 -3 16 105
use FILL  FILL_5801
timestamp 1677677812
transform 1 0 3360 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_35
timestamp 1677677812
transform -1 0 3400 0 1 2370
box -8 -3 40 105
use FILL  FILL_5802
timestamp 1677677812
transform 1 0 3400 0 1 2370
box -8 -3 16 105
use FILL  FILL_5803
timestamp 1677677812
transform 1 0 3408 0 1 2370
box -8 -3 16 105
use FILL  FILL_5804
timestamp 1677677812
transform 1 0 3416 0 1 2370
box -8 -3 16 105
use FILL  FILL_5805
timestamp 1677677812
transform 1 0 3424 0 1 2370
box -8 -3 16 105
use FILL  FILL_5810
timestamp 1677677812
transform 1 0 3432 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_234
timestamp 1677677812
transform 1 0 3440 0 1 2370
box -8 -3 46 105
use FILL  FILL_5812
timestamp 1677677812
transform 1 0 3480 0 1 2370
box -8 -3 16 105
use FILL  FILL_5813
timestamp 1677677812
transform 1 0 3488 0 1 2370
box -8 -3 16 105
use FILL  FILL_5814
timestamp 1677677812
transform 1 0 3496 0 1 2370
box -8 -3 16 105
use FILL  FILL_5815
timestamp 1677677812
transform 1 0 3504 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_331
timestamp 1677677812
transform 1 0 3512 0 1 2370
box -8 -3 104 105
use FILL  FILL_5820
timestamp 1677677812
transform 1 0 3608 0 1 2370
box -8 -3 16 105
use FILL  FILL_5821
timestamp 1677677812
transform 1 0 3616 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_220
timestamp 1677677812
transform 1 0 3624 0 1 2370
box -8 -3 46 105
use FILL  FILL_5822
timestamp 1677677812
transform 1 0 3664 0 1 2370
box -8 -3 16 105
use FILL  FILL_5823
timestamp 1677677812
transform 1 0 3672 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_332
timestamp 1677677812
transform 1 0 3680 0 1 2370
box -8 -3 104 105
use FILL  FILL_5824
timestamp 1677677812
transform 1 0 3776 0 1 2370
box -8 -3 16 105
use FILL  FILL_5825
timestamp 1677677812
transform 1 0 3784 0 1 2370
box -8 -3 16 105
use FILL  FILL_5826
timestamp 1677677812
transform 1 0 3792 0 1 2370
box -8 -3 16 105
use FILL  FILL_5827
timestamp 1677677812
transform 1 0 3800 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_379
timestamp 1677677812
transform 1 0 3808 0 1 2370
box -9 -3 26 105
use FILL  FILL_5828
timestamp 1677677812
transform 1 0 3824 0 1 2370
box -8 -3 16 105
use FILL  FILL_5838
timestamp 1677677812
transform 1 0 3832 0 1 2370
box -8 -3 16 105
use FILL  FILL_5839
timestamp 1677677812
transform 1 0 3840 0 1 2370
box -8 -3 16 105
use FILL  FILL_5840
timestamp 1677677812
transform 1 0 3848 0 1 2370
box -8 -3 16 105
use BUFX2  BUFX2_57
timestamp 1677677812
transform 1 0 3856 0 1 2370
box -5 -3 28 105
use FILL  FILL_5841
timestamp 1677677812
transform 1 0 3880 0 1 2370
box -8 -3 16 105
use FILL  FILL_5842
timestamp 1677677812
transform 1 0 3888 0 1 2370
box -8 -3 16 105
use FILL  FILL_5843
timestamp 1677677812
transform 1 0 3896 0 1 2370
box -8 -3 16 105
use FILL  FILL_5844
timestamp 1677677812
transform 1 0 3904 0 1 2370
box -8 -3 16 105
use FILL  FILL_5845
timestamp 1677677812
transform 1 0 3912 0 1 2370
box -8 -3 16 105
use FILL  FILL_5846
timestamp 1677677812
transform 1 0 3920 0 1 2370
box -8 -3 16 105
use FILL  FILL_5847
timestamp 1677677812
transform 1 0 3928 0 1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_222
timestamp 1677677812
transform 1 0 3936 0 1 2370
box -8 -3 46 105
use FILL  FILL_5849
timestamp 1677677812
transform 1 0 3976 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_336
timestamp 1677677812
transform -1 0 4080 0 1 2370
box -8 -3 104 105
use INVX2  INVX2_381
timestamp 1677677812
transform 1 0 4080 0 1 2370
box -9 -3 26 105
use FILL  FILL_5850
timestamp 1677677812
transform 1 0 4096 0 1 2370
box -8 -3 16 105
use FILL  FILL_5851
timestamp 1677677812
transform 1 0 4104 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_382
timestamp 1677677812
transform -1 0 4128 0 1 2370
box -9 -3 26 105
use FILL  FILL_5852
timestamp 1677677812
transform 1 0 4128 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_337
timestamp 1677677812
transform -1 0 4232 0 1 2370
box -8 -3 104 105
use OAI22X1  OAI22X1_223
timestamp 1677677812
transform 1 0 4232 0 1 2370
box -8 -3 46 105
use FILL  FILL_5853
timestamp 1677677812
transform 1 0 4272 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_383
timestamp 1677677812
transform 1 0 4280 0 1 2370
box -9 -3 26 105
use FILL  FILL_5854
timestamp 1677677812
transform 1 0 4296 0 1 2370
box -8 -3 16 105
use FILL  FILL_5855
timestamp 1677677812
transform 1 0 4304 0 1 2370
box -8 -3 16 105
use FILL  FILL_5856
timestamp 1677677812
transform 1 0 4312 0 1 2370
box -8 -3 16 105
use FILL  FILL_5857
timestamp 1677677812
transform 1 0 4320 0 1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_36
timestamp 1677677812
transform -1 0 4360 0 1 2370
box -8 -3 40 105
use FILL  FILL_5858
timestamp 1677677812
transform 1 0 4360 0 1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_340
timestamp 1677677812
transform 1 0 4368 0 1 2370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_341
timestamp 1677677812
transform 1 0 4464 0 1 2370
box -8 -3 104 105
use FILL  FILL_5875
timestamp 1677677812
transform 1 0 4560 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_384
timestamp 1677677812
transform 1 0 4568 0 1 2370
box -9 -3 26 105
use FILL  FILL_5876
timestamp 1677677812
transform 1 0 4584 0 1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_237
timestamp 1677677812
transform 1 0 4592 0 1 2370
box -8 -3 46 105
use FILL  FILL_5881
timestamp 1677677812
transform 1 0 4632 0 1 2370
box -8 -3 16 105
use FILL  FILL_5883
timestamp 1677677812
transform 1 0 4640 0 1 2370
box -8 -3 16 105
use FILL  FILL_5885
timestamp 1677677812
transform 1 0 4648 0 1 2370
box -8 -3 16 105
use FILL  FILL_5887
timestamp 1677677812
transform 1 0 4656 0 1 2370
box -8 -3 16 105
use INVX2  INVX2_386
timestamp 1677677812
transform -1 0 4680 0 1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_343
timestamp 1677677812
transform 1 0 4680 0 1 2370
box -8 -3 104 105
use FILL  FILL_5888
timestamp 1677677812
transform 1 0 4776 0 1 2370
box -8 -3 16 105
use FILL  FILL_5891
timestamp 1677677812
transform 1 0 4784 0 1 2370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_47
timestamp 1677677812
transform 1 0 4819 0 1 2370
box -10 -3 10 3
use M2_M1  M2_M1_4950
timestamp 1677677812
transform 1 0 84 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5038
timestamp 1677677812
transform 1 0 124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5039
timestamp 1677677812
transform 1 0 164 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5040
timestamp 1677677812
transform 1 0 172 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4542
timestamp 1677677812
transform 1 0 164 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4951
timestamp 1677677812
transform 1 0 188 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4952
timestamp 1677677812
transform 1 0 196 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4953
timestamp 1677677812
transform 1 0 212 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4438
timestamp 1677677812
transform 1 0 236 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4954
timestamp 1677677812
transform 1 0 236 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4507
timestamp 1677677812
transform 1 0 260 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5041
timestamp 1677677812
transform 1 0 180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5042
timestamp 1677677812
transform 1 0 188 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5043
timestamp 1677677812
transform 1 0 204 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5044
timestamp 1677677812
transform 1 0 228 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5045
timestamp 1677677812
transform 1 0 244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5046
timestamp 1677677812
transform 1 0 260 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4543
timestamp 1677677812
transform 1 0 196 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4569
timestamp 1677677812
transform 1 0 212 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4570
timestamp 1677677812
transform 1 0 260 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_4955
timestamp 1677677812
transform 1 0 300 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4482
timestamp 1677677812
transform 1 0 332 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4439
timestamp 1677677812
transform 1 0 364 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4956
timestamp 1677677812
transform 1 0 332 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4957
timestamp 1677677812
transform 1 0 348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5047
timestamp 1677677812
transform 1 0 324 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5048
timestamp 1677677812
transform 1 0 340 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4508
timestamp 1677677812
transform 1 0 356 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4958
timestamp 1677677812
transform 1 0 364 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4544
timestamp 1677677812
transform 1 0 348 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5049
timestamp 1677677812
transform 1 0 364 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4440
timestamp 1677677812
transform 1 0 396 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_4959
timestamp 1677677812
transform 1 0 380 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4960
timestamp 1677677812
transform 1 0 396 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4961
timestamp 1677677812
transform 1 0 404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5050
timestamp 1677677812
transform 1 0 388 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4514
timestamp 1677677812
transform 1 0 396 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4509
timestamp 1677677812
transform 1 0 412 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5051
timestamp 1677677812
transform 1 0 412 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4962
timestamp 1677677812
transform 1 0 460 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4963
timestamp 1677677812
transform 1 0 548 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5052
timestamp 1677677812
transform 1 0 444 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5053
timestamp 1677677812
transform 1 0 484 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4515
timestamp 1677677812
transform 1 0 532 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5054
timestamp 1677677812
transform 1 0 540 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4545
timestamp 1677677812
transform 1 0 444 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4546
timestamp 1677677812
transform 1 0 484 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4571
timestamp 1677677812
transform 1 0 508 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4572
timestamp 1677677812
transform 1 0 564 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5055
timestamp 1677677812
transform 1 0 580 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4441
timestamp 1677677812
transform 1 0 612 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4442
timestamp 1677677812
transform 1 0 636 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4483
timestamp 1677677812
transform 1 0 628 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4947
timestamp 1677677812
transform 1 0 636 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_5056
timestamp 1677677812
transform 1 0 636 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4547
timestamp 1677677812
transform 1 0 636 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4454
timestamp 1677677812
transform 1 0 660 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4484
timestamp 1677677812
transform 1 0 676 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4964
timestamp 1677677812
transform 1 0 668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5057
timestamp 1677677812
transform 1 0 676 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4573
timestamp 1677677812
transform 1 0 676 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_4965
timestamp 1677677812
transform 1 0 692 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5058
timestamp 1677677812
transform 1 0 716 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5059
timestamp 1677677812
transform 1 0 788 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4596
timestamp 1677677812
transform 1 0 796 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4597
timestamp 1677677812
transform 1 0 820 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4455
timestamp 1677677812
transform 1 0 852 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4485
timestamp 1677677812
transform 1 0 852 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4966
timestamp 1677677812
transform 1 0 852 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5060
timestamp 1677677812
transform 1 0 836 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4967
timestamp 1677677812
transform 1 0 876 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5061
timestamp 1677677812
transform 1 0 868 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5137
timestamp 1677677812
transform 1 0 908 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4598
timestamp 1677677812
transform 1 0 900 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4456
timestamp 1677677812
transform 1 0 940 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4510
timestamp 1677677812
transform 1 0 932 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4968
timestamp 1677677812
transform 1 0 940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5062
timestamp 1677677812
transform 1 0 932 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4548
timestamp 1677677812
transform 1 0 932 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4969
timestamp 1677677812
transform 1 0 956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5138
timestamp 1677677812
transform 1 0 956 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4457
timestamp 1677677812
transform 1 0 980 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4970
timestamp 1677677812
transform 1 0 988 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4549
timestamp 1677677812
transform 1 0 1012 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4592
timestamp 1677677812
transform 1 0 1004 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4443
timestamp 1677677812
transform 1 0 1124 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4458
timestamp 1677677812
transform 1 0 1084 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4486
timestamp 1677677812
transform 1 0 1044 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4487
timestamp 1677677812
transform 1 0 1060 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4971
timestamp 1677677812
transform 1 0 1044 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4459
timestamp 1677677812
transform 1 0 1140 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4460
timestamp 1677677812
transform 1 0 1156 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4488
timestamp 1677677812
transform 1 0 1132 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4489
timestamp 1677677812
transform 1 0 1172 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4972
timestamp 1677677812
transform 1 0 1140 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4973
timestamp 1677677812
transform 1 0 1148 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4974
timestamp 1677677812
transform 1 0 1164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4975
timestamp 1677677812
transform 1 0 1172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5063
timestamp 1677677812
transform 1 0 1084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5064
timestamp 1677677812
transform 1 0 1124 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5065
timestamp 1677677812
transform 1 0 1132 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4550
timestamp 1677677812
transform 1 0 1084 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4574
timestamp 1677677812
transform 1 0 1132 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5066
timestamp 1677677812
transform 1 0 1156 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5067
timestamp 1677677812
transform 1 0 1180 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4551
timestamp 1677677812
transform 1 0 1180 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4516
timestamp 1677677812
transform 1 0 1196 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4461
timestamp 1677677812
transform 1 0 1212 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4976
timestamp 1677677812
transform 1 0 1228 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4517
timestamp 1677677812
transform 1 0 1228 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_4977
timestamp 1677677812
transform 1 0 1236 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5139
timestamp 1677677812
transform 1 0 1284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5068
timestamp 1677677812
transform 1 0 1324 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4462
timestamp 1677677812
transform 1 0 1364 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4978
timestamp 1677677812
transform 1 0 1364 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4444
timestamp 1677677812
transform 1 0 1388 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4490
timestamp 1677677812
transform 1 0 1436 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4979
timestamp 1677677812
transform 1 0 1388 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4518
timestamp 1677677812
transform 1 0 1388 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5069
timestamp 1677677812
transform 1 0 1436 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4519
timestamp 1677677812
transform 1 0 1452 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5070
timestamp 1677677812
transform 1 0 1492 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4445
timestamp 1677677812
transform 1 0 1524 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4491
timestamp 1677677812
transform 1 0 1548 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4980
timestamp 1677677812
transform 1 0 1532 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4981
timestamp 1677677812
transform 1 0 1548 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4599
timestamp 1677677812
transform 1 0 1524 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5071
timestamp 1677677812
transform 1 0 1540 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5072
timestamp 1677677812
transform 1 0 1556 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4575
timestamp 1677677812
transform 1 0 1548 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4600
timestamp 1677677812
transform 1 0 1548 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4982
timestamp 1677677812
transform 1 0 1580 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5073
timestamp 1677677812
transform 1 0 1604 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4463
timestamp 1677677812
transform 1 0 1676 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4983
timestamp 1677677812
transform 1 0 1652 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4984
timestamp 1677677812
transform 1 0 1668 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4985
timestamp 1677677812
transform 1 0 1684 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5074
timestamp 1677677812
transform 1 0 1676 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4552
timestamp 1677677812
transform 1 0 1652 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4464
timestamp 1677677812
transform 1 0 1740 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4446
timestamp 1677677812
transform 1 0 1828 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4492
timestamp 1677677812
transform 1 0 1748 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4986
timestamp 1677677812
transform 1 0 1748 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5075
timestamp 1677677812
transform 1 0 1788 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4520
timestamp 1677677812
transform 1 0 1820 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5076
timestamp 1677677812
transform 1 0 1828 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5077
timestamp 1677677812
transform 1 0 1836 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4576
timestamp 1677677812
transform 1 0 1788 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4577
timestamp 1677677812
transform 1 0 1836 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4465
timestamp 1677677812
transform 1 0 1876 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4447
timestamp 1677677812
transform 1 0 1916 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4466
timestamp 1677677812
transform 1 0 1908 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4521
timestamp 1677677812
transform 1 0 1916 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4448
timestamp 1677677812
transform 1 0 1932 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4467
timestamp 1677677812
transform 1 0 1964 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4468
timestamp 1677677812
transform 1 0 2020 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4493
timestamp 1677677812
transform 1 0 1980 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_4987
timestamp 1677677812
transform 1 0 1932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4988
timestamp 1677677812
transform 1 0 1940 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4989
timestamp 1677677812
transform 1 0 1956 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4990
timestamp 1677677812
transform 1 0 1964 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4991
timestamp 1677677812
transform 1 0 1980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5078
timestamp 1677677812
transform 1 0 1932 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4522
timestamp 1677677812
transform 1 0 1940 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5079
timestamp 1677677812
transform 1 0 1948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5080
timestamp 1677677812
transform 1 0 2028 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4523
timestamp 1677677812
transform 1 0 2052 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5081
timestamp 1677677812
transform 1 0 2060 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5082
timestamp 1677677812
transform 1 0 2068 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4578
timestamp 1677677812
transform 1 0 2028 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4579
timestamp 1677677812
transform 1 0 2068 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_4992
timestamp 1677677812
transform 1 0 2164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4993
timestamp 1677677812
transform 1 0 2172 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5083
timestamp 1677677812
transform 1 0 2164 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4524
timestamp 1677677812
transform 1 0 2172 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5084
timestamp 1677677812
transform 1 0 2180 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5085
timestamp 1677677812
transform 1 0 2196 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4994
timestamp 1677677812
transform 1 0 2212 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5086
timestamp 1677677812
transform 1 0 2220 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4995
timestamp 1677677812
transform 1 0 2244 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4601
timestamp 1677677812
transform 1 0 2252 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5140
timestamp 1677677812
transform 1 0 2268 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4449
timestamp 1677677812
transform 1 0 2284 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4469
timestamp 1677677812
transform 1 0 2292 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4996
timestamp 1677677812
transform 1 0 2292 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_4997
timestamp 1677677812
transform 1 0 2308 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4494
timestamp 1677677812
transform 1 0 2332 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5087
timestamp 1677677812
transform 1 0 2332 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4602
timestamp 1677677812
transform 1 0 2332 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_4998
timestamp 1677677812
transform 1 0 2348 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5088
timestamp 1677677812
transform 1 0 2356 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4470
timestamp 1677677812
transform 1 0 2396 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_4999
timestamp 1677677812
transform 1 0 2404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5089
timestamp 1677677812
transform 1 0 2388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5090
timestamp 1677677812
transform 1 0 2396 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4471
timestamp 1677677812
transform 1 0 2420 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4472
timestamp 1677677812
transform 1 0 2516 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5000
timestamp 1677677812
transform 1 0 2516 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5091
timestamp 1677677812
transform 1 0 2476 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4495
timestamp 1677677812
transform 1 0 2532 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5092
timestamp 1677677812
transform 1 0 2580 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4525
timestamp 1677677812
transform 1 0 2652 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5093
timestamp 1677677812
transform 1 0 2684 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4580
timestamp 1677677812
transform 1 0 2684 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4496
timestamp 1677677812
transform 1 0 2700 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5001
timestamp 1677677812
transform 1 0 2700 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4526
timestamp 1677677812
transform 1 0 2700 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5094
timestamp 1677677812
transform 1 0 2724 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4581
timestamp 1677677812
transform 1 0 2724 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4450
timestamp 1677677812
transform 1 0 2788 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5095
timestamp 1677677812
transform 1 0 2788 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5096
timestamp 1677677812
transform 1 0 2844 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_4948
timestamp 1677677812
transform 1 0 2868 0 1 2345
box -2 -2 2 2
use M3_M2  M3_M2_4527
timestamp 1677677812
transform 1 0 2892 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5141
timestamp 1677677812
transform 1 0 2892 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5002
timestamp 1677677812
transform 1 0 2908 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5003
timestamp 1677677812
transform 1 0 2932 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5097
timestamp 1677677812
transform 1 0 2924 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4528
timestamp 1677677812
transform 1 0 2932 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5142
timestamp 1677677812
transform 1 0 2932 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_4949
timestamp 1677677812
transform 1 0 2964 0 1 2345
box -2 -2 2 2
use M2_M1  M2_M1_5143
timestamp 1677677812
transform 1 0 2956 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4582
timestamp 1677677812
transform 1 0 2948 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5098
timestamp 1677677812
transform 1 0 2996 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4583
timestamp 1677677812
transform 1 0 2996 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5004
timestamp 1677677812
transform 1 0 3020 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4584
timestamp 1677677812
transform 1 0 3036 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5005
timestamp 1677677812
transform 1 0 3060 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4529
timestamp 1677677812
transform 1 0 3060 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5099
timestamp 1677677812
transform 1 0 3092 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4530
timestamp 1677677812
transform 1 0 3108 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4603
timestamp 1677677812
transform 1 0 3068 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4604
timestamp 1677677812
transform 1 0 3092 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4531
timestamp 1677677812
transform 1 0 3156 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4553
timestamp 1677677812
transform 1 0 3156 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4473
timestamp 1677677812
transform 1 0 3172 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4497
timestamp 1677677812
transform 1 0 3188 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5006
timestamp 1677677812
transform 1 0 3188 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4532
timestamp 1677677812
transform 1 0 3180 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5100
timestamp 1677677812
transform 1 0 3188 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4585
timestamp 1677677812
transform 1 0 3172 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4554
timestamp 1677677812
transform 1 0 3204 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_4945
timestamp 1677677812
transform 1 0 3228 0 1 2355
box -2 -2 2 2
use M3_M2  M3_M2_4498
timestamp 1677677812
transform 1 0 3220 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5101
timestamp 1677677812
transform 1 0 3244 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4555
timestamp 1677677812
transform 1 0 3244 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4451
timestamp 1677677812
transform 1 0 3268 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5102
timestamp 1677677812
transform 1 0 3284 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4511
timestamp 1677677812
transform 1 0 3324 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_4946
timestamp 1677677812
transform 1 0 3348 0 1 2355
box -2 -2 2 2
use M2_M1  M2_M1_5007
timestamp 1677677812
transform 1 0 3388 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5008
timestamp 1677677812
transform 1 0 3404 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5103
timestamp 1677677812
transform 1 0 3396 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4556
timestamp 1677677812
transform 1 0 3396 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4605
timestamp 1677677812
transform 1 0 3388 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5009
timestamp 1677677812
transform 1 0 3428 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4533
timestamp 1677677812
transform 1 0 3428 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4474
timestamp 1677677812
transform 1 0 3444 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5010
timestamp 1677677812
transform 1 0 3444 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4557
timestamp 1677677812
transform 1 0 3444 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4475
timestamp 1677677812
transform 1 0 3492 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4499
timestamp 1677677812
transform 1 0 3468 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4500
timestamp 1677677812
transform 1 0 3500 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5104
timestamp 1677677812
transform 1 0 3460 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5105
timestamp 1677677812
transform 1 0 3468 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5106
timestamp 1677677812
transform 1 0 3484 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5107
timestamp 1677677812
transform 1 0 3500 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4586
timestamp 1677677812
transform 1 0 3468 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4476
timestamp 1677677812
transform 1 0 3524 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5011
timestamp 1677677812
transform 1 0 3524 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4587
timestamp 1677677812
transform 1 0 3516 0 1 2305
box -3 -3 3 3
use M2_M1  M2_M1_5012
timestamp 1677677812
transform 1 0 3540 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5013
timestamp 1677677812
transform 1 0 3628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5108
timestamp 1677677812
transform 1 0 3572 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5109
timestamp 1677677812
transform 1 0 3620 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4588
timestamp 1677677812
transform 1 0 3532 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4589
timestamp 1677677812
transform 1 0 3572 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4606
timestamp 1677677812
transform 1 0 3580 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4534
timestamp 1677677812
transform 1 0 3628 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4477
timestamp 1677677812
transform 1 0 3668 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5014
timestamp 1677677812
transform 1 0 3660 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5015
timestamp 1677677812
transform 1 0 3676 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5110
timestamp 1677677812
transform 1 0 3644 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5111
timestamp 1677677812
transform 1 0 3668 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4558
timestamp 1677677812
transform 1 0 3660 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5016
timestamp 1677677812
transform 1 0 3716 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5112
timestamp 1677677812
transform 1 0 3740 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4559
timestamp 1677677812
transform 1 0 3740 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4452
timestamp 1677677812
transform 1 0 3820 0 1 2365
box -3 -3 3 3
use M3_M2  M3_M2_4478
timestamp 1677677812
transform 1 0 3812 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5113
timestamp 1677677812
transform 1 0 3812 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4590
timestamp 1677677812
transform 1 0 3828 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4453
timestamp 1677677812
transform 1 0 3844 0 1 2365
box -3 -3 3 3
use M2_M1  M2_M1_5017
timestamp 1677677812
transform 1 0 3844 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5114
timestamp 1677677812
transform 1 0 3892 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5115
timestamp 1677677812
transform 1 0 3924 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4560
timestamp 1677677812
transform 1 0 3892 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5018
timestamp 1677677812
transform 1 0 3940 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4535
timestamp 1677677812
transform 1 0 3940 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5019
timestamp 1677677812
transform 1 0 3964 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5020
timestamp 1677677812
transform 1 0 3980 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5021
timestamp 1677677812
transform 1 0 3988 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5116
timestamp 1677677812
transform 1 0 3948 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5117
timestamp 1677677812
transform 1 0 3972 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4561
timestamp 1677677812
transform 1 0 3964 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4591
timestamp 1677677812
transform 1 0 3948 0 1 2305
box -3 -3 3 3
use M3_M2  M3_M2_4607
timestamp 1677677812
transform 1 0 3940 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4536
timestamp 1677677812
transform 1 0 3988 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4501
timestamp 1677677812
transform 1 0 4020 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5022
timestamp 1677677812
transform 1 0 4020 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5118
timestamp 1677677812
transform 1 0 4012 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5119
timestamp 1677677812
transform 1 0 4028 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4608
timestamp 1677677812
transform 1 0 4028 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5023
timestamp 1677677812
transform 1 0 4044 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5024
timestamp 1677677812
transform 1 0 4060 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4502
timestamp 1677677812
transform 1 0 4116 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5025
timestamp 1677677812
transform 1 0 4164 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5120
timestamp 1677677812
transform 1 0 4084 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5121
timestamp 1677677812
transform 1 0 4116 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4537
timestamp 1677677812
transform 1 0 4164 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4562
timestamp 1677677812
transform 1 0 4100 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4609
timestamp 1677677812
transform 1 0 4180 0 1 2285
box -3 -3 3 3
use M3_M2  M3_M2_4479
timestamp 1677677812
transform 1 0 4236 0 1 2355
box -3 -3 3 3
use M2_M1  M2_M1_5026
timestamp 1677677812
transform 1 0 4196 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4538
timestamp 1677677812
transform 1 0 4196 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4539
timestamp 1677677812
transform 1 0 4220 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5122
timestamp 1677677812
transform 1 0 4244 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5123
timestamp 1677677812
transform 1 0 4276 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4610
timestamp 1677677812
transform 1 0 4252 0 1 2285
box -3 -3 3 3
use M2_M1  M2_M1_5144
timestamp 1677677812
transform 1 0 4284 0 1 2315
box -2 -2 2 2
use M2_M1  M2_M1_5146
timestamp 1677677812
transform 1 0 4284 0 1 2305
box -2 -2 2 2
use M3_M2  M3_M2_4593
timestamp 1677677812
transform 1 0 4284 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5124
timestamp 1677677812
transform 1 0 4308 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4563
timestamp 1677677812
transform 1 0 4308 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5027
timestamp 1677677812
transform 1 0 4340 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5125
timestamp 1677677812
transform 1 0 4356 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5145
timestamp 1677677812
transform 1 0 4364 0 1 2315
box -2 -2 2 2
use M3_M2  M3_M2_4594
timestamp 1677677812
transform 1 0 4364 0 1 2295
box -3 -3 3 3
use M3_M2  M3_M2_4480
timestamp 1677677812
transform 1 0 4420 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4503
timestamp 1677677812
transform 1 0 4436 0 1 2345
box -3 -3 3 3
use M3_M2  M3_M2_4504
timestamp 1677677812
transform 1 0 4492 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5028
timestamp 1677677812
transform 1 0 4412 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5029
timestamp 1677677812
transform 1 0 4420 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5030
timestamp 1677677812
transform 1 0 4436 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5031
timestamp 1677677812
transform 1 0 4452 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5032
timestamp 1677677812
transform 1 0 4468 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5126
timestamp 1677677812
transform 1 0 4388 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5127
timestamp 1677677812
transform 1 0 4404 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5128
timestamp 1677677812
transform 1 0 4420 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5129
timestamp 1677677812
transform 1 0 4444 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4564
timestamp 1677677812
transform 1 0 4412 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4565
timestamp 1677677812
transform 1 0 4444 0 1 2315
box -3 -3 3 3
use M2_M1  M2_M1_5130
timestamp 1677677812
transform 1 0 4492 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4595
timestamp 1677677812
transform 1 0 4460 0 1 2295
box -3 -3 3 3
use M2_M1  M2_M1_5131
timestamp 1677677812
transform 1 0 4564 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5132
timestamp 1677677812
transform 1 0 4572 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4566
timestamp 1677677812
transform 1 0 4564 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4481
timestamp 1677677812
transform 1 0 4596 0 1 2355
box -3 -3 3 3
use M3_M2  M3_M2_4505
timestamp 1677677812
transform 1 0 4612 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5033
timestamp 1677677812
transform 1 0 4596 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5034
timestamp 1677677812
transform 1 0 4612 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4512
timestamp 1677677812
transform 1 0 4620 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5035
timestamp 1677677812
transform 1 0 4628 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5036
timestamp 1677677812
transform 1 0 4636 0 1 2335
box -2 -2 2 2
use M2_M1  M2_M1_5133
timestamp 1677677812
transform 1 0 4604 0 1 2325
box -2 -2 2 2
use M2_M1  M2_M1_5134
timestamp 1677677812
transform 1 0 4620 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4567
timestamp 1677677812
transform 1 0 4604 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4540
timestamp 1677677812
transform 1 0 4644 0 1 2325
box -3 -3 3 3
use M3_M2  M3_M2_4568
timestamp 1677677812
transform 1 0 4636 0 1 2315
box -3 -3 3 3
use M3_M2  M3_M2_4506
timestamp 1677677812
transform 1 0 4692 0 1 2345
box -3 -3 3 3
use M2_M1  M2_M1_5037
timestamp 1677677812
transform 1 0 4668 0 1 2335
box -2 -2 2 2
use M3_M2  M3_M2_4541
timestamp 1677677812
transform 1 0 4668 0 1 2325
box -3 -3 3 3
use M2_M1  M2_M1_5135
timestamp 1677677812
transform 1 0 4692 0 1 2325
box -2 -2 2 2
use M3_M2  M3_M2_4513
timestamp 1677677812
transform 1 0 4764 0 1 2335
box -3 -3 3 3
use M2_M1  M2_M1_5136
timestamp 1677677812
transform 1 0 4764 0 1 2325
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_48
timestamp 1677677812
transform 1 0 24 0 1 2270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_315
timestamp 1677677812
transform 1 0 72 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_365
timestamp 1677677812
transform -1 0 184 0 -1 2370
box -9 -3 26 105
use AOI22X1  AOI22X1_223
timestamp 1677677812
transform -1 0 224 0 -1 2370
box -8 -3 46 105
use AOI22X1  AOI22X1_224
timestamp 1677677812
transform 1 0 224 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5400
timestamp 1677677812
transform 1 0 264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5402
timestamp 1677677812
transform 1 0 272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5404
timestamp 1677677812
transform 1 0 280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5417
timestamp 1677677812
transform 1 0 288 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5418
timestamp 1677677812
transform 1 0 296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5419
timestamp 1677677812
transform 1 0 304 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_211
timestamp 1677677812
transform 1 0 312 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5420
timestamp 1677677812
transform 1 0 352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5421
timestamp 1677677812
transform 1 0 360 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_226
timestamp 1677677812
transform 1 0 368 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5422
timestamp 1677677812
transform 1 0 408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5423
timestamp 1677677812
transform 1 0 416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5424
timestamp 1677677812
transform 1 0 424 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_367
timestamp 1677677812
transform 1 0 432 0 -1 2370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_317
timestamp 1677677812
transform 1 0 448 0 -1 2370
box -8 -3 104 105
use BUFX2  BUFX2_49
timestamp 1677677812
transform -1 0 568 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5425
timestamp 1677677812
transform 1 0 568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5427
timestamp 1677677812
transform 1 0 576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5429
timestamp 1677677812
transform 1 0 584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5434
timestamp 1677677812
transform 1 0 592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5435
timestamp 1677677812
transform 1 0 600 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_50
timestamp 1677677812
transform -1 0 632 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5436
timestamp 1677677812
transform 1 0 632 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_55
timestamp 1677677812
transform 1 0 640 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5437
timestamp 1677677812
transform 1 0 664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5438
timestamp 1677677812
transform 1 0 672 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_319
timestamp 1677677812
transform 1 0 680 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5439
timestamp 1677677812
transform 1 0 776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5441
timestamp 1677677812
transform 1 0 784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5443
timestamp 1677677812
transform 1 0 792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5445
timestamp 1677677812
transform 1 0 800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5449
timestamp 1677677812
transform 1 0 808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5450
timestamp 1677677812
transform 1 0 816 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_109
timestamp 1677677812
transform 1 0 824 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5451
timestamp 1677677812
transform 1 0 856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5453
timestamp 1677677812
transform 1 0 864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5455
timestamp 1677677812
transform 1 0 872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5457
timestamp 1677677812
transform 1 0 880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5459
timestamp 1677677812
transform 1 0 888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5461
timestamp 1677677812
transform 1 0 896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5463
timestamp 1677677812
transform 1 0 904 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_227
timestamp 1677677812
transform 1 0 912 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5470
timestamp 1677677812
transform 1 0 952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5472
timestamp 1677677812
transform 1 0 960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5474
timestamp 1677677812
transform 1 0 968 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5476
timestamp 1677677812
transform 1 0 976 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5478
timestamp 1677677812
transform 1 0 984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5480
timestamp 1677677812
transform 1 0 992 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5482
timestamp 1677677812
transform 1 0 1000 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5484
timestamp 1677677812
transform 1 0 1008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5486
timestamp 1677677812
transform 1 0 1016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5488
timestamp 1677677812
transform 1 0 1024 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_320
timestamp 1677677812
transform 1 0 1032 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5502
timestamp 1677677812
transform 1 0 1128 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_228
timestamp 1677677812
transform 1 0 1136 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5506
timestamp 1677677812
transform 1 0 1176 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5507
timestamp 1677677812
transform 1 0 1184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5508
timestamp 1677677812
transform 1 0 1192 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5509
timestamp 1677677812
transform 1 0 1200 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_369
timestamp 1677677812
transform -1 0 1224 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5510
timestamp 1677677812
transform 1 0 1224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5511
timestamp 1677677812
transform 1 0 1232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5512
timestamp 1677677812
transform 1 0 1240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5513
timestamp 1677677812
transform 1 0 1248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5514
timestamp 1677677812
transform 1 0 1256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5515
timestamp 1677677812
transform 1 0 1264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5517
timestamp 1677677812
transform 1 0 1272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5519
timestamp 1677677812
transform 1 0 1280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5521
timestamp 1677677812
transform 1 0 1288 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_111
timestamp 1677677812
transform -1 0 1328 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5523
timestamp 1677677812
transform 1 0 1328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5525
timestamp 1677677812
transform 1 0 1336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5527
timestamp 1677677812
transform 1 0 1344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5529
timestamp 1677677812
transform 1 0 1352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5531
timestamp 1677677812
transform 1 0 1360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5533
timestamp 1677677812
transform 1 0 1368 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_322
timestamp 1677677812
transform 1 0 1376 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5542
timestamp 1677677812
transform 1 0 1472 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5543
timestamp 1677677812
transform 1 0 1480 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5545
timestamp 1677677812
transform 1 0 1488 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5547
timestamp 1677677812
transform 1 0 1496 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5549
timestamp 1677677812
transform 1 0 1504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5551
timestamp 1677677812
transform 1 0 1512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5553
timestamp 1677677812
transform 1 0 1520 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_214
timestamp 1677677812
transform -1 0 1568 0 -1 2370
box -8 -3 46 105
use M3_M2  M3_M2_4611
timestamp 1677677812
transform 1 0 1580 0 1 2275
box -3 -3 3 3
use FILL  FILL_5555
timestamp 1677677812
transform 1 0 1568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5557
timestamp 1677677812
transform 1 0 1576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5559
timestamp 1677677812
transform 1 0 1584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5561
timestamp 1677677812
transform 1 0 1592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5563
timestamp 1677677812
transform 1 0 1600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5565
timestamp 1677677812
transform 1 0 1608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5567
timestamp 1677677812
transform 1 0 1616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5568
timestamp 1677677812
transform 1 0 1624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5569
timestamp 1677677812
transform 1 0 1632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5570
timestamp 1677677812
transform 1 0 1640 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_215
timestamp 1677677812
transform 1 0 1648 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5571
timestamp 1677677812
transform 1 0 1688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5572
timestamp 1677677812
transform 1 0 1696 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5573
timestamp 1677677812
transform 1 0 1704 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5574
timestamp 1677677812
transform 1 0 1712 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5576
timestamp 1677677812
transform 1 0 1720 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5586
timestamp 1677677812
transform 1 0 1728 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_324
timestamp 1677677812
transform 1 0 1736 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5587
timestamp 1677677812
transform 1 0 1832 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5589
timestamp 1677677812
transform 1 0 1840 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5591
timestamp 1677677812
transform 1 0 1848 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5593
timestamp 1677677812
transform 1 0 1856 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5615
timestamp 1677677812
transform 1 0 1864 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_372
timestamp 1677677812
transform -1 0 1888 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5616
timestamp 1677677812
transform 1 0 1888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5617
timestamp 1677677812
transform 1 0 1896 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5618
timestamp 1677677812
transform 1 0 1904 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5619
timestamp 1677677812
transform 1 0 1912 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5620
timestamp 1677677812
transform 1 0 1920 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_229
timestamp 1677677812
transform -1 0 1968 0 -1 2370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_325
timestamp 1677677812
transform 1 0 1968 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5621
timestamp 1677677812
transform 1 0 2064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5622
timestamp 1677677812
transform 1 0 2072 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5623
timestamp 1677677812
transform 1 0 2080 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_373
timestamp 1677677812
transform -1 0 2104 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5624
timestamp 1677677812
transform 1 0 2104 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5626
timestamp 1677677812
transform 1 0 2112 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5628
timestamp 1677677812
transform 1 0 2120 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4612
timestamp 1677677812
transform 1 0 2140 0 1 2275
box -3 -3 3 3
use FILL  FILL_5630
timestamp 1677677812
transform 1 0 2128 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5632
timestamp 1677677812
transform 1 0 2136 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5634
timestamp 1677677812
transform 1 0 2144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5642
timestamp 1677677812
transform 1 0 2152 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_230
timestamp 1677677812
transform -1 0 2200 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5643
timestamp 1677677812
transform 1 0 2200 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5645
timestamp 1677677812
transform 1 0 2208 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5647
timestamp 1677677812
transform 1 0 2216 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5649
timestamp 1677677812
transform 1 0 2224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5651
timestamp 1677677812
transform 1 0 2232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5653
timestamp 1677677812
transform 1 0 2240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5655
timestamp 1677677812
transform 1 0 2248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5657
timestamp 1677677812
transform 1 0 2256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5658
timestamp 1677677812
transform 1 0 2264 0 -1 2370
box -8 -3 16 105
use BUFX2  BUFX2_52
timestamp 1677677812
transform 1 0 2272 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5659
timestamp 1677677812
transform 1 0 2296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5661
timestamp 1677677812
transform 1 0 2304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5663
timestamp 1677677812
transform 1 0 2312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5665
timestamp 1677677812
transform 1 0 2320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5667
timestamp 1677677812
transform 1 0 2328 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_232
timestamp 1677677812
transform 1 0 2336 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5672
timestamp 1677677812
transform 1 0 2376 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5674
timestamp 1677677812
transform 1 0 2384 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5676
timestamp 1677677812
transform 1 0 2392 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5682
timestamp 1677677812
transform 1 0 2400 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5683
timestamp 1677677812
transform 1 0 2408 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5684
timestamp 1677677812
transform 1 0 2416 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5685
timestamp 1677677812
transform 1 0 2424 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_327
timestamp 1677677812
transform -1 0 2528 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5686
timestamp 1677677812
transform 1 0 2528 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5688
timestamp 1677677812
transform 1 0 2536 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5690
timestamp 1677677812
transform 1 0 2544 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5692
timestamp 1677677812
transform 1 0 2552 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5693
timestamp 1677677812
transform 1 0 2560 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5694
timestamp 1677677812
transform 1 0 2568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5695
timestamp 1677677812
transform 1 0 2576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5696
timestamp 1677677812
transform 1 0 2584 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5697
timestamp 1677677812
transform 1 0 2592 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5699
timestamp 1677677812
transform 1 0 2600 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5701
timestamp 1677677812
transform 1 0 2608 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5703
timestamp 1677677812
transform 1 0 2616 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5705
timestamp 1677677812
transform 1 0 2624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5707
timestamp 1677677812
transform 1 0 2632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5709
timestamp 1677677812
transform 1 0 2640 0 -1 2370
box -8 -3 16 105
use INVX2  INVX2_376
timestamp 1677677812
transform 1 0 2648 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5711
timestamp 1677677812
transform 1 0 2664 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5713
timestamp 1677677812
transform 1 0 2672 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5715
timestamp 1677677812
transform 1 0 2680 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_329
timestamp 1677677812
transform 1 0 2688 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5717
timestamp 1677677812
transform 1 0 2784 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5719
timestamp 1677677812
transform 1 0 2792 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5721
timestamp 1677677812
transform 1 0 2800 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5727
timestamp 1677677812
transform 1 0 2808 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5728
timestamp 1677677812
transform 1 0 2816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5729
timestamp 1677677812
transform 1 0 2824 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_113
timestamp 1677677812
transform 1 0 2832 0 -1 2370
box -8 -3 34 105
use FILL  FILL_5730
timestamp 1677677812
transform 1 0 2864 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5732
timestamp 1677677812
transform 1 0 2872 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5734
timestamp 1677677812
transform 1 0 2880 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5737
timestamp 1677677812
transform 1 0 2888 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5738
timestamp 1677677812
transform 1 0 2896 0 -1 2370
box -8 -3 16 105
use NOR2X1  NOR2X1_57
timestamp 1677677812
transform 1 0 2904 0 -1 2370
box -8 -3 32 105
use FILL  FILL_5739
timestamp 1677677812
transform 1 0 2928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5741
timestamp 1677677812
transform 1 0 2936 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5743
timestamp 1677677812
transform 1 0 2944 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5745
timestamp 1677677812
transform 1 0 2952 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5747
timestamp 1677677812
transform 1 0 2960 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5749
timestamp 1677677812
transform 1 0 2968 0 -1 2370
box -8 -3 16 105
use OAI21X1  OAI21X1_116
timestamp 1677677812
transform -1 0 3008 0 -1 2370
box -8 -3 34 105
use M3_M2  M3_M2_4613
timestamp 1677677812
transform 1 0 3020 0 1 2275
box -3 -3 3 3
use FILL  FILL_5751
timestamp 1677677812
transform 1 0 3008 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5753
timestamp 1677677812
transform 1 0 3016 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5755
timestamp 1677677812
transform 1 0 3024 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5757
timestamp 1677677812
transform 1 0 3032 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4614
timestamp 1677677812
transform 1 0 3076 0 1 2275
box -3 -3 3 3
use FILL  FILL_5759
timestamp 1677677812
transform 1 0 3040 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_330
timestamp 1677677812
transform 1 0 3048 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5766
timestamp 1677677812
transform 1 0 3144 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5768
timestamp 1677677812
transform 1 0 3152 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5770
timestamp 1677677812
transform 1 0 3160 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4615
timestamp 1677677812
transform 1 0 3188 0 1 2275
box -3 -3 3 3
use INVX2  INVX2_378
timestamp 1677677812
transform 1 0 3168 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5774
timestamp 1677677812
transform 1 0 3184 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5777
timestamp 1677677812
transform 1 0 3192 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4616
timestamp 1677677812
transform 1 0 3212 0 1 2275
box -3 -3 3 3
use BUFX2  BUFX2_54
timestamp 1677677812
transform -1 0 3224 0 -1 2370
box -5 -3 28 105
use FILL  FILL_5778
timestamp 1677677812
transform 1 0 3224 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5780
timestamp 1677677812
transform 1 0 3232 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5782
timestamp 1677677812
transform 1 0 3240 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5785
timestamp 1677677812
transform 1 0 3248 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5786
timestamp 1677677812
transform 1 0 3256 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5787
timestamp 1677677812
transform 1 0 3264 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5788
timestamp 1677677812
transform 1 0 3272 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5789
timestamp 1677677812
transform 1 0 3280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5790
timestamp 1677677812
transform 1 0 3288 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4617
timestamp 1677677812
transform 1 0 3308 0 1 2275
box -3 -3 3 3
use FILL  FILL_5791
timestamp 1677677812
transform 1 0 3296 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5792
timestamp 1677677812
transform 1 0 3304 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5793
timestamp 1677677812
transform 1 0 3312 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5794
timestamp 1677677812
transform 1 0 3320 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5795
timestamp 1677677812
transform 1 0 3328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5796
timestamp 1677677812
transform 1 0 3336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5798
timestamp 1677677812
transform 1 0 3344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5800
timestamp 1677677812
transform 1 0 3352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5806
timestamp 1677677812
transform 1 0 3360 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5807
timestamp 1677677812
transform 1 0 3368 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5808
timestamp 1677677812
transform 1 0 3376 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_219
timestamp 1677677812
transform -1 0 3424 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5809
timestamp 1677677812
transform 1 0 3424 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5811
timestamp 1677677812
transform 1 0 3432 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5816
timestamp 1677677812
transform 1 0 3440 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5817
timestamp 1677677812
transform 1 0 3448 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5818
timestamp 1677677812
transform 1 0 3456 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_235
timestamp 1677677812
transform -1 0 3504 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5819
timestamp 1677677812
transform 1 0 3504 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5829
timestamp 1677677812
transform 1 0 3512 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5830
timestamp 1677677812
transform 1 0 3520 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_333
timestamp 1677677812
transform 1 0 3528 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5831
timestamp 1677677812
transform 1 0 3624 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5832
timestamp 1677677812
transform 1 0 3632 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_221
timestamp 1677677812
transform 1 0 3640 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5833
timestamp 1677677812
transform 1 0 3680 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5834
timestamp 1677677812
transform 1 0 3688 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5835
timestamp 1677677812
transform 1 0 3696 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_334
timestamp 1677677812
transform 1 0 3704 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_380
timestamp 1677677812
transform 1 0 3800 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5836
timestamp 1677677812
transform 1 0 3816 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5837
timestamp 1677677812
transform 1 0 3824 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4618
timestamp 1677677812
transform 1 0 3892 0 1 2275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_335
timestamp 1677677812
transform 1 0 3832 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5848
timestamp 1677677812
transform 1 0 3928 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5859
timestamp 1677677812
transform 1 0 3936 0 -1 2370
box -8 -3 16 105
use M3_M2  M3_M2_4619
timestamp 1677677812
transform 1 0 3980 0 1 2275
box -3 -3 3 3
use OAI22X1  OAI22X1_224
timestamp 1677677812
transform 1 0 3944 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5860
timestamp 1677677812
transform 1 0 3984 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5861
timestamp 1677677812
transform 1 0 3992 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_225
timestamp 1677677812
transform 1 0 4000 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5862
timestamp 1677677812
transform 1 0 4040 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5863
timestamp 1677677812
transform 1 0 4048 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5864
timestamp 1677677812
transform 1 0 4056 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5865
timestamp 1677677812
transform 1 0 4064 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5866
timestamp 1677677812
transform 1 0 4072 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_338
timestamp 1677677812
transform -1 0 4176 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5867
timestamp 1677677812
transform 1 0 4176 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_339
timestamp 1677677812
transform 1 0 4184 0 -1 2370
box -8 -3 104 105
use FILL  FILL_5868
timestamp 1677677812
transform 1 0 4280 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5869
timestamp 1677677812
transform 1 0 4288 0 -1 2370
box -8 -3 16 105
use NAND3X1  NAND3X1_37
timestamp 1677677812
transform 1 0 4296 0 -1 2370
box -8 -3 40 105
use FILL  FILL_5870
timestamp 1677677812
transform 1 0 4328 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5871
timestamp 1677677812
transform 1 0 4336 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5872
timestamp 1677677812
transform 1 0 4344 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5873
timestamp 1677677812
transform 1 0 4352 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5874
timestamp 1677677812
transform 1 0 4360 0 -1 2370
box -8 -3 16 105
use AOI22X1  AOI22X1_236
timestamp 1677677812
transform 1 0 4368 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5877
timestamp 1677677812
transform 1 0 4408 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_226
timestamp 1677677812
transform 1 0 4416 0 -1 2370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_342
timestamp 1677677812
transform 1 0 4456 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_385
timestamp 1677677812
transform 1 0 4552 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5878
timestamp 1677677812
transform 1 0 4568 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5879
timestamp 1677677812
transform 1 0 4576 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5880
timestamp 1677677812
transform 1 0 4584 0 -1 2370
box -8 -3 16 105
use OAI22X1  OAI22X1_227
timestamp 1677677812
transform 1 0 4592 0 -1 2370
box -8 -3 46 105
use FILL  FILL_5882
timestamp 1677677812
transform 1 0 4632 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5884
timestamp 1677677812
transform 1 0 4640 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5886
timestamp 1677677812
transform 1 0 4648 0 -1 2370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_344
timestamp 1677677812
transform 1 0 4656 0 -1 2370
box -8 -3 104 105
use INVX2  INVX2_387
timestamp 1677677812
transform 1 0 4752 0 -1 2370
box -9 -3 26 105
use FILL  FILL_5889
timestamp 1677677812
transform 1 0 4768 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5890
timestamp 1677677812
transform 1 0 4776 0 -1 2370
box -8 -3 16 105
use FILL  FILL_5892
timestamp 1677677812
transform 1 0 4784 0 -1 2370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_49
timestamp 1677677812
transform 1 0 4843 0 1 2270
box -10 -3 10 3
use M3_M2  M3_M2_4667
timestamp 1677677812
transform 1 0 132 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4655
timestamp 1677677812
transform 1 0 180 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4668
timestamp 1677677812
transform 1 0 172 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5161
timestamp 1677677812
transform 1 0 132 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5162
timestamp 1677677812
transform 1 0 164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5271
timestamp 1677677812
transform 1 0 84 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5272
timestamp 1677677812
transform 1 0 180 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4786
timestamp 1677677812
transform 1 0 188 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4669
timestamp 1677677812
transform 1 0 204 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5163
timestamp 1677677812
transform 1 0 204 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4627
timestamp 1677677812
transform 1 0 228 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4628
timestamp 1677677812
transform 1 0 252 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4633
timestamp 1677677812
transform 1 0 292 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4656
timestamp 1677677812
transform 1 0 244 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4670
timestamp 1677677812
transform 1 0 244 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5164
timestamp 1677677812
transform 1 0 244 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5165
timestamp 1677677812
transform 1 0 300 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5273
timestamp 1677677812
transform 1 0 220 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4751
timestamp 1677677812
transform 1 0 220 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4752
timestamp 1677677812
transform 1 0 292 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4787
timestamp 1677677812
transform 1 0 212 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5166
timestamp 1677677812
transform 1 0 324 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5167
timestamp 1677677812
transform 1 0 372 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4671
timestamp 1677677812
transform 1 0 420 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4707
timestamp 1677677812
transform 1 0 396 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5168
timestamp 1677677812
transform 1 0 404 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5169
timestamp 1677677812
transform 1 0 420 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5274
timestamp 1677677812
transform 1 0 388 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5275
timestamp 1677677812
transform 1 0 396 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5276
timestamp 1677677812
transform 1 0 412 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5277
timestamp 1677677812
transform 1 0 420 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4634
timestamp 1677677812
transform 1 0 460 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4657
timestamp 1677677812
transform 1 0 460 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4708
timestamp 1677677812
transform 1 0 452 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5278
timestamp 1677677812
transform 1 0 452 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4672
timestamp 1677677812
transform 1 0 492 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5170
timestamp 1677677812
transform 1 0 476 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4709
timestamp 1677677812
transform 1 0 484 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5171
timestamp 1677677812
transform 1 0 492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5279
timestamp 1677677812
transform 1 0 484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5280
timestamp 1677677812
transform 1 0 492 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4658
timestamp 1677677812
transform 1 0 620 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4673
timestamp 1677677812
transform 1 0 556 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4674
timestamp 1677677812
transform 1 0 596 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5172
timestamp 1677677812
transform 1 0 556 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5173
timestamp 1677677812
transform 1 0 564 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4710
timestamp 1677677812
transform 1 0 572 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5174
timestamp 1677677812
transform 1 0 596 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4711
timestamp 1677677812
transform 1 0 644 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5281
timestamp 1677677812
transform 1 0 644 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4753
timestamp 1677677812
transform 1 0 620 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4754
timestamp 1677677812
transform 1 0 644 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4675
timestamp 1677677812
transform 1 0 692 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5282
timestamp 1677677812
transform 1 0 692 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4755
timestamp 1677677812
transform 1 0 692 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5175
timestamp 1677677812
transform 1 0 716 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4712
timestamp 1677677812
transform 1 0 756 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4676
timestamp 1677677812
transform 1 0 772 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4659
timestamp 1677677812
transform 1 0 804 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5176
timestamp 1677677812
transform 1 0 780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5177
timestamp 1677677812
transform 1 0 796 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5178
timestamp 1677677812
transform 1 0 812 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5283
timestamp 1677677812
transform 1 0 788 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5284
timestamp 1677677812
transform 1 0 812 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4756
timestamp 1677677812
transform 1 0 796 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4788
timestamp 1677677812
transform 1 0 780 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4660
timestamp 1677677812
transform 1 0 828 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5285
timestamp 1677677812
transform 1 0 836 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5179
timestamp 1677677812
transform 1 0 860 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4757
timestamp 1677677812
transform 1 0 860 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4789
timestamp 1677677812
transform 1 0 860 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4635
timestamp 1677677812
transform 1 0 892 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4661
timestamp 1677677812
transform 1 0 900 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4636
timestamp 1677677812
transform 1 0 924 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5180
timestamp 1677677812
transform 1 0 900 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5181
timestamp 1677677812
transform 1 0 916 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5286
timestamp 1677677812
transform 1 0 908 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4727
timestamp 1677677812
transform 1 0 916 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4713
timestamp 1677677812
transform 1 0 940 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5287
timestamp 1677677812
transform 1 0 940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5182
timestamp 1677677812
transform 1 0 980 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5183
timestamp 1677677812
transform 1 0 1004 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5184
timestamp 1677677812
transform 1 0 1020 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5185
timestamp 1677677812
transform 1 0 1028 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4758
timestamp 1677677812
transform 1 0 1028 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4677
timestamp 1677677812
transform 1 0 1044 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5288
timestamp 1677677812
transform 1 0 1052 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4790
timestamp 1677677812
transform 1 0 1044 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4728
timestamp 1677677812
transform 1 0 1068 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4759
timestamp 1677677812
transform 1 0 1068 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4729
timestamp 1677677812
transform 1 0 1108 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5289
timestamp 1677677812
transform 1 0 1124 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4629
timestamp 1677677812
transform 1 0 1164 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4678
timestamp 1677677812
transform 1 0 1156 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4730
timestamp 1677677812
transform 1 0 1148 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4679
timestamp 1677677812
transform 1 0 1212 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5186
timestamp 1677677812
transform 1 0 1172 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5187
timestamp 1677677812
transform 1 0 1180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5188
timestamp 1677677812
transform 1 0 1196 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4714
timestamp 1677677812
transform 1 0 1204 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4731
timestamp 1677677812
transform 1 0 1196 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5290
timestamp 1677677812
transform 1 0 1204 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5291
timestamp 1677677812
transform 1 0 1212 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4760
timestamp 1677677812
transform 1 0 1212 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4715
timestamp 1677677812
transform 1 0 1228 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4620
timestamp 1677677812
transform 1 0 1284 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4637
timestamp 1677677812
transform 1 0 1292 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5151
timestamp 1677677812
transform 1 0 1284 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5189
timestamp 1677677812
transform 1 0 1284 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4638
timestamp 1677677812
transform 1 0 1308 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4680
timestamp 1677677812
transform 1 0 1324 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5190
timestamp 1677677812
transform 1 0 1324 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4791
timestamp 1677677812
transform 1 0 1332 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4621
timestamp 1677677812
transform 1 0 1364 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_5152
timestamp 1677677812
transform 1 0 1364 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5292
timestamp 1677677812
transform 1 0 1404 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4761
timestamp 1677677812
transform 1 0 1404 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4681
timestamp 1677677812
transform 1 0 1436 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5191
timestamp 1677677812
transform 1 0 1436 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5293
timestamp 1677677812
transform 1 0 1420 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4682
timestamp 1677677812
transform 1 0 1484 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5294
timestamp 1677677812
transform 1 0 1484 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5295
timestamp 1677677812
transform 1 0 1492 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5192
timestamp 1677677812
transform 1 0 1540 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5296
timestamp 1677677812
transform 1 0 1532 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4639
timestamp 1677677812
transform 1 0 1604 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5193
timestamp 1677677812
transform 1 0 1580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5194
timestamp 1677677812
transform 1 0 1604 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5297
timestamp 1677677812
transform 1 0 1588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4762
timestamp 1677677812
transform 1 0 1580 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5298
timestamp 1677677812
transform 1 0 1652 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4640
timestamp 1677677812
transform 1 0 1692 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4683
timestamp 1677677812
transform 1 0 1676 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5195
timestamp 1677677812
transform 1 0 1676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5196
timestamp 1677677812
transform 1 0 1692 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5299
timestamp 1677677812
transform 1 0 1668 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5300
timestamp 1677677812
transform 1 0 1684 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4763
timestamp 1677677812
transform 1 0 1684 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4684
timestamp 1677677812
transform 1 0 1708 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4622
timestamp 1677677812
transform 1 0 1724 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4623
timestamp 1677677812
transform 1 0 1748 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_5197
timestamp 1677677812
transform 1 0 1740 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5301
timestamp 1677677812
transform 1 0 1732 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4685
timestamp 1677677812
transform 1 0 1780 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4686
timestamp 1677677812
transform 1 0 1804 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5198
timestamp 1677677812
transform 1 0 1780 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5302
timestamp 1677677812
transform 1 0 1828 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4764
timestamp 1677677812
transform 1 0 1780 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4765
timestamp 1677677812
transform 1 0 1812 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5199
timestamp 1677677812
transform 1 0 1844 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4766
timestamp 1677677812
transform 1 0 1844 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4641
timestamp 1677677812
transform 1 0 1932 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5200
timestamp 1677677812
transform 1 0 1932 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4624
timestamp 1677677812
transform 1 0 1964 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_5201
timestamp 1677677812
transform 1 0 1956 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4716
timestamp 1677677812
transform 1 0 1972 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5303
timestamp 1677677812
transform 1 0 1940 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5304
timestamp 1677677812
transform 1 0 1948 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5305
timestamp 1677677812
transform 1 0 1964 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5202
timestamp 1677677812
transform 1 0 1988 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4767
timestamp 1677677812
transform 1 0 1980 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4687
timestamp 1677677812
transform 1 0 2052 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4717
timestamp 1677677812
transform 1 0 2004 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4688
timestamp 1677677812
transform 1 0 2092 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5203
timestamp 1677677812
transform 1 0 2052 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5204
timestamp 1677677812
transform 1 0 2084 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5205
timestamp 1677677812
transform 1 0 2092 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5306
timestamp 1677677812
transform 1 0 2004 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4732
timestamp 1677677812
transform 1 0 2084 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4768
timestamp 1677677812
transform 1 0 2004 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4642
timestamp 1677677812
transform 1 0 2108 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5206
timestamp 1677677812
transform 1 0 2108 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4643
timestamp 1677677812
transform 1 0 2164 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5207
timestamp 1677677812
transform 1 0 2164 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4718
timestamp 1677677812
transform 1 0 2180 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4625
timestamp 1677677812
transform 1 0 2212 0 1 2265
box -3 -3 3 3
use M2_M1  M2_M1_5208
timestamp 1677677812
transform 1 0 2188 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5209
timestamp 1677677812
transform 1 0 2204 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5307
timestamp 1677677812
transform 1 0 2172 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5308
timestamp 1677677812
transform 1 0 2180 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5309
timestamp 1677677812
transform 1 0 2212 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4769
timestamp 1677677812
transform 1 0 2212 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4689
timestamp 1677677812
transform 1 0 2276 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5310
timestamp 1677677812
transform 1 0 2276 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5311
timestamp 1677677812
transform 1 0 2292 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4792
timestamp 1677677812
transform 1 0 2284 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5210
timestamp 1677677812
transform 1 0 2308 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4644
timestamp 1677677812
transform 1 0 2324 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5211
timestamp 1677677812
transform 1 0 2324 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4645
timestamp 1677677812
transform 1 0 2356 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4690
timestamp 1677677812
transform 1 0 2348 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5212
timestamp 1677677812
transform 1 0 2348 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5312
timestamp 1677677812
transform 1 0 2364 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4770
timestamp 1677677812
transform 1 0 2364 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4646
timestamp 1677677812
transform 1 0 2388 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5213
timestamp 1677677812
transform 1 0 2380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5313
timestamp 1677677812
transform 1 0 2388 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4793
timestamp 1677677812
transform 1 0 2420 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4771
timestamp 1677677812
transform 1 0 2460 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5214
timestamp 1677677812
transform 1 0 2476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5215
timestamp 1677677812
transform 1 0 2492 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5216
timestamp 1677677812
transform 1 0 2580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5217
timestamp 1677677812
transform 1 0 2596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5314
timestamp 1677677812
transform 1 0 2572 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4719
timestamp 1677677812
transform 1 0 2628 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5315
timestamp 1677677812
transform 1 0 2628 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5218
timestamp 1677677812
transform 1 0 2676 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5219
timestamp 1677677812
transform 1 0 2732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5316
timestamp 1677677812
transform 1 0 2652 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4720
timestamp 1677677812
transform 1 0 2788 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5220
timestamp 1677677812
transform 1 0 2804 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5317
timestamp 1677677812
transform 1 0 2828 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5153
timestamp 1677677812
transform 1 0 2868 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4721
timestamp 1677677812
transform 1 0 2868 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4722
timestamp 1677677812
transform 1 0 2892 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5318
timestamp 1677677812
transform 1 0 2884 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5319
timestamp 1677677812
transform 1 0 2892 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4772
timestamp 1677677812
transform 1 0 2884 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5154
timestamp 1677677812
transform 1 0 2916 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5155
timestamp 1677677812
transform 1 0 2924 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5221
timestamp 1677677812
transform 1 0 2924 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4733
timestamp 1677677812
transform 1 0 2924 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5222
timestamp 1677677812
transform 1 0 2948 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4734
timestamp 1677677812
transform 1 0 2980 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4773
timestamp 1677677812
transform 1 0 3012 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4626
timestamp 1677677812
transform 1 0 3052 0 1 2265
box -3 -3 3 3
use M3_M2  M3_M2_4691
timestamp 1677677812
transform 1 0 3044 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5223
timestamp 1677677812
transform 1 0 3036 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5224
timestamp 1677677812
transform 1 0 3076 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5320
timestamp 1677677812
transform 1 0 3044 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5321
timestamp 1677677812
transform 1 0 3052 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5322
timestamp 1677677812
transform 1 0 3068 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5323
timestamp 1677677812
transform 1 0 3084 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4774
timestamp 1677677812
transform 1 0 3052 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4692
timestamp 1677677812
transform 1 0 3164 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4693
timestamp 1677677812
transform 1 0 3188 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5225
timestamp 1677677812
transform 1 0 3164 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5226
timestamp 1677677812
transform 1 0 3180 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5227
timestamp 1677677812
transform 1 0 3188 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5324
timestamp 1677677812
transform 1 0 3148 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4735
timestamp 1677677812
transform 1 0 3156 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5325
timestamp 1677677812
transform 1 0 3172 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4736
timestamp 1677677812
transform 1 0 3180 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5326
timestamp 1677677812
transform 1 0 3188 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5327
timestamp 1677677812
transform 1 0 3212 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5228
timestamp 1677677812
transform 1 0 3260 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4630
timestamp 1677677812
transform 1 0 3276 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5328
timestamp 1677677812
transform 1 0 3284 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5156
timestamp 1677677812
transform 1 0 3308 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5147
timestamp 1677677812
transform 1 0 3324 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5229
timestamp 1677677812
transform 1 0 3348 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4737
timestamp 1677677812
transform 1 0 3348 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5230
timestamp 1677677812
transform 1 0 3388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5231
timestamp 1677677812
transform 1 0 3396 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4647
timestamp 1677677812
transform 1 0 3420 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5148
timestamp 1677677812
transform 1 0 3420 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5157
timestamp 1677677812
transform 1 0 3420 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4723
timestamp 1677677812
transform 1 0 3420 0 1 2215
box -3 -3 3 3
use M3_M2  M3_M2_4694
timestamp 1677677812
transform 1 0 3460 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4648
timestamp 1677677812
transform 1 0 3484 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5232
timestamp 1677677812
transform 1 0 3476 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5329
timestamp 1677677812
transform 1 0 3468 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4775
timestamp 1677677812
transform 1 0 3476 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4695
timestamp 1677677812
transform 1 0 3524 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5233
timestamp 1677677812
transform 1 0 3500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5234
timestamp 1677677812
transform 1 0 3516 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5235
timestamp 1677677812
transform 1 0 3524 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5330
timestamp 1677677812
transform 1 0 3492 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4738
timestamp 1677677812
transform 1 0 3500 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4776
timestamp 1677677812
transform 1 0 3492 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4696
timestamp 1677677812
transform 1 0 3540 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4739
timestamp 1677677812
transform 1 0 3532 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4649
timestamp 1677677812
transform 1 0 3596 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4697
timestamp 1677677812
transform 1 0 3572 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4698
timestamp 1677677812
transform 1 0 3588 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5236
timestamp 1677677812
transform 1 0 3572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5237
timestamp 1677677812
transform 1 0 3588 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5331
timestamp 1677677812
transform 1 0 3540 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5332
timestamp 1677677812
transform 1 0 3548 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4740
timestamp 1677677812
transform 1 0 3556 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5333
timestamp 1677677812
transform 1 0 3564 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5334
timestamp 1677677812
transform 1 0 3580 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4794
timestamp 1677677812
transform 1 0 3548 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4650
timestamp 1677677812
transform 1 0 3636 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5335
timestamp 1677677812
transform 1 0 3620 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5336
timestamp 1677677812
transform 1 0 3628 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4795
timestamp 1677677812
transform 1 0 3628 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5238
timestamp 1677677812
transform 1 0 3644 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5239
timestamp 1677677812
transform 1 0 3660 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5337
timestamp 1677677812
transform 1 0 3652 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4741
timestamp 1677677812
transform 1 0 3660 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4777
timestamp 1677677812
transform 1 0 3652 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5338
timestamp 1677677812
transform 1 0 3684 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5240
timestamp 1677677812
transform 1 0 3732 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5339
timestamp 1677677812
transform 1 0 3708 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4778
timestamp 1677677812
transform 1 0 3732 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5241
timestamp 1677677812
transform 1 0 3804 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4742
timestamp 1677677812
transform 1 0 3804 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4796
timestamp 1677677812
transform 1 0 3804 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5363
timestamp 1677677812
transform 1 0 3812 0 1 2185
box -2 -2 2 2
use M2_M1  M2_M1_5242
timestamp 1677677812
transform 1 0 3828 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5243
timestamp 1677677812
transform 1 0 3844 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4651
timestamp 1677677812
transform 1 0 3900 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5244
timestamp 1677677812
transform 1 0 3868 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5245
timestamp 1677677812
transform 1 0 3884 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5340
timestamp 1677677812
transform 1 0 3836 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5341
timestamp 1677677812
transform 1 0 3852 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5342
timestamp 1677677812
transform 1 0 3860 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4743
timestamp 1677677812
transform 1 0 3868 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5343
timestamp 1677677812
transform 1 0 3876 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4779
timestamp 1677677812
transform 1 0 3876 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4652
timestamp 1677677812
transform 1 0 3924 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4699
timestamp 1677677812
transform 1 0 3924 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4653
timestamp 1677677812
transform 1 0 3964 0 1 2245
box -3 -3 3 3
use M2_M1  M2_M1_5246
timestamp 1677677812
transform 1 0 3932 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5247
timestamp 1677677812
transform 1 0 3948 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5344
timestamp 1677677812
transform 1 0 3924 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4780
timestamp 1677677812
transform 1 0 3916 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4724
timestamp 1677677812
transform 1 0 3956 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5248
timestamp 1677677812
transform 1 0 3964 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5249
timestamp 1677677812
transform 1 0 3972 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5345
timestamp 1677677812
transform 1 0 3940 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4744
timestamp 1677677812
transform 1 0 3964 0 1 2205
box -3 -3 3 3
use M3_M2  M3_M2_4781
timestamp 1677677812
transform 1 0 3940 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4700
timestamp 1677677812
transform 1 0 4028 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5250
timestamp 1677677812
transform 1 0 3996 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5251
timestamp 1677677812
transform 1 0 4012 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5252
timestamp 1677677812
transform 1 0 4028 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5346
timestamp 1677677812
transform 1 0 3996 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5347
timestamp 1677677812
transform 1 0 4020 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4797
timestamp 1677677812
transform 1 0 3988 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4745
timestamp 1677677812
transform 1 0 4028 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5253
timestamp 1677677812
transform 1 0 4044 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5348
timestamp 1677677812
transform 1 0 4060 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5254
timestamp 1677677812
transform 1 0 4116 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4746
timestamp 1677677812
transform 1 0 4116 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5349
timestamp 1677677812
transform 1 0 4164 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4662
timestamp 1677677812
transform 1 0 4228 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5149
timestamp 1677677812
transform 1 0 4236 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5158
timestamp 1677677812
transform 1 0 4228 0 1 2225
box -2 -2 2 2
use M3_M2  M3_M2_4782
timestamp 1677677812
transform 1 0 4228 0 1 2195
box -3 -3 3 3
use M2_M1  M2_M1_5159
timestamp 1677677812
transform 1 0 4252 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5150
timestamp 1677677812
transform 1 0 4308 0 1 2235
box -2 -2 2 2
use M2_M1  M2_M1_5255
timestamp 1677677812
transform 1 0 4308 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4747
timestamp 1677677812
transform 1 0 4308 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5160
timestamp 1677677812
transform 1 0 4324 0 1 2225
box -2 -2 2 2
use M2_M1  M2_M1_5256
timestamp 1677677812
transform 1 0 4332 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4725
timestamp 1677677812
transform 1 0 4340 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5257
timestamp 1677677812
transform 1 0 4348 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4726
timestamp 1677677812
transform 1 0 4356 0 1 2215
box -3 -3 3 3
use M2_M1  M2_M1_5350
timestamp 1677677812
transform 1 0 4332 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4654
timestamp 1677677812
transform 1 0 4380 0 1 2245
box -3 -3 3 3
use M3_M2  M3_M2_4701
timestamp 1677677812
transform 1 0 4396 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5258
timestamp 1677677812
transform 1 0 4380 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5259
timestamp 1677677812
transform 1 0 4388 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5351
timestamp 1677677812
transform 1 0 4396 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4783
timestamp 1677677812
transform 1 0 4396 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4702
timestamp 1677677812
transform 1 0 4428 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5260
timestamp 1677677812
transform 1 0 4412 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5261
timestamp 1677677812
transform 1 0 4428 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5352
timestamp 1677677812
transform 1 0 4420 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5353
timestamp 1677677812
transform 1 0 4436 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4784
timestamp 1677677812
transform 1 0 4420 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4798
timestamp 1677677812
transform 1 0 4420 0 1 2185
box -3 -3 3 3
use M2_M1  M2_M1_5354
timestamp 1677677812
transform 1 0 4452 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4631
timestamp 1677677812
transform 1 0 4508 0 1 2255
box -3 -3 3 3
use M2_M1  M2_M1_5262
timestamp 1677677812
transform 1 0 4500 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5355
timestamp 1677677812
transform 1 0 4476 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4785
timestamp 1677677812
transform 1 0 4500 0 1 2195
box -3 -3 3 3
use M3_M2  M3_M2_4663
timestamp 1677677812
transform 1 0 4588 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4664
timestamp 1677677812
transform 1 0 4612 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4703
timestamp 1677677812
transform 1 0 4572 0 1 2225
box -3 -3 3 3
use M3_M2  M3_M2_4704
timestamp 1677677812
transform 1 0 4604 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5263
timestamp 1677677812
transform 1 0 4572 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5264
timestamp 1677677812
transform 1 0 4580 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5265
timestamp 1677677812
transform 1 0 4596 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5266
timestamp 1677677812
transform 1 0 4612 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5356
timestamp 1677677812
transform 1 0 4588 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4748
timestamp 1677677812
transform 1 0 4596 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5357
timestamp 1677677812
transform 1 0 4604 0 1 2205
box -2 -2 2 2
use M2_M1  M2_M1_5267
timestamp 1677677812
transform 1 0 4636 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5358
timestamp 1677677812
transform 1 0 4628 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4749
timestamp 1677677812
transform 1 0 4644 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5359
timestamp 1677677812
transform 1 0 4652 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4665
timestamp 1677677812
transform 1 0 4668 0 1 2235
box -3 -3 3 3
use M3_M2  M3_M2_4705
timestamp 1677677812
transform 1 0 4684 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5268
timestamp 1677677812
transform 1 0 4668 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5269
timestamp 1677677812
transform 1 0 4684 0 1 2215
box -2 -2 2 2
use M3_M2  M3_M2_4750
timestamp 1677677812
transform 1 0 4668 0 1 2205
box -3 -3 3 3
use M2_M1  M2_M1_5360
timestamp 1677677812
transform 1 0 4676 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4706
timestamp 1677677812
transform 1 0 4700 0 1 2225
box -3 -3 3 3
use M2_M1  M2_M1_5270
timestamp 1677677812
transform 1 0 4700 0 1 2215
box -2 -2 2 2
use M2_M1  M2_M1_5361
timestamp 1677677812
transform 1 0 4708 0 1 2205
box -2 -2 2 2
use M3_M2  M3_M2_4799
timestamp 1677677812
transform 1 0 4716 0 1 2185
box -3 -3 3 3
use M3_M2  M3_M2_4632
timestamp 1677677812
transform 1 0 4740 0 1 2255
box -3 -3 3 3
use M3_M2  M3_M2_4666
timestamp 1677677812
transform 1 0 4732 0 1 2235
box -3 -3 3 3
use M2_M1  M2_M1_5362
timestamp 1677677812
transform 1 0 4788 0 1 2205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_50
timestamp 1677677812
transform 1 0 48 0 1 2170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_345
timestamp 1677677812
transform 1 0 72 0 1 2170
box -8 -3 104 105
use FILL  FILL_5893
timestamp 1677677812
transform 1 0 168 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_389
timestamp 1677677812
transform 1 0 176 0 1 2170
box -9 -3 26 105
use FILL  FILL_5905
timestamp 1677677812
transform 1 0 192 0 1 2170
box -8 -3 16 105
use FILL  FILL_5909
timestamp 1677677812
transform 1 0 200 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_346
timestamp 1677677812
transform 1 0 208 0 1 2170
box -8 -3 104 105
use FILL  FILL_5911
timestamp 1677677812
transform 1 0 304 0 1 2170
box -8 -3 16 105
use FILL  FILL_5912
timestamp 1677677812
transform 1 0 312 0 1 2170
box -8 -3 16 105
use FILL  FILL_5913
timestamp 1677677812
transform 1 0 320 0 1 2170
box -8 -3 16 105
use FILL  FILL_5914
timestamp 1677677812
transform 1 0 328 0 1 2170
box -8 -3 16 105
use FILL  FILL_5915
timestamp 1677677812
transform 1 0 336 0 1 2170
box -8 -3 16 105
use FILL  FILL_5916
timestamp 1677677812
transform 1 0 344 0 1 2170
box -8 -3 16 105
use FILL  FILL_5917
timestamp 1677677812
transform 1 0 352 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_390
timestamp 1677677812
transform -1 0 376 0 1 2170
box -9 -3 26 105
use FILL  FILL_5918
timestamp 1677677812
transform 1 0 376 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_238
timestamp 1677677812
transform 1 0 384 0 1 2170
box -8 -3 46 105
use FILL  FILL_5927
timestamp 1677677812
transform 1 0 424 0 1 2170
box -8 -3 16 105
use FILL  FILL_5928
timestamp 1677677812
transform 1 0 432 0 1 2170
box -8 -3 16 105
use FILL  FILL_5929
timestamp 1677677812
transform 1 0 440 0 1 2170
box -8 -3 16 105
use FILL  FILL_5930
timestamp 1677677812
transform 1 0 448 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_239
timestamp 1677677812
transform 1 0 456 0 1 2170
box -8 -3 46 105
use FILL  FILL_5931
timestamp 1677677812
transform 1 0 496 0 1 2170
box -8 -3 16 105
use FILL  FILL_5942
timestamp 1677677812
transform 1 0 504 0 1 2170
box -8 -3 16 105
use FILL  FILL_5944
timestamp 1677677812
transform 1 0 512 0 1 2170
box -8 -3 16 105
use FILL  FILL_5945
timestamp 1677677812
transform 1 0 520 0 1 2170
box -8 -3 16 105
use FILL  FILL_5946
timestamp 1677677812
transform 1 0 528 0 1 2170
box -8 -3 16 105
use FILL  FILL_5947
timestamp 1677677812
transform 1 0 536 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_392
timestamp 1677677812
transform 1 0 544 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_348
timestamp 1677677812
transform -1 0 656 0 1 2170
box -8 -3 104 105
use FILL  FILL_5948
timestamp 1677677812
transform 1 0 656 0 1 2170
box -8 -3 16 105
use FILL  FILL_5949
timestamp 1677677812
transform 1 0 664 0 1 2170
box -8 -3 16 105
use FILL  FILL_5958
timestamp 1677677812
transform 1 0 672 0 1 2170
box -8 -3 16 105
use FILL  FILL_5960
timestamp 1677677812
transform 1 0 680 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_393
timestamp 1677677812
transform 1 0 688 0 1 2170
box -9 -3 26 105
use FILL  FILL_5962
timestamp 1677677812
transform 1 0 704 0 1 2170
box -8 -3 16 105
use FILL  FILL_5963
timestamp 1677677812
transform 1 0 712 0 1 2170
box -8 -3 16 105
use FILL  FILL_5964
timestamp 1677677812
transform 1 0 720 0 1 2170
box -8 -3 16 105
use FILL  FILL_5965
timestamp 1677677812
transform 1 0 728 0 1 2170
box -8 -3 16 105
use FILL  FILL_5966
timestamp 1677677812
transform 1 0 736 0 1 2170
box -8 -3 16 105
use FILL  FILL_5970
timestamp 1677677812
transform 1 0 744 0 1 2170
box -8 -3 16 105
use FILL  FILL_5972
timestamp 1677677812
transform 1 0 752 0 1 2170
box -8 -3 16 105
use FILL  FILL_5974
timestamp 1677677812
transform 1 0 760 0 1 2170
box -8 -3 16 105
use FILL  FILL_5976
timestamp 1677677812
transform 1 0 768 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_240
timestamp 1677677812
transform -1 0 816 0 1 2170
box -8 -3 46 105
use FILL  FILL_5977
timestamp 1677677812
transform 1 0 816 0 1 2170
box -8 -3 16 105
use FILL  FILL_5985
timestamp 1677677812
transform 1 0 824 0 1 2170
box -8 -3 16 105
use FILL  FILL_5986
timestamp 1677677812
transform 1 0 832 0 1 2170
box -8 -3 16 105
use FILL  FILL_5987
timestamp 1677677812
transform 1 0 840 0 1 2170
box -8 -3 16 105
use FILL  FILL_5988
timestamp 1677677812
transform 1 0 848 0 1 2170
box -8 -3 16 105
use FILL  FILL_5989
timestamp 1677677812
transform 1 0 856 0 1 2170
box -8 -3 16 105
use FILL  FILL_5990
timestamp 1677677812
transform 1 0 864 0 1 2170
box -8 -3 16 105
use FILL  FILL_5992
timestamp 1677677812
transform 1 0 872 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_242
timestamp 1677677812
transform -1 0 920 0 1 2170
box -8 -3 46 105
use FILL  FILL_5993
timestamp 1677677812
transform 1 0 920 0 1 2170
box -8 -3 16 105
use FILL  FILL_5994
timestamp 1677677812
transform 1 0 928 0 1 2170
box -8 -3 16 105
use FILL  FILL_5995
timestamp 1677677812
transform 1 0 936 0 1 2170
box -8 -3 16 105
use FILL  FILL_6002
timestamp 1677677812
transform 1 0 944 0 1 2170
box -8 -3 16 105
use FILL  FILL_6004
timestamp 1677677812
transform 1 0 952 0 1 2170
box -8 -3 16 105
use FILL  FILL_6006
timestamp 1677677812
transform 1 0 960 0 1 2170
box -8 -3 16 105
use FILL  FILL_6008
timestamp 1677677812
transform 1 0 968 0 1 2170
box -8 -3 16 105
use FILL  FILL_6010
timestamp 1677677812
transform 1 0 976 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_243
timestamp 1677677812
transform 1 0 984 0 1 2170
box -8 -3 46 105
use FILL  FILL_6011
timestamp 1677677812
transform 1 0 1024 0 1 2170
box -8 -3 16 105
use FILL  FILL_6015
timestamp 1677677812
transform 1 0 1032 0 1 2170
box -8 -3 16 105
use FILL  FILL_6017
timestamp 1677677812
transform 1 0 1040 0 1 2170
box -8 -3 16 105
use FILL  FILL_6019
timestamp 1677677812
transform 1 0 1048 0 1 2170
box -8 -3 16 105
use FILL  FILL_6021
timestamp 1677677812
transform 1 0 1056 0 1 2170
box -8 -3 16 105
use FILL  FILL_6023
timestamp 1677677812
transform 1 0 1064 0 1 2170
box -8 -3 16 105
use FILL  FILL_6024
timestamp 1677677812
transform 1 0 1072 0 1 2170
box -8 -3 16 105
use FILL  FILL_6025
timestamp 1677677812
transform 1 0 1080 0 1 2170
box -8 -3 16 105
use FILL  FILL_6026
timestamp 1677677812
transform 1 0 1088 0 1 2170
box -8 -3 16 105
use FILL  FILL_6027
timestamp 1677677812
transform 1 0 1096 0 1 2170
box -8 -3 16 105
use FILL  FILL_6028
timestamp 1677677812
transform 1 0 1104 0 1 2170
box -8 -3 16 105
use FILL  FILL_6031
timestamp 1677677812
transform 1 0 1112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6033
timestamp 1677677812
transform 1 0 1120 0 1 2170
box -8 -3 16 105
use FILL  FILL_6035
timestamp 1677677812
transform 1 0 1128 0 1 2170
box -8 -3 16 105
use FILL  FILL_6037
timestamp 1677677812
transform 1 0 1136 0 1 2170
box -8 -3 16 105
use FILL  FILL_6039
timestamp 1677677812
transform 1 0 1144 0 1 2170
box -8 -3 16 105
use FILL  FILL_6041
timestamp 1677677812
transform 1 0 1152 0 1 2170
box -8 -3 16 105
use FILL  FILL_6043
timestamp 1677677812
transform 1 0 1160 0 1 2170
box -8 -3 16 105
use FILL  FILL_6045
timestamp 1677677812
transform 1 0 1168 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4800
timestamp 1677677812
transform 1 0 1204 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_244
timestamp 1677677812
transform -1 0 1216 0 1 2170
box -8 -3 46 105
use FILL  FILL_6046
timestamp 1677677812
transform 1 0 1216 0 1 2170
box -8 -3 16 105
use FILL  FILL_6054
timestamp 1677677812
transform 1 0 1224 0 1 2170
box -8 -3 16 105
use FILL  FILL_6056
timestamp 1677677812
transform 1 0 1232 0 1 2170
box -8 -3 16 105
use FILL  FILL_6058
timestamp 1677677812
transform 1 0 1240 0 1 2170
box -8 -3 16 105
use FILL  FILL_6059
timestamp 1677677812
transform 1 0 1248 0 1 2170
box -8 -3 16 105
use FILL  FILL_6060
timestamp 1677677812
transform 1 0 1256 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4801
timestamp 1677677812
transform 1 0 1276 0 1 2175
box -3 -3 3 3
use FILL  FILL_6061
timestamp 1677677812
transform 1 0 1264 0 1 2170
box -8 -3 16 105
use FILL  FILL_6062
timestamp 1677677812
transform 1 0 1272 0 1 2170
box -8 -3 16 105
use FILL  FILL_6063
timestamp 1677677812
transform 1 0 1280 0 1 2170
box -8 -3 16 105
use FILL  FILL_6064
timestamp 1677677812
transform 1 0 1288 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_119
timestamp 1677677812
transform -1 0 1328 0 1 2170
box -8 -3 34 105
use FILL  FILL_6065
timestamp 1677677812
transform 1 0 1328 0 1 2170
box -8 -3 16 105
use FILL  FILL_6073
timestamp 1677677812
transform 1 0 1336 0 1 2170
box -8 -3 16 105
use FILL  FILL_6075
timestamp 1677677812
transform 1 0 1344 0 1 2170
box -8 -3 16 105
use FILL  FILL_6077
timestamp 1677677812
transform 1 0 1352 0 1 2170
box -8 -3 16 105
use FILL  FILL_6079
timestamp 1677677812
transform 1 0 1360 0 1 2170
box -8 -3 16 105
use FILL  FILL_6081
timestamp 1677677812
transform 1 0 1368 0 1 2170
box -8 -3 16 105
use FILL  FILL_6083
timestamp 1677677812
transform 1 0 1376 0 1 2170
box -8 -3 16 105
use FILL  FILL_6085
timestamp 1677677812
transform 1 0 1384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6086
timestamp 1677677812
transform 1 0 1392 0 1 2170
box -8 -3 16 105
use FILL  FILL_6087
timestamp 1677677812
transform 1 0 1400 0 1 2170
box -8 -3 16 105
use FILL  FILL_6088
timestamp 1677677812
transform 1 0 1408 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4802
timestamp 1677677812
transform 1 0 1436 0 1 2175
box -3 -3 3 3
use OAI21X1  OAI21X1_120
timestamp 1677677812
transform -1 0 1448 0 1 2170
box -8 -3 34 105
use FILL  FILL_6089
timestamp 1677677812
transform 1 0 1448 0 1 2170
box -8 -3 16 105
use FILL  FILL_6095
timestamp 1677677812
transform 1 0 1456 0 1 2170
box -8 -3 16 105
use FILL  FILL_6097
timestamp 1677677812
transform 1 0 1464 0 1 2170
box -8 -3 16 105
use FILL  FILL_6099
timestamp 1677677812
transform 1 0 1472 0 1 2170
box -8 -3 16 105
use FILL  FILL_6101
timestamp 1677677812
transform 1 0 1480 0 1 2170
box -8 -3 16 105
use FILL  FILL_6103
timestamp 1677677812
transform 1 0 1488 0 1 2170
box -8 -3 16 105
use FILL  FILL_6105
timestamp 1677677812
transform 1 0 1496 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_394
timestamp 1677677812
transform 1 0 1504 0 1 2170
box -9 -3 26 105
use FILL  FILL_6106
timestamp 1677677812
transform 1 0 1520 0 1 2170
box -8 -3 16 105
use FILL  FILL_6108
timestamp 1677677812
transform 1 0 1528 0 1 2170
box -8 -3 16 105
use FILL  FILL_6110
timestamp 1677677812
transform 1 0 1536 0 1 2170
box -8 -3 16 105
use FILL  FILL_6112
timestamp 1677677812
transform 1 0 1544 0 1 2170
box -8 -3 16 105
use FILL  FILL_6113
timestamp 1677677812
transform 1 0 1552 0 1 2170
box -8 -3 16 105
use FILL  FILL_6114
timestamp 1677677812
transform 1 0 1560 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_230
timestamp 1677677812
transform -1 0 1608 0 1 2170
box -8 -3 46 105
use FILL  FILL_6115
timestamp 1677677812
transform 1 0 1608 0 1 2170
box -8 -3 16 105
use FILL  FILL_6116
timestamp 1677677812
transform 1 0 1616 0 1 2170
box -8 -3 16 105
use FILL  FILL_6117
timestamp 1677677812
transform 1 0 1624 0 1 2170
box -8 -3 16 105
use FILL  FILL_6118
timestamp 1677677812
transform 1 0 1632 0 1 2170
box -8 -3 16 105
use FILL  FILL_6119
timestamp 1677677812
transform 1 0 1640 0 1 2170
box -8 -3 16 105
use FILL  FILL_6121
timestamp 1677677812
transform 1 0 1648 0 1 2170
box -8 -3 16 105
use FILL  FILL_6123
timestamp 1677677812
transform 1 0 1656 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_231
timestamp 1677677812
transform -1 0 1704 0 1 2170
box -8 -3 46 105
use FILL  FILL_6124
timestamp 1677677812
transform 1 0 1704 0 1 2170
box -8 -3 16 105
use FILL  FILL_6125
timestamp 1677677812
transform 1 0 1712 0 1 2170
box -8 -3 16 105
use FILL  FILL_6126
timestamp 1677677812
transform 1 0 1720 0 1 2170
box -8 -3 16 105
use FILL  FILL_6127
timestamp 1677677812
transform 1 0 1728 0 1 2170
box -8 -3 16 105
use FILL  FILL_6132
timestamp 1677677812
transform 1 0 1736 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_350
timestamp 1677677812
transform -1 0 1840 0 1 2170
box -8 -3 104 105
use FILL  FILL_6133
timestamp 1677677812
transform 1 0 1840 0 1 2170
box -8 -3 16 105
use FILL  FILL_6134
timestamp 1677677812
transform 1 0 1848 0 1 2170
box -8 -3 16 105
use FILL  FILL_6138
timestamp 1677677812
transform 1 0 1856 0 1 2170
box -8 -3 16 105
use FILL  FILL_6140
timestamp 1677677812
transform 1 0 1864 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_396
timestamp 1677677812
transform -1 0 1888 0 1 2170
box -9 -3 26 105
use FILL  FILL_6141
timestamp 1677677812
transform 1 0 1888 0 1 2170
box -8 -3 16 105
use FILL  FILL_6146
timestamp 1677677812
transform 1 0 1896 0 1 2170
box -8 -3 16 105
use FILL  FILL_6148
timestamp 1677677812
transform 1 0 1904 0 1 2170
box -8 -3 16 105
use FILL  FILL_6149
timestamp 1677677812
transform 1 0 1912 0 1 2170
box -8 -3 16 105
use FILL  FILL_6150
timestamp 1677677812
transform 1 0 1920 0 1 2170
box -8 -3 16 105
use FILL  FILL_6151
timestamp 1677677812
transform 1 0 1928 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_246
timestamp 1677677812
transform -1 0 1976 0 1 2170
box -8 -3 46 105
use FILL  FILL_6152
timestamp 1677677812
transform 1 0 1976 0 1 2170
box -8 -3 16 105
use FILL  FILL_6158
timestamp 1677677812
transform 1 0 1984 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_352
timestamp 1677677812
transform 1 0 1992 0 1 2170
box -8 -3 104 105
use FILL  FILL_6160
timestamp 1677677812
transform 1 0 2088 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_397
timestamp 1677677812
transform -1 0 2112 0 1 2170
box -9 -3 26 105
use FILL  FILL_6161
timestamp 1677677812
transform 1 0 2112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6173
timestamp 1677677812
transform 1 0 2120 0 1 2170
box -8 -3 16 105
use FILL  FILL_6175
timestamp 1677677812
transform 1 0 2128 0 1 2170
box -8 -3 16 105
use FILL  FILL_6177
timestamp 1677677812
transform 1 0 2136 0 1 2170
box -8 -3 16 105
use FILL  FILL_6179
timestamp 1677677812
transform 1 0 2144 0 1 2170
box -8 -3 16 105
use FILL  FILL_6181
timestamp 1677677812
transform 1 0 2152 0 1 2170
box -8 -3 16 105
use FILL  FILL_6183
timestamp 1677677812
transform 1 0 2160 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_247
timestamp 1677677812
transform -1 0 2208 0 1 2170
box -8 -3 46 105
use FILL  FILL_6184
timestamp 1677677812
transform 1 0 2208 0 1 2170
box -8 -3 16 105
use FILL  FILL_6187
timestamp 1677677812
transform 1 0 2216 0 1 2170
box -8 -3 16 105
use FILL  FILL_6189
timestamp 1677677812
transform 1 0 2224 0 1 2170
box -8 -3 16 105
use FILL  FILL_6191
timestamp 1677677812
transform 1 0 2232 0 1 2170
box -8 -3 16 105
use FILL  FILL_6193
timestamp 1677677812
transform 1 0 2240 0 1 2170
box -8 -3 16 105
use FILL  FILL_6195
timestamp 1677677812
transform 1 0 2248 0 1 2170
box -8 -3 16 105
use FILL  FILL_6197
timestamp 1677677812
transform 1 0 2256 0 1 2170
box -8 -3 16 105
use FILL  FILL_6199
timestamp 1677677812
transform 1 0 2264 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_398
timestamp 1677677812
transform 1 0 2272 0 1 2170
box -9 -3 26 105
use FILL  FILL_6201
timestamp 1677677812
transform 1 0 2288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6202
timestamp 1677677812
transform 1 0 2296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6203
timestamp 1677677812
transform 1 0 2304 0 1 2170
box -8 -3 16 105
use FILL  FILL_6204
timestamp 1677677812
transform 1 0 2312 0 1 2170
box -8 -3 16 105
use FILL  FILL_6205
timestamp 1677677812
transform 1 0 2320 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_248
timestamp 1677677812
transform -1 0 2368 0 1 2170
box -8 -3 46 105
use FILL  FILL_6206
timestamp 1677677812
transform 1 0 2368 0 1 2170
box -8 -3 16 105
use FILL  FILL_6208
timestamp 1677677812
transform 1 0 2376 0 1 2170
box -8 -3 16 105
use FILL  FILL_6210
timestamp 1677677812
transform 1 0 2384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6212
timestamp 1677677812
transform 1 0 2392 0 1 2170
box -8 -3 16 105
use FILL  FILL_6214
timestamp 1677677812
transform 1 0 2400 0 1 2170
box -8 -3 16 105
use FILL  FILL_6216
timestamp 1677677812
transform 1 0 2408 0 1 2170
box -8 -3 16 105
use FILL  FILL_6217
timestamp 1677677812
transform 1 0 2416 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_399
timestamp 1677677812
transform 1 0 2424 0 1 2170
box -9 -3 26 105
use FILL  FILL_6218
timestamp 1677677812
transform 1 0 2440 0 1 2170
box -8 -3 16 105
use FILL  FILL_6219
timestamp 1677677812
transform 1 0 2448 0 1 2170
box -8 -3 16 105
use FILL  FILL_6222
timestamp 1677677812
transform 1 0 2456 0 1 2170
box -8 -3 16 105
use FILL  FILL_6224
timestamp 1677677812
transform 1 0 2464 0 1 2170
box -8 -3 16 105
use FILL  FILL_6226
timestamp 1677677812
transform 1 0 2472 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4803
timestamp 1677677812
transform 1 0 2492 0 1 2175
box -3 -3 3 3
use FILL  FILL_6228
timestamp 1677677812
transform 1 0 2480 0 1 2170
box -8 -3 16 105
use FILL  FILL_6229
timestamp 1677677812
transform 1 0 2488 0 1 2170
box -8 -3 16 105
use FILL  FILL_6230
timestamp 1677677812
transform 1 0 2496 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4804
timestamp 1677677812
transform 1 0 2516 0 1 2175
box -3 -3 3 3
use FILL  FILL_6231
timestamp 1677677812
transform 1 0 2504 0 1 2170
box -8 -3 16 105
use FILL  FILL_6232
timestamp 1677677812
transform 1 0 2512 0 1 2170
box -8 -3 16 105
use FILL  FILL_6233
timestamp 1677677812
transform 1 0 2520 0 1 2170
box -8 -3 16 105
use FILL  FILL_6236
timestamp 1677677812
transform 1 0 2528 0 1 2170
box -8 -3 16 105
use FILL  FILL_6238
timestamp 1677677812
transform 1 0 2536 0 1 2170
box -8 -3 16 105
use FILL  FILL_6240
timestamp 1677677812
transform 1 0 2544 0 1 2170
box -8 -3 16 105
use FILL  FILL_6242
timestamp 1677677812
transform 1 0 2552 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_249
timestamp 1677677812
transform 1 0 2560 0 1 2170
box -8 -3 46 105
use FILL  FILL_6244
timestamp 1677677812
transform 1 0 2600 0 1 2170
box -8 -3 16 105
use FILL  FILL_6249
timestamp 1677677812
transform 1 0 2608 0 1 2170
box -8 -3 16 105
use FILL  FILL_6251
timestamp 1677677812
transform 1 0 2616 0 1 2170
box -8 -3 16 105
use FILL  FILL_6253
timestamp 1677677812
transform 1 0 2624 0 1 2170
box -8 -3 16 105
use FILL  FILL_6254
timestamp 1677677812
transform 1 0 2632 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_354
timestamp 1677677812
transform 1 0 2640 0 1 2170
box -8 -3 104 105
use FILL  FILL_6255
timestamp 1677677812
transform 1 0 2736 0 1 2170
box -8 -3 16 105
use FILL  FILL_6266
timestamp 1677677812
transform 1 0 2744 0 1 2170
box -8 -3 16 105
use FILL  FILL_6268
timestamp 1677677812
transform 1 0 2752 0 1 2170
box -8 -3 16 105
use FILL  FILL_6269
timestamp 1677677812
transform 1 0 2760 0 1 2170
box -8 -3 16 105
use FILL  FILL_6270
timestamp 1677677812
transform 1 0 2768 0 1 2170
box -8 -3 16 105
use FILL  FILL_6271
timestamp 1677677812
transform 1 0 2776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6273
timestamp 1677677812
transform 1 0 2784 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_122
timestamp 1677677812
transform 1 0 2792 0 1 2170
box -8 -3 34 105
use FILL  FILL_6275
timestamp 1677677812
transform 1 0 2824 0 1 2170
box -8 -3 16 105
use FILL  FILL_6281
timestamp 1677677812
transform 1 0 2832 0 1 2170
box -8 -3 16 105
use FILL  FILL_6283
timestamp 1677677812
transform 1 0 2840 0 1 2170
box -8 -3 16 105
use FILL  FILL_6284
timestamp 1677677812
transform 1 0 2848 0 1 2170
box -8 -3 16 105
use FILL  FILL_6285
timestamp 1677677812
transform 1 0 2856 0 1 2170
box -8 -3 16 105
use FILL  FILL_6286
timestamp 1677677812
transform 1 0 2864 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_401
timestamp 1677677812
transform -1 0 2888 0 1 2170
box -9 -3 26 105
use M3_M2  M3_M2_4805
timestamp 1677677812
transform 1 0 2900 0 1 2175
box -3 -3 3 3
use FILL  FILL_6287
timestamp 1677677812
transform 1 0 2888 0 1 2170
box -8 -3 16 105
use FILL  FILL_6292
timestamp 1677677812
transform 1 0 2896 0 1 2170
box -8 -3 16 105
use FILL  FILL_6293
timestamp 1677677812
transform 1 0 2904 0 1 2170
box -8 -3 16 105
use FILL  FILL_6294
timestamp 1677677812
transform 1 0 2912 0 1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_123
timestamp 1677677812
transform -1 0 2952 0 1 2170
box -8 -3 34 105
use FILL  FILL_6295
timestamp 1677677812
transform 1 0 2952 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4806
timestamp 1677677812
transform 1 0 2972 0 1 2175
box -3 -3 3 3
use FILL  FILL_6300
timestamp 1677677812
transform 1 0 2960 0 1 2170
box -8 -3 16 105
use FILL  FILL_6301
timestamp 1677677812
transform 1 0 2968 0 1 2170
box -8 -3 16 105
use FILL  FILL_6302
timestamp 1677677812
transform 1 0 2976 0 1 2170
box -8 -3 16 105
use FILL  FILL_6303
timestamp 1677677812
transform 1 0 2984 0 1 2170
box -8 -3 16 105
use FILL  FILL_6304
timestamp 1677677812
transform 1 0 2992 0 1 2170
box -8 -3 16 105
use FILL  FILL_6305
timestamp 1677677812
transform 1 0 3000 0 1 2170
box -8 -3 16 105
use FILL  FILL_6306
timestamp 1677677812
transform 1 0 3008 0 1 2170
box -8 -3 16 105
use FILL  FILL_6309
timestamp 1677677812
transform 1 0 3016 0 1 2170
box -8 -3 16 105
use FILL  FILL_6310
timestamp 1677677812
transform 1 0 3024 0 1 2170
box -8 -3 16 105
use FILL  FILL_6311
timestamp 1677677812
transform 1 0 3032 0 1 2170
box -8 -3 16 105
use FILL  FILL_6312
timestamp 1677677812
transform 1 0 3040 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4807
timestamp 1677677812
transform 1 0 3084 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_236
timestamp 1677677812
transform 1 0 3048 0 1 2170
box -8 -3 46 105
use FILL  FILL_6313
timestamp 1677677812
transform 1 0 3088 0 1 2170
box -8 -3 16 105
use FILL  FILL_6314
timestamp 1677677812
transform 1 0 3096 0 1 2170
box -8 -3 16 105
use FILL  FILL_6315
timestamp 1677677812
transform 1 0 3104 0 1 2170
box -8 -3 16 105
use FILL  FILL_6316
timestamp 1677677812
transform 1 0 3112 0 1 2170
box -8 -3 16 105
use FILL  FILL_6317
timestamp 1677677812
transform 1 0 3120 0 1 2170
box -8 -3 16 105
use FILL  FILL_6318
timestamp 1677677812
transform 1 0 3128 0 1 2170
box -8 -3 16 105
use FILL  FILL_6319
timestamp 1677677812
transform 1 0 3136 0 1 2170
box -8 -3 16 105
use FILL  FILL_6320
timestamp 1677677812
transform 1 0 3144 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_237
timestamp 1677677812
transform -1 0 3192 0 1 2170
box -8 -3 46 105
use FILL  FILL_6321
timestamp 1677677812
transform 1 0 3192 0 1 2170
box -8 -3 16 105
use FILL  FILL_6322
timestamp 1677677812
transform 1 0 3200 0 1 2170
box -8 -3 16 105
use FILL  FILL_6323
timestamp 1677677812
transform 1 0 3208 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_402
timestamp 1677677812
transform 1 0 3216 0 1 2170
box -9 -3 26 105
use FILL  FILL_6324
timestamp 1677677812
transform 1 0 3232 0 1 2170
box -8 -3 16 105
use FILL  FILL_6325
timestamp 1677677812
transform 1 0 3240 0 1 2170
box -8 -3 16 105
use FILL  FILL_6326
timestamp 1677677812
transform 1 0 3248 0 1 2170
box -8 -3 16 105
use FILL  FILL_6327
timestamp 1677677812
transform 1 0 3256 0 1 2170
box -8 -3 16 105
use BUFX2  BUFX2_61
timestamp 1677677812
transform 1 0 3264 0 1 2170
box -5 -3 28 105
use FILL  FILL_6328
timestamp 1677677812
transform 1 0 3288 0 1 2170
box -8 -3 16 105
use FILL  FILL_6329
timestamp 1677677812
transform 1 0 3296 0 1 2170
box -8 -3 16 105
use FILL  FILL_6335
timestamp 1677677812
transform 1 0 3304 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_39
timestamp 1677677812
transform -1 0 3344 0 1 2170
box -8 -3 40 105
use FILL  FILL_6336
timestamp 1677677812
transform 1 0 3344 0 1 2170
box -8 -3 16 105
use FILL  FILL_6337
timestamp 1677677812
transform 1 0 3352 0 1 2170
box -8 -3 16 105
use FILL  FILL_6338
timestamp 1677677812
transform 1 0 3360 0 1 2170
box -8 -3 16 105
use FILL  FILL_6343
timestamp 1677677812
transform 1 0 3368 0 1 2170
box -8 -3 16 105
use FILL  FILL_6345
timestamp 1677677812
transform 1 0 3376 0 1 2170
box -8 -3 16 105
use FILL  FILL_6346
timestamp 1677677812
transform 1 0 3384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6347
timestamp 1677677812
transform 1 0 3392 0 1 2170
box -8 -3 16 105
use FILL  FILL_6348
timestamp 1677677812
transform 1 0 3400 0 1 2170
box -8 -3 16 105
use FILL  FILL_6349
timestamp 1677677812
transform 1 0 3408 0 1 2170
box -8 -3 16 105
use FILL  FILL_6350
timestamp 1677677812
transform 1 0 3416 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_403
timestamp 1677677812
transform -1 0 3440 0 1 2170
box -9 -3 26 105
use FILL  FILL_6351
timestamp 1677677812
transform 1 0 3440 0 1 2170
box -8 -3 16 105
use FILL  FILL_6352
timestamp 1677677812
transform 1 0 3448 0 1 2170
box -8 -3 16 105
use FILL  FILL_6353
timestamp 1677677812
transform 1 0 3456 0 1 2170
box -8 -3 16 105
use FILL  FILL_6354
timestamp 1677677812
transform 1 0 3464 0 1 2170
box -8 -3 16 105
use FILL  FILL_6355
timestamp 1677677812
transform 1 0 3472 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_251
timestamp 1677677812
transform 1 0 3480 0 1 2170
box -8 -3 46 105
use FILL  FILL_6357
timestamp 1677677812
transform 1 0 3520 0 1 2170
box -8 -3 16 105
use FILL  FILL_6358
timestamp 1677677812
transform 1 0 3528 0 1 2170
box -8 -3 16 105
use FILL  FILL_6359
timestamp 1677677812
transform 1 0 3536 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_239
timestamp 1677677812
transform 1 0 3544 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_404
timestamp 1677677812
transform -1 0 3600 0 1 2170
box -9 -3 26 105
use FILL  FILL_6363
timestamp 1677677812
transform 1 0 3600 0 1 2170
box -8 -3 16 105
use FILL  FILL_6364
timestamp 1677677812
transform 1 0 3608 0 1 2170
box -8 -3 16 105
use FILL  FILL_6365
timestamp 1677677812
transform 1 0 3616 0 1 2170
box -8 -3 16 105
use FILL  FILL_6371
timestamp 1677677812
transform 1 0 3624 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_241
timestamp 1677677812
transform 1 0 3632 0 1 2170
box -8 -3 46 105
use FILL  FILL_6373
timestamp 1677677812
transform 1 0 3672 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4808
timestamp 1677677812
transform 1 0 3692 0 1 2175
box -3 -3 3 3
use FILL  FILL_6374
timestamp 1677677812
transform 1 0 3680 0 1 2170
box -8 -3 16 105
use FILL  FILL_6375
timestamp 1677677812
transform 1 0 3688 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4809
timestamp 1677677812
transform 1 0 3724 0 1 2175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_358
timestamp 1677677812
transform 1 0 3696 0 1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4810
timestamp 1677677812
transform 1 0 3804 0 1 2175
box -3 -3 3 3
use INVX2  INVX2_405
timestamp 1677677812
transform 1 0 3792 0 1 2170
box -9 -3 26 105
use FILL  FILL_6379
timestamp 1677677812
transform 1 0 3808 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4811
timestamp 1677677812
transform 1 0 3852 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_243
timestamp 1677677812
transform 1 0 3816 0 1 2170
box -8 -3 46 105
use FILL  FILL_6380
timestamp 1677677812
transform 1 0 3856 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4812
timestamp 1677677812
transform 1 0 3892 0 1 2175
box -3 -3 3 3
use AOI22X1  AOI22X1_252
timestamp 1677677812
transform -1 0 3904 0 1 2170
box -8 -3 46 105
use FILL  FILL_6381
timestamp 1677677812
transform 1 0 3904 0 1 2170
box -8 -3 16 105
use FILL  FILL_6382
timestamp 1677677812
transform 1 0 3912 0 1 2170
box -8 -3 16 105
use FILL  FILL_6383
timestamp 1677677812
transform 1 0 3920 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_253
timestamp 1677677812
transform 1 0 3928 0 1 2170
box -8 -3 46 105
use FILL  FILL_6395
timestamp 1677677812
transform 1 0 3968 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4813
timestamp 1677677812
transform 1 0 3988 0 1 2175
box -3 -3 3 3
use FILL  FILL_6396
timestamp 1677677812
transform 1 0 3976 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_407
timestamp 1677677812
transform -1 0 4000 0 1 2170
box -9 -3 26 105
use OAI22X1  OAI22X1_244
timestamp 1677677812
transform 1 0 4000 0 1 2170
box -8 -3 46 105
use FILL  FILL_6397
timestamp 1677677812
transform 1 0 4040 0 1 2170
box -8 -3 16 105
use FILL  FILL_6398
timestamp 1677677812
transform 1 0 4048 0 1 2170
box -8 -3 16 105
use FILL  FILL_6399
timestamp 1677677812
transform 1 0 4056 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_408
timestamp 1677677812
transform -1 0 4080 0 1 2170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_360
timestamp 1677677812
transform -1 0 4176 0 1 2170
box -8 -3 104 105
use FILL  FILL_6400
timestamp 1677677812
transform 1 0 4176 0 1 2170
box -8 -3 16 105
use FILL  FILL_6401
timestamp 1677677812
transform 1 0 4184 0 1 2170
box -8 -3 16 105
use FILL  FILL_6402
timestamp 1677677812
transform 1 0 4192 0 1 2170
box -8 -3 16 105
use FILL  FILL_6403
timestamp 1677677812
transform 1 0 4200 0 1 2170
box -8 -3 16 105
use FILL  FILL_6404
timestamp 1677677812
transform 1 0 4208 0 1 2170
box -8 -3 16 105
use FILL  FILL_6405
timestamp 1677677812
transform 1 0 4216 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_41
timestamp 1677677812
transform -1 0 4256 0 1 2170
box -8 -3 40 105
use FILL  FILL_6406
timestamp 1677677812
transform 1 0 4256 0 1 2170
box -8 -3 16 105
use FILL  FILL_6423
timestamp 1677677812
transform 1 0 4264 0 1 2170
box -8 -3 16 105
use FILL  FILL_6425
timestamp 1677677812
transform 1 0 4272 0 1 2170
box -8 -3 16 105
use FILL  FILL_6427
timestamp 1677677812
transform 1 0 4280 0 1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_42
timestamp 1677677812
transform -1 0 4320 0 1 2170
box -8 -3 40 105
use FILL  FILL_6428
timestamp 1677677812
transform 1 0 4320 0 1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_254
timestamp 1677677812
transform 1 0 4328 0 1 2170
box -8 -3 46 105
use FILL  FILL_6435
timestamp 1677677812
transform 1 0 4368 0 1 2170
box -8 -3 16 105
use FILL  FILL_6436
timestamp 1677677812
transform 1 0 4376 0 1 2170
box -8 -3 16 105
use FILL  FILL_6437
timestamp 1677677812
transform 1 0 4384 0 1 2170
box -8 -3 16 105
use FILL  FILL_6438
timestamp 1677677812
transform 1 0 4392 0 1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4814
timestamp 1677677812
transform 1 0 4436 0 1 2175
box -3 -3 3 3
use OAI22X1  OAI22X1_248
timestamp 1677677812
transform 1 0 4400 0 1 2170
box -8 -3 46 105
use FILL  FILL_6443
timestamp 1677677812
transform 1 0 4440 0 1 2170
box -8 -3 16 105
use FILL  FILL_6444
timestamp 1677677812
transform 1 0 4448 0 1 2170
box -8 -3 16 105
use FILL  FILL_6445
timestamp 1677677812
transform 1 0 4456 0 1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_362
timestamp 1677677812
transform 1 0 4464 0 1 2170
box -8 -3 104 105
use INVX2  INVX2_411
timestamp 1677677812
transform 1 0 4560 0 1 2170
box -9 -3 26 105
use AOI22X1  AOI22X1_255
timestamp 1677677812
transform 1 0 4576 0 1 2170
box -8 -3 46 105
use INVX2  INVX2_412
timestamp 1677677812
transform -1 0 4632 0 1 2170
box -9 -3 26 105
use FILL  FILL_6446
timestamp 1677677812
transform 1 0 4632 0 1 2170
box -8 -3 16 105
use FILL  FILL_6460
timestamp 1677677812
transform 1 0 4640 0 1 2170
box -8 -3 16 105
use FILL  FILL_6462
timestamp 1677677812
transform 1 0 4648 0 1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_250
timestamp 1677677812
transform 1 0 4656 0 1 2170
box -8 -3 46 105
use FILL  FILL_6464
timestamp 1677677812
transform 1 0 4696 0 1 2170
box -8 -3 16 105
use FILL  FILL_6465
timestamp 1677677812
transform 1 0 4704 0 1 2170
box -8 -3 16 105
use FILL  FILL_6466
timestamp 1677677812
transform 1 0 4712 0 1 2170
box -8 -3 16 105
use FILL  FILL_6467
timestamp 1677677812
transform 1 0 4720 0 1 2170
box -8 -3 16 105
use FILL  FILL_6468
timestamp 1677677812
transform 1 0 4728 0 1 2170
box -8 -3 16 105
use FILL  FILL_6469
timestamp 1677677812
transform 1 0 4736 0 1 2170
box -8 -3 16 105
use FILL  FILL_6470
timestamp 1677677812
transform 1 0 4744 0 1 2170
box -8 -3 16 105
use INVX2  INVX2_415
timestamp 1677677812
transform -1 0 4768 0 1 2170
box -9 -3 26 105
use FILL  FILL_6471
timestamp 1677677812
transform 1 0 4768 0 1 2170
box -8 -3 16 105
use FILL  FILL_6472
timestamp 1677677812
transform 1 0 4776 0 1 2170
box -8 -3 16 105
use FILL  FILL_6473
timestamp 1677677812
transform 1 0 4784 0 1 2170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_51
timestamp 1677677812
transform 1 0 4819 0 1 2170
box -10 -3 10 3
use M2_M1  M2_M1_5452
timestamp 1677677812
transform 1 0 108 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5453
timestamp 1677677812
transform 1 0 196 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5366
timestamp 1677677812
transform 1 0 228 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4892
timestamp 1677677812
transform 1 0 252 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5454
timestamp 1677677812
transform 1 0 268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5367
timestamp 1677677812
transform 1 0 292 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4893
timestamp 1677677812
transform 1 0 292 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5455
timestamp 1677677812
transform 1 0 324 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4951
timestamp 1677677812
transform 1 0 364 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5368
timestamp 1677677812
transform 1 0 412 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4851
timestamp 1677677812
transform 1 0 452 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5369
timestamp 1677677812
transform 1 0 436 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5370
timestamp 1677677812
transform 1 0 452 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5371
timestamp 1677677812
transform 1 0 460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5456
timestamp 1677677812
transform 1 0 428 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5457
timestamp 1677677812
transform 1 0 444 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4909
timestamp 1677677812
transform 1 0 428 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4934
timestamp 1677677812
transform 1 0 436 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4946
timestamp 1677677812
transform 1 0 444 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4815
timestamp 1677677812
transform 1 0 516 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4834
timestamp 1677677812
transform 1 0 508 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4816
timestamp 1677677812
transform 1 0 548 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4835
timestamp 1677677812
transform 1 0 556 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4872
timestamp 1677677812
transform 1 0 532 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5372
timestamp 1677677812
transform 1 0 540 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5458
timestamp 1677677812
transform 1 0 532 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5459
timestamp 1677677812
transform 1 0 548 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5460
timestamp 1677677812
transform 1 0 556 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4910
timestamp 1677677812
transform 1 0 524 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4911
timestamp 1677677812
transform 1 0 548 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4947
timestamp 1677677812
transform 1 0 532 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5373
timestamp 1677677812
transform 1 0 572 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4894
timestamp 1677677812
transform 1 0 572 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4817
timestamp 1677677812
transform 1 0 596 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5461
timestamp 1677677812
transform 1 0 596 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4818
timestamp 1677677812
transform 1 0 612 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5374
timestamp 1677677812
transform 1 0 612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5375
timestamp 1677677812
transform 1 0 620 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4895
timestamp 1677677812
transform 1 0 612 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4836
timestamp 1677677812
transform 1 0 636 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4837
timestamp 1677677812
transform 1 0 676 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4852
timestamp 1677677812
transform 1 0 676 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5462
timestamp 1677677812
transform 1 0 676 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5538
timestamp 1677677812
transform 1 0 676 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5376
timestamp 1677677812
transform 1 0 732 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4873
timestamp 1677677812
transform 1 0 740 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5463
timestamp 1677677812
transform 1 0 724 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4896
timestamp 1677677812
transform 1 0 732 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5464
timestamp 1677677812
transform 1 0 788 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4952
timestamp 1677677812
transform 1 0 788 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5377
timestamp 1677677812
transform 1 0 812 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4853
timestamp 1677677812
transform 1 0 852 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5378
timestamp 1677677812
transform 1 0 852 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5379
timestamp 1677677812
transform 1 0 868 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5465
timestamp 1677677812
transform 1 0 844 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5466
timestamp 1677677812
transform 1 0 860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5467
timestamp 1677677812
transform 1 0 932 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4838
timestamp 1677677812
transform 1 0 948 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4854
timestamp 1677677812
transform 1 0 948 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5380
timestamp 1677677812
transform 1 0 948 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4839
timestamp 1677677812
transform 1 0 980 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5468
timestamp 1677677812
transform 1 0 988 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4953
timestamp 1677677812
transform 1 0 988 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5381
timestamp 1677677812
transform 1 0 1012 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5382
timestamp 1677677812
transform 1 0 1036 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4897
timestamp 1677677812
transform 1 0 1060 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5539
timestamp 1677677812
transform 1 0 1060 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5540
timestamp 1677677812
transform 1 0 1068 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5469
timestamp 1677677812
transform 1 0 1092 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4935
timestamp 1677677812
transform 1 0 1100 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4954
timestamp 1677677812
transform 1 0 1092 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5383
timestamp 1677677812
transform 1 0 1124 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4955
timestamp 1677677812
transform 1 0 1132 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5470
timestamp 1677677812
transform 1 0 1180 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4840
timestamp 1677677812
transform 1 0 1212 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4898
timestamp 1677677812
transform 1 0 1236 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4819
timestamp 1677677812
transform 1 0 1284 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4841
timestamp 1677677812
transform 1 0 1276 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4855
timestamp 1677677812
transform 1 0 1260 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4856
timestamp 1677677812
transform 1 0 1284 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5384
timestamp 1677677812
transform 1 0 1260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5385
timestamp 1677677812
transform 1 0 1276 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5386
timestamp 1677677812
transform 1 0 1284 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5471
timestamp 1677677812
transform 1 0 1268 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5472
timestamp 1677677812
transform 1 0 1308 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4820
timestamp 1677677812
transform 1 0 1380 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5541
timestamp 1677677812
transform 1 0 1372 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5387
timestamp 1677677812
transform 1 0 1388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5473
timestamp 1677677812
transform 1 0 1396 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4936
timestamp 1677677812
transform 1 0 1388 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5542
timestamp 1677677812
transform 1 0 1420 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4937
timestamp 1677677812
transform 1 0 1420 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5388
timestamp 1677677812
transform 1 0 1436 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4956
timestamp 1677677812
transform 1 0 1452 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5474
timestamp 1677677812
transform 1 0 1500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5389
timestamp 1677677812
transform 1 0 1516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5390
timestamp 1677677812
transform 1 0 1532 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4821
timestamp 1677677812
transform 1 0 1580 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5391
timestamp 1677677812
transform 1 0 1556 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5475
timestamp 1677677812
transform 1 0 1588 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4957
timestamp 1677677812
transform 1 0 1556 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4822
timestamp 1677677812
transform 1 0 1676 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5476
timestamp 1677677812
transform 1 0 1676 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5477
timestamp 1677677812
transform 1 0 1684 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4842
timestamp 1677677812
transform 1 0 1732 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4857
timestamp 1677677812
transform 1 0 1724 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5392
timestamp 1677677812
transform 1 0 1724 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5478
timestamp 1677677812
transform 1 0 1716 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5393
timestamp 1677677812
transform 1 0 1764 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5479
timestamp 1677677812
transform 1 0 1812 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4948
timestamp 1677677812
transform 1 0 1860 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4874
timestamp 1677677812
transform 1 0 1900 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5480
timestamp 1677677812
transform 1 0 1900 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5394
timestamp 1677677812
transform 1 0 1916 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5395
timestamp 1677677812
transform 1 0 1932 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4875
timestamp 1677677812
transform 1 0 1940 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5396
timestamp 1677677812
transform 1 0 1948 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5481
timestamp 1677677812
transform 1 0 1924 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5482
timestamp 1677677812
transform 1 0 1940 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4899
timestamp 1677677812
transform 1 0 1948 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4912
timestamp 1677677812
transform 1 0 1924 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4938
timestamp 1677677812
transform 1 0 1932 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5397
timestamp 1677677812
transform 1 0 2036 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4858
timestamp 1677677812
transform 1 0 2060 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5398
timestamp 1677677812
transform 1 0 2060 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5483
timestamp 1677677812
transform 1 0 2052 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4900
timestamp 1677677812
transform 1 0 2060 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5484
timestamp 1677677812
transform 1 0 2068 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4913
timestamp 1677677812
transform 1 0 2044 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4949
timestamp 1677677812
transform 1 0 2052 0 1 2095
box -3 -3 3 3
use M2_M1  M2_M1_5399
timestamp 1677677812
transform 1 0 2084 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4901
timestamp 1677677812
transform 1 0 2148 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4823
timestamp 1677677812
transform 1 0 2164 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5400
timestamp 1677677812
transform 1 0 2164 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5401
timestamp 1677677812
transform 1 0 2180 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5485
timestamp 1677677812
transform 1 0 2188 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4950
timestamp 1677677812
transform 1 0 2188 0 1 2095
box -3 -3 3 3
use M3_M2  M3_M2_4902
timestamp 1677677812
transform 1 0 2204 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5402
timestamp 1677677812
transform 1 0 2252 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4824
timestamp 1677677812
transform 1 0 2292 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4825
timestamp 1677677812
transform 1 0 2364 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5403
timestamp 1677677812
transform 1 0 2284 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5486
timestamp 1677677812
transform 1 0 2308 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5487
timestamp 1677677812
transform 1 0 2364 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4914
timestamp 1677677812
transform 1 0 2364 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5488
timestamp 1677677812
transform 1 0 2388 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4915
timestamp 1677677812
transform 1 0 2388 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4903
timestamp 1677677812
transform 1 0 2412 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4876
timestamp 1677677812
transform 1 0 2436 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5404
timestamp 1677677812
transform 1 0 2444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5489
timestamp 1677677812
transform 1 0 2436 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5490
timestamp 1677677812
transform 1 0 2460 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4916
timestamp 1677677812
transform 1 0 2468 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4877
timestamp 1677677812
transform 1 0 2508 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5405
timestamp 1677677812
transform 1 0 2516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5491
timestamp 1677677812
transform 1 0 2508 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4917
timestamp 1677677812
transform 1 0 2508 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5406
timestamp 1677677812
transform 1 0 2564 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4918
timestamp 1677677812
transform 1 0 2564 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5407
timestamp 1677677812
transform 1 0 2580 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4904
timestamp 1677677812
transform 1 0 2580 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4958
timestamp 1677677812
transform 1 0 2572 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4878
timestamp 1677677812
transform 1 0 2620 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5492
timestamp 1677677812
transform 1 0 2620 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4859
timestamp 1677677812
transform 1 0 2660 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5364
timestamp 1677677812
transform 1 0 2668 0 1 2145
box -2 -2 2 2
use M2_M1  M2_M1_5408
timestamp 1677677812
transform 1 0 2636 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5493
timestamp 1677677812
transform 1 0 2644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5494
timestamp 1677677812
transform 1 0 2660 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4919
timestamp 1677677812
transform 1 0 2644 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4959
timestamp 1677677812
transform 1 0 2636 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4879
timestamp 1677677812
transform 1 0 2676 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4880
timestamp 1677677812
transform 1 0 2716 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5409
timestamp 1677677812
transform 1 0 2732 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5365
timestamp 1677677812
transform 1 0 2772 0 1 2145
box -2 -2 2 2
use M3_M2  M3_M2_4939
timestamp 1677677812
transform 1 0 2772 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5495
timestamp 1677677812
transform 1 0 2828 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4826
timestamp 1677677812
transform 1 0 2844 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5410
timestamp 1677677812
transform 1 0 2844 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5496
timestamp 1677677812
transform 1 0 2860 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5411
timestamp 1677677812
transform 1 0 2892 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5412
timestamp 1677677812
transform 1 0 2900 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4905
timestamp 1677677812
transform 1 0 2892 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4881
timestamp 1677677812
transform 1 0 2908 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5497
timestamp 1677677812
transform 1 0 2908 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5498
timestamp 1677677812
transform 1 0 2956 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4960
timestamp 1677677812
transform 1 0 2956 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5413
timestamp 1677677812
transform 1 0 2972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5414
timestamp 1677677812
transform 1 0 2988 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4882
timestamp 1677677812
transform 1 0 2996 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4860
timestamp 1677677812
transform 1 0 3020 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5415
timestamp 1677677812
transform 1 0 3020 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5499
timestamp 1677677812
transform 1 0 2980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5500
timestamp 1677677812
transform 1 0 3004 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5501
timestamp 1677677812
transform 1 0 3012 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4920
timestamp 1677677812
transform 1 0 2972 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4921
timestamp 1677677812
transform 1 0 2988 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4922
timestamp 1677677812
transform 1 0 3004 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4940
timestamp 1677677812
transform 1 0 3004 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4843
timestamp 1677677812
transform 1 0 3108 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4883
timestamp 1677677812
transform 1 0 3060 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5416
timestamp 1677677812
transform 1 0 3108 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5502
timestamp 1677677812
transform 1 0 3060 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4923
timestamp 1677677812
transform 1 0 3036 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4941
timestamp 1677677812
transform 1 0 3028 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4844
timestamp 1677677812
transform 1 0 3132 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5417
timestamp 1677677812
transform 1 0 3132 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5503
timestamp 1677677812
transform 1 0 3172 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5504
timestamp 1677677812
transform 1 0 3212 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5505
timestamp 1677677812
transform 1 0 3220 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4924
timestamp 1677677812
transform 1 0 3132 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4925
timestamp 1677677812
transform 1 0 3172 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4884
timestamp 1677677812
transform 1 0 3236 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4942
timestamp 1677677812
transform 1 0 3228 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5418
timestamp 1677677812
transform 1 0 3260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5543
timestamp 1677677812
transform 1 0 3260 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4943
timestamp 1677677812
transform 1 0 3260 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4885
timestamp 1677677812
transform 1 0 3300 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5544
timestamp 1677677812
transform 1 0 3292 0 1 2115
box -2 -2 2 2
use M2_M1  M2_M1_5546
timestamp 1677677812
transform 1 0 3276 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4827
timestamp 1677677812
transform 1 0 3324 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4886
timestamp 1677677812
transform 1 0 3324 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4906
timestamp 1677677812
transform 1 0 3340 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5506
timestamp 1677677812
transform 1 0 3348 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5547
timestamp 1677677812
transform 1 0 3340 0 1 2105
box -2 -2 2 2
use M3_M2  M3_M2_4887
timestamp 1677677812
transform 1 0 3364 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4907
timestamp 1677677812
transform 1 0 3372 0 1 2125
box -3 -3 3 3
use M2_M1  M2_M1_5545
timestamp 1677677812
transform 1 0 3372 0 1 2115
box -2 -2 2 2
use M3_M2  M3_M2_4961
timestamp 1677677812
transform 1 0 3372 0 1 2085
box -3 -3 3 3
use M2_M1  M2_M1_5419
timestamp 1677677812
transform 1 0 3388 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4845
timestamp 1677677812
transform 1 0 3476 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5420
timestamp 1677677812
transform 1 0 3476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5507
timestamp 1677677812
transform 1 0 3412 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5508
timestamp 1677677812
transform 1 0 3468 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5509
timestamp 1677677812
transform 1 0 3476 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5421
timestamp 1677677812
transform 1 0 3516 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5422
timestamp 1677677812
transform 1 0 3532 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5510
timestamp 1677677812
transform 1 0 3524 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4962
timestamp 1677677812
transform 1 0 3532 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4861
timestamp 1677677812
transform 1 0 3548 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4862
timestamp 1677677812
transform 1 0 3564 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4846
timestamp 1677677812
transform 1 0 3612 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4863
timestamp 1677677812
transform 1 0 3596 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5423
timestamp 1677677812
transform 1 0 3572 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5424
timestamp 1677677812
transform 1 0 3580 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5425
timestamp 1677677812
transform 1 0 3596 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5426
timestamp 1677677812
transform 1 0 3612 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5427
timestamp 1677677812
transform 1 0 3620 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5511
timestamp 1677677812
transform 1 0 3588 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4926
timestamp 1677677812
transform 1 0 3580 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5512
timestamp 1677677812
transform 1 0 3644 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5428
timestamp 1677677812
transform 1 0 3668 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5429
timestamp 1677677812
transform 1 0 3684 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5430
timestamp 1677677812
transform 1 0 3692 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5513
timestamp 1677677812
transform 1 0 3676 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4927
timestamp 1677677812
transform 1 0 3684 0 1 2115
box -3 -3 3 3
use M2_M1  M2_M1_5514
timestamp 1677677812
transform 1 0 3724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5515
timestamp 1677677812
transform 1 0 3804 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4828
timestamp 1677677812
transform 1 0 3828 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4829
timestamp 1677677812
transform 1 0 3852 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4830
timestamp 1677677812
transform 1 0 3900 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5431
timestamp 1677677812
transform 1 0 3820 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5516
timestamp 1677677812
transform 1 0 3844 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4908
timestamp 1677677812
transform 1 0 3884 0 1 2125
box -3 -3 3 3
use M3_M2  M3_M2_4847
timestamp 1677677812
transform 1 0 3924 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5432
timestamp 1677677812
transform 1 0 3924 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5517
timestamp 1677677812
transform 1 0 3916 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5518
timestamp 1677677812
transform 1 0 3932 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4963
timestamp 1677677812
transform 1 0 3948 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4831
timestamp 1677677812
transform 1 0 3996 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5433
timestamp 1677677812
transform 1 0 3972 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5434
timestamp 1677677812
transform 1 0 3988 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5519
timestamp 1677677812
transform 1 0 3980 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5520
timestamp 1677677812
transform 1 0 3996 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4964
timestamp 1677677812
transform 1 0 3980 0 1 2085
box -3 -3 3 3
use M3_M2  M3_M2_4864
timestamp 1677677812
transform 1 0 4004 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5521
timestamp 1677677812
transform 1 0 4012 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4865
timestamp 1677677812
transform 1 0 4036 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4866
timestamp 1677677812
transform 1 0 4068 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5435
timestamp 1677677812
transform 1 0 4028 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5436
timestamp 1677677812
transform 1 0 4036 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5437
timestamp 1677677812
transform 1 0 4052 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4888
timestamp 1677677812
transform 1 0 4060 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5438
timestamp 1677677812
transform 1 0 4068 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5522
timestamp 1677677812
transform 1 0 4044 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5523
timestamp 1677677812
transform 1 0 4060 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4928
timestamp 1677677812
transform 1 0 4060 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4944
timestamp 1677677812
transform 1 0 4044 0 1 2105
box -3 -3 3 3
use M2_M1  M2_M1_5439
timestamp 1677677812
transform 1 0 4156 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4889
timestamp 1677677812
transform 1 0 4180 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5524
timestamp 1677677812
transform 1 0 4180 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4867
timestamp 1677677812
transform 1 0 4260 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5440
timestamp 1677677812
transform 1 0 4260 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5525
timestamp 1677677812
transform 1 0 4252 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4929
timestamp 1677677812
transform 1 0 4252 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4930
timestamp 1677677812
transform 1 0 4332 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4848
timestamp 1677677812
transform 1 0 4388 0 1 2155
box -3 -3 3 3
use M2_M1  M2_M1_5441
timestamp 1677677812
transform 1 0 4372 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5442
timestamp 1677677812
transform 1 0 4388 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5443
timestamp 1677677812
transform 1 0 4396 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5526
timestamp 1677677812
transform 1 0 4364 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5527
timestamp 1677677812
transform 1 0 4380 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4931
timestamp 1677677812
transform 1 0 4364 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4945
timestamp 1677677812
transform 1 0 4380 0 1 2105
box -3 -3 3 3
use M3_M2  M3_M2_4868
timestamp 1677677812
transform 1 0 4444 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5444
timestamp 1677677812
transform 1 0 4444 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5445
timestamp 1677677812
transform 1 0 4460 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5528
timestamp 1677677812
transform 1 0 4460 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4932
timestamp 1677677812
transform 1 0 4460 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4869
timestamp 1677677812
transform 1 0 4476 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5446
timestamp 1677677812
transform 1 0 4476 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5529
timestamp 1677677812
transform 1 0 4484 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5530
timestamp 1677677812
transform 1 0 4500 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5447
timestamp 1677677812
transform 1 0 4524 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5531
timestamp 1677677812
transform 1 0 4524 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5532
timestamp 1677677812
transform 1 0 4540 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5533
timestamp 1677677812
transform 1 0 4556 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4933
timestamp 1677677812
transform 1 0 4540 0 1 2115
box -3 -3 3 3
use M3_M2  M3_M2_4870
timestamp 1677677812
transform 1 0 4588 0 1 2145
box -3 -3 3 3
use M3_M2  M3_M2_4849
timestamp 1677677812
transform 1 0 4620 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4871
timestamp 1677677812
transform 1 0 4628 0 1 2145
box -3 -3 3 3
use M2_M1  M2_M1_5448
timestamp 1677677812
transform 1 0 4588 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5449
timestamp 1677677812
transform 1 0 4604 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5450
timestamp 1677677812
transform 1 0 4620 0 1 2135
box -2 -2 2 2
use M2_M1  M2_M1_5534
timestamp 1677677812
transform 1 0 4596 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5535
timestamp 1677677812
transform 1 0 4636 0 1 2125
box -2 -2 2 2
use M3_M2  M3_M2_4850
timestamp 1677677812
transform 1 0 4652 0 1 2155
box -3 -3 3 3
use M3_M2  M3_M2_4890
timestamp 1677677812
transform 1 0 4676 0 1 2135
box -3 -3 3 3
use M3_M2  M3_M2_4832
timestamp 1677677812
transform 1 0 4700 0 1 2165
box -3 -3 3 3
use M3_M2  M3_M2_4833
timestamp 1677677812
transform 1 0 4756 0 1 2165
box -3 -3 3 3
use M2_M1  M2_M1_5451
timestamp 1677677812
transform 1 0 4700 0 1 2135
box -2 -2 2 2
use M3_M2  M3_M2_4891
timestamp 1677677812
transform 1 0 4724 0 1 2135
box -3 -3 3 3
use M2_M1  M2_M1_5536
timestamp 1677677812
transform 1 0 4724 0 1 2125
box -2 -2 2 2
use M2_M1  M2_M1_5537
timestamp 1677677812
transform 1 0 4788 0 1 2125
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_52
timestamp 1677677812
transform 1 0 24 0 1 2070
box -10 -3 10 3
use FILL  FILL_5894
timestamp 1677677812
transform 1 0 72 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5895
timestamp 1677677812
transform 1 0 80 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5896
timestamp 1677677812
transform 1 0 88 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5897
timestamp 1677677812
transform 1 0 96 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_388
timestamp 1677677812
transform -1 0 120 0 -1 2170
box -9 -3 26 105
use FILL  FILL_5898
timestamp 1677677812
transform 1 0 120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5899
timestamp 1677677812
transform 1 0 128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5900
timestamp 1677677812
transform 1 0 136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5901
timestamp 1677677812
transform 1 0 144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5902
timestamp 1677677812
transform 1 0 152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5903
timestamp 1677677812
transform 1 0 160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5904
timestamp 1677677812
transform 1 0 168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5906
timestamp 1677677812
transform 1 0 176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5907
timestamp 1677677812
transform 1 0 184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5908
timestamp 1677677812
transform 1 0 192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5910
timestamp 1677677812
transform 1 0 200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5919
timestamp 1677677812
transform 1 0 208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5920
timestamp 1677677812
transform 1 0 216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5921
timestamp 1677677812
transform 1 0 224 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_391
timestamp 1677677812
transform -1 0 248 0 -1 2170
box -9 -3 26 105
use FILL  FILL_5922
timestamp 1677677812
transform 1 0 248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5923
timestamp 1677677812
transform 1 0 256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5924
timestamp 1677677812
transform 1 0 264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5925
timestamp 1677677812
transform 1 0 272 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_347
timestamp 1677677812
transform 1 0 280 0 -1 2170
box -8 -3 104 105
use FILL  FILL_5926
timestamp 1677677812
transform 1 0 376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5932
timestamp 1677677812
transform 1 0 384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5933
timestamp 1677677812
transform 1 0 392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5934
timestamp 1677677812
transform 1 0 400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5935
timestamp 1677677812
transform 1 0 408 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_228
timestamp 1677677812
transform 1 0 416 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5936
timestamp 1677677812
transform 1 0 456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5937
timestamp 1677677812
transform 1 0 464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5938
timestamp 1677677812
transform 1 0 472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5939
timestamp 1677677812
transform 1 0 480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5940
timestamp 1677677812
transform 1 0 488 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5941
timestamp 1677677812
transform 1 0 496 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5943
timestamp 1677677812
transform 1 0 504 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5950
timestamp 1677677812
transform 1 0 512 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_229
timestamp 1677677812
transform -1 0 560 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5951
timestamp 1677677812
transform 1 0 560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5952
timestamp 1677677812
transform 1 0 568 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_11
timestamp 1677677812
transform -1 0 608 0 -1 2170
box -8 -3 40 105
use FILL  FILL_5953
timestamp 1677677812
transform 1 0 608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5954
timestamp 1677677812
transform 1 0 616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5955
timestamp 1677677812
transform 1 0 624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5956
timestamp 1677677812
transform 1 0 632 0 -1 2170
box -8 -3 16 105
use BUFX2  BUFX2_58
timestamp 1677677812
transform -1 0 664 0 -1 2170
box -5 -3 28 105
use FILL  FILL_5957
timestamp 1677677812
transform 1 0 664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5959
timestamp 1677677812
transform 1 0 672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5961
timestamp 1677677812
transform 1 0 680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5967
timestamp 1677677812
transform 1 0 688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5968
timestamp 1677677812
transform 1 0 696 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_12
timestamp 1677677812
transform -1 0 736 0 -1 2170
box -8 -3 40 105
use FILL  FILL_5969
timestamp 1677677812
transform 1 0 736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5971
timestamp 1677677812
transform 1 0 744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5973
timestamp 1677677812
transform 1 0 752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5975
timestamp 1677677812
transform 1 0 760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5978
timestamp 1677677812
transform 1 0 768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5979
timestamp 1677677812
transform 1 0 776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5980
timestamp 1677677812
transform 1 0 784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5981
timestamp 1677677812
transform 1 0 792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5982
timestamp 1677677812
transform 1 0 800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5983
timestamp 1677677812
transform 1 0 808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5984
timestamp 1677677812
transform 1 0 816 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_241
timestamp 1677677812
transform 1 0 824 0 -1 2170
box -8 -3 46 105
use FILL  FILL_5991
timestamp 1677677812
transform 1 0 864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5996
timestamp 1677677812
transform 1 0 872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5997
timestamp 1677677812
transform 1 0 880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5998
timestamp 1677677812
transform 1 0 888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_5999
timestamp 1677677812
transform 1 0 896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6000
timestamp 1677677812
transform 1 0 904 0 -1 2170
box -8 -3 16 105
use BUFX2  BUFX2_59
timestamp 1677677812
transform -1 0 936 0 -1 2170
box -5 -3 28 105
use FILL  FILL_6001
timestamp 1677677812
transform 1 0 936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6003
timestamp 1677677812
transform 1 0 944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6005
timestamp 1677677812
transform 1 0 952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6007
timestamp 1677677812
transform 1 0 960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6009
timestamp 1677677812
transform 1 0 968 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_117
timestamp 1677677812
transform 1 0 976 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6012
timestamp 1677677812
transform 1 0 1008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6013
timestamp 1677677812
transform 1 0 1016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6014
timestamp 1677677812
transform 1 0 1024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6016
timestamp 1677677812
transform 1 0 1032 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6018
timestamp 1677677812
transform 1 0 1040 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6020
timestamp 1677677812
transform 1 0 1048 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6022
timestamp 1677677812
transform 1 0 1056 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6029
timestamp 1677677812
transform 1 0 1064 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_118
timestamp 1677677812
transform -1 0 1104 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6030
timestamp 1677677812
transform 1 0 1104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6032
timestamp 1677677812
transform 1 0 1112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6034
timestamp 1677677812
transform 1 0 1120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6036
timestamp 1677677812
transform 1 0 1128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6038
timestamp 1677677812
transform 1 0 1136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6040
timestamp 1677677812
transform 1 0 1144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6042
timestamp 1677677812
transform 1 0 1152 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6044
timestamp 1677677812
transform 1 0 1160 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6047
timestamp 1677677812
transform 1 0 1168 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6048
timestamp 1677677812
transform 1 0 1176 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6049
timestamp 1677677812
transform 1 0 1184 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6050
timestamp 1677677812
transform 1 0 1192 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6051
timestamp 1677677812
transform 1 0 1200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6052
timestamp 1677677812
transform 1 0 1208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6053
timestamp 1677677812
transform 1 0 1216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6055
timestamp 1677677812
transform 1 0 1224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6057
timestamp 1677677812
transform 1 0 1232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6066
timestamp 1677677812
transform 1 0 1240 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_245
timestamp 1677677812
transform -1 0 1288 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6067
timestamp 1677677812
transform 1 0 1288 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4965
timestamp 1677677812
transform 1 0 1308 0 1 2075
box -3 -3 3 3
use FILL  FILL_6068
timestamp 1677677812
transform 1 0 1296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6069
timestamp 1677677812
transform 1 0 1304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6070
timestamp 1677677812
transform 1 0 1312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6071
timestamp 1677677812
transform 1 0 1320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6072
timestamp 1677677812
transform 1 0 1328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6074
timestamp 1677677812
transform 1 0 1336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6076
timestamp 1677677812
transform 1 0 1344 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6078
timestamp 1677677812
transform 1 0 1352 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6080
timestamp 1677677812
transform 1 0 1360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6082
timestamp 1677677812
transform 1 0 1368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6084
timestamp 1677677812
transform 1 0 1376 0 -1 2170
box -8 -3 16 105
use OAI21X1  OAI21X1_121
timestamp 1677677812
transform 1 0 1384 0 -1 2170
box -8 -3 34 105
use FILL  FILL_6090
timestamp 1677677812
transform 1 0 1416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6091
timestamp 1677677812
transform 1 0 1424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6092
timestamp 1677677812
transform 1 0 1432 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6093
timestamp 1677677812
transform 1 0 1440 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6094
timestamp 1677677812
transform 1 0 1448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6096
timestamp 1677677812
transform 1 0 1456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6098
timestamp 1677677812
transform 1 0 1464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6100
timestamp 1677677812
transform 1 0 1472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6102
timestamp 1677677812
transform 1 0 1480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6104
timestamp 1677677812
transform 1 0 1488 0 -1 2170
box -8 -3 16 105
use BUFX2  BUFX2_60
timestamp 1677677812
transform 1 0 1496 0 -1 2170
box -5 -3 28 105
use FILL  FILL_6107
timestamp 1677677812
transform 1 0 1520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6109
timestamp 1677677812
transform 1 0 1528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6111
timestamp 1677677812
transform 1 0 1536 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_349
timestamp 1677677812
transform 1 0 1544 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6120
timestamp 1677677812
transform 1 0 1640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6122
timestamp 1677677812
transform 1 0 1648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6128
timestamp 1677677812
transform 1 0 1656 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_395
timestamp 1677677812
transform 1 0 1664 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6129
timestamp 1677677812
transform 1 0 1680 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4966
timestamp 1677677812
transform 1 0 1700 0 1 2075
box -3 -3 3 3
use FILL  FILL_6130
timestamp 1677677812
transform 1 0 1688 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_13
timestamp 1677677812
transform -1 0 1728 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6131
timestamp 1677677812
transform 1 0 1728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6135
timestamp 1677677812
transform 1 0 1736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6136
timestamp 1677677812
transform 1 0 1744 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_351
timestamp 1677677812
transform 1 0 1752 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6137
timestamp 1677677812
transform 1 0 1848 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6139
timestamp 1677677812
transform 1 0 1856 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6142
timestamp 1677677812
transform 1 0 1864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6143
timestamp 1677677812
transform 1 0 1872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6144
timestamp 1677677812
transform 1 0 1880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6145
timestamp 1677677812
transform 1 0 1888 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6147
timestamp 1677677812
transform 1 0 1896 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6153
timestamp 1677677812
transform 1 0 1904 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_232
timestamp 1677677812
transform -1 0 1952 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6154
timestamp 1677677812
transform 1 0 1952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6155
timestamp 1677677812
transform 1 0 1960 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6156
timestamp 1677677812
transform 1 0 1968 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6157
timestamp 1677677812
transform 1 0 1976 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6159
timestamp 1677677812
transform 1 0 1984 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6162
timestamp 1677677812
transform 1 0 1992 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6163
timestamp 1677677812
transform 1 0 2000 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6164
timestamp 1677677812
transform 1 0 2008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6165
timestamp 1677677812
transform 1 0 2016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6166
timestamp 1677677812
transform 1 0 2024 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6167
timestamp 1677677812
transform 1 0 2032 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_233
timestamp 1677677812
transform -1 0 2080 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6168
timestamp 1677677812
transform 1 0 2080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6169
timestamp 1677677812
transform 1 0 2088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6170
timestamp 1677677812
transform 1 0 2096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6171
timestamp 1677677812
transform 1 0 2104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6172
timestamp 1677677812
transform 1 0 2112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6174
timestamp 1677677812
transform 1 0 2120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6176
timestamp 1677677812
transform 1 0 2128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6178
timestamp 1677677812
transform 1 0 2136 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6180
timestamp 1677677812
transform 1 0 2144 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6182
timestamp 1677677812
transform 1 0 2152 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_234
timestamp 1677677812
transform 1 0 2160 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6185
timestamp 1677677812
transform 1 0 2200 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6186
timestamp 1677677812
transform 1 0 2208 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6188
timestamp 1677677812
transform 1 0 2216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6190
timestamp 1677677812
transform 1 0 2224 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6192
timestamp 1677677812
transform 1 0 2232 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6194
timestamp 1677677812
transform 1 0 2240 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6196
timestamp 1677677812
transform 1 0 2248 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6198
timestamp 1677677812
transform 1 0 2256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6200
timestamp 1677677812
transform 1 0 2264 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_353
timestamp 1677677812
transform 1 0 2272 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6207
timestamp 1677677812
transform 1 0 2368 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6209
timestamp 1677677812
transform 1 0 2376 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6211
timestamp 1677677812
transform 1 0 2384 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6213
timestamp 1677677812
transform 1 0 2392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6215
timestamp 1677677812
transform 1 0 2400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6220
timestamp 1677677812
transform 1 0 2408 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_14
timestamp 1677677812
transform -1 0 2448 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6221
timestamp 1677677812
transform 1 0 2448 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6223
timestamp 1677677812
transform 1 0 2456 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6225
timestamp 1677677812
transform 1 0 2464 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6227
timestamp 1677677812
transform 1 0 2472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6234
timestamp 1677677812
transform 1 0 2480 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_15
timestamp 1677677812
transform -1 0 2520 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6235
timestamp 1677677812
transform 1 0 2520 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6237
timestamp 1677677812
transform 1 0 2528 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6239
timestamp 1677677812
transform 1 0 2536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6241
timestamp 1677677812
transform 1 0 2544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6243
timestamp 1677677812
transform 1 0 2552 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_400
timestamp 1677677812
transform 1 0 2560 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6245
timestamp 1677677812
transform 1 0 2576 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6246
timestamp 1677677812
transform 1 0 2584 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6247
timestamp 1677677812
transform 1 0 2592 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6248
timestamp 1677677812
transform 1 0 2600 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6250
timestamp 1677677812
transform 1 0 2608 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6252
timestamp 1677677812
transform 1 0 2616 0 -1 2170
box -8 -3 16 105
use AOI22X1  AOI22X1_250
timestamp 1677677812
transform 1 0 2624 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6256
timestamp 1677677812
transform 1 0 2664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6257
timestamp 1677677812
transform 1 0 2672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6258
timestamp 1677677812
transform 1 0 2680 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6259
timestamp 1677677812
transform 1 0 2688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6260
timestamp 1677677812
transform 1 0 2696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6261
timestamp 1677677812
transform 1 0 2704 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6262
timestamp 1677677812
transform 1 0 2712 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6263
timestamp 1677677812
transform 1 0 2720 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6264
timestamp 1677677812
transform 1 0 2728 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6265
timestamp 1677677812
transform 1 0 2736 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6267
timestamp 1677677812
transform 1 0 2744 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_58
timestamp 1677677812
transform 1 0 2752 0 -1 2170
box -8 -3 32 105
use FILL  FILL_6272
timestamp 1677677812
transform 1 0 2776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6274
timestamp 1677677812
transform 1 0 2784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6276
timestamp 1677677812
transform 1 0 2792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6277
timestamp 1677677812
transform 1 0 2800 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6278
timestamp 1677677812
transform 1 0 2808 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6279
timestamp 1677677812
transform 1 0 2816 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6280
timestamp 1677677812
transform 1 0 2824 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6282
timestamp 1677677812
transform 1 0 2832 0 -1 2170
box -8 -3 16 105
use NOR2X1  NOR2X1_59
timestamp 1677677812
transform 1 0 2840 0 -1 2170
box -8 -3 32 105
use FILL  FILL_6288
timestamp 1677677812
transform 1 0 2864 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6289
timestamp 1677677812
transform 1 0 2872 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6290
timestamp 1677677812
transform 1 0 2880 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6291
timestamp 1677677812
transform 1 0 2888 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_16
timestamp 1677677812
transform 1 0 2896 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6296
timestamp 1677677812
transform 1 0 2928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6297
timestamp 1677677812
transform 1 0 2936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6298
timestamp 1677677812
transform 1 0 2944 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6299
timestamp 1677677812
transform 1 0 2952 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6307
timestamp 1677677812
transform 1 0 2960 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_235
timestamp 1677677812
transform -1 0 3008 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6308
timestamp 1677677812
transform 1 0 3008 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6330
timestamp 1677677812
transform 1 0 3016 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_355
timestamp 1677677812
transform -1 0 3120 0 -1 2170
box -8 -3 104 105
use M3_M2  M3_M2_4967
timestamp 1677677812
transform 1 0 3220 0 1 2075
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_356
timestamp 1677677812
transform 1 0 3120 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6331
timestamp 1677677812
transform 1 0 3216 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6332
timestamp 1677677812
transform 1 0 3224 0 -1 2170
box -8 -3 16 105
use BUFX2  BUFX2_62
timestamp 1677677812
transform 1 0 3232 0 -1 2170
box -5 -3 28 105
use FILL  FILL_6333
timestamp 1677677812
transform 1 0 3256 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_38
timestamp 1677677812
transform -1 0 3296 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6334
timestamp 1677677812
transform 1 0 3296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6339
timestamp 1677677812
transform 1 0 3304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6340
timestamp 1677677812
transform 1 0 3312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6341
timestamp 1677677812
transform 1 0 3320 0 -1 2170
box -8 -3 16 105
use NAND3X1  NAND3X1_40
timestamp 1677677812
transform -1 0 3360 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6342
timestamp 1677677812
transform 1 0 3360 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6344
timestamp 1677677812
transform 1 0 3368 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_357
timestamp 1677677812
transform 1 0 3376 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6356
timestamp 1677677812
transform 1 0 3472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6360
timestamp 1677677812
transform 1 0 3480 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6361
timestamp 1677677812
transform 1 0 3488 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_238
timestamp 1677677812
transform 1 0 3496 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6362
timestamp 1677677812
transform 1 0 3536 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6366
timestamp 1677677812
transform 1 0 3544 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6367
timestamp 1677677812
transform 1 0 3552 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6368
timestamp 1677677812
transform 1 0 3560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6369
timestamp 1677677812
transform 1 0 3568 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_240
timestamp 1677677812
transform -1 0 3616 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6370
timestamp 1677677812
transform 1 0 3616 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6372
timestamp 1677677812
transform 1 0 3624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6376
timestamp 1677677812
transform 1 0 3632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6377
timestamp 1677677812
transform 1 0 3640 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_242
timestamp 1677677812
transform 1 0 3648 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6378
timestamp 1677677812
transform 1 0 3688 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6384
timestamp 1677677812
transform 1 0 3696 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6385
timestamp 1677677812
transform 1 0 3704 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_17
timestamp 1677677812
transform 1 0 3712 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6386
timestamp 1677677812
transform 1 0 3744 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6387
timestamp 1677677812
transform 1 0 3752 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6388
timestamp 1677677812
transform 1 0 3760 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6389
timestamp 1677677812
transform 1 0 3768 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6390
timestamp 1677677812
transform 1 0 3776 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6391
timestamp 1677677812
transform 1 0 3784 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6392
timestamp 1677677812
transform 1 0 3792 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6393
timestamp 1677677812
transform 1 0 3800 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_359
timestamp 1677677812
transform 1 0 3808 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_406
timestamp 1677677812
transform 1 0 3904 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6394
timestamp 1677677812
transform 1 0 3920 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6407
timestamp 1677677812
transform 1 0 3928 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6408
timestamp 1677677812
transform 1 0 3936 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6409
timestamp 1677677812
transform 1 0 3944 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_245
timestamp 1677677812
transform 1 0 3952 0 -1 2170
box -8 -3 46 105
use INVX2  INVX2_409
timestamp 1677677812
transform -1 0 4008 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6410
timestamp 1677677812
transform 1 0 4008 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4968
timestamp 1677677812
transform 1 0 4028 0 1 2075
box -3 -3 3 3
use FILL  FILL_6411
timestamp 1677677812
transform 1 0 4016 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6412
timestamp 1677677812
transform 1 0 4024 0 -1 2170
box -8 -3 16 105
use M3_M2  M3_M2_4969
timestamp 1677677812
transform 1 0 4044 0 1 2075
box -3 -3 3 3
use OAI22X1  OAI22X1_246
timestamp 1677677812
transform 1 0 4032 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6413
timestamp 1677677812
transform 1 0 4072 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6414
timestamp 1677677812
transform 1 0 4080 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6415
timestamp 1677677812
transform 1 0 4088 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6416
timestamp 1677677812
transform 1 0 4096 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6417
timestamp 1677677812
transform 1 0 4104 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6418
timestamp 1677677812
transform 1 0 4112 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6419
timestamp 1677677812
transform 1 0 4120 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6420
timestamp 1677677812
transform 1 0 4128 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6421
timestamp 1677677812
transform 1 0 4136 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_361
timestamp 1677677812
transform 1 0 4144 0 -1 2170
box -8 -3 104 105
use INVX2  INVX2_410
timestamp 1677677812
transform 1 0 4240 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6422
timestamp 1677677812
transform 1 0 4256 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6424
timestamp 1677677812
transform 1 0 4264 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6426
timestamp 1677677812
transform 1 0 4272 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6429
timestamp 1677677812
transform 1 0 4280 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6430
timestamp 1677677812
transform 1 0 4288 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6431
timestamp 1677677812
transform 1 0 4296 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6432
timestamp 1677677812
transform 1 0 4304 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6433
timestamp 1677677812
transform 1 0 4312 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6434
timestamp 1677677812
transform 1 0 4320 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6439
timestamp 1677677812
transform 1 0 4328 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6440
timestamp 1677677812
transform 1 0 4336 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6441
timestamp 1677677812
transform 1 0 4344 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_247
timestamp 1677677812
transform -1 0 4392 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6442
timestamp 1677677812
transform 1 0 4392 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6447
timestamp 1677677812
transform 1 0 4400 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6448
timestamp 1677677812
transform 1 0 4408 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6449
timestamp 1677677812
transform 1 0 4416 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6450
timestamp 1677677812
transform 1 0 4424 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6451
timestamp 1677677812
transform 1 0 4432 0 -1 2170
box -8 -3 16 105
use INVX2  INVX2_413
timestamp 1677677812
transform 1 0 4440 0 -1 2170
box -9 -3 26 105
use INVX2  INVX2_414
timestamp 1677677812
transform 1 0 4456 0 -1 2170
box -9 -3 26 105
use FILL  FILL_6452
timestamp 1677677812
transform 1 0 4472 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6453
timestamp 1677677812
transform 1 0 4480 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_18
timestamp 1677677812
transform 1 0 4488 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6454
timestamp 1677677812
transform 1 0 4520 0 -1 2170
box -8 -3 16 105
use AND2X2  AND2X2_19
timestamp 1677677812
transform 1 0 4528 0 -1 2170
box -8 -3 40 105
use FILL  FILL_6455
timestamp 1677677812
transform 1 0 4560 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6456
timestamp 1677677812
transform 1 0 4568 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6457
timestamp 1677677812
transform 1 0 4576 0 -1 2170
box -8 -3 16 105
use OAI22X1  OAI22X1_249
timestamp 1677677812
transform -1 0 4624 0 -1 2170
box -8 -3 46 105
use FILL  FILL_6458
timestamp 1677677812
transform 1 0 4624 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6459
timestamp 1677677812
transform 1 0 4632 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6461
timestamp 1677677812
transform 1 0 4640 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6463
timestamp 1677677812
transform 1 0 4648 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6474
timestamp 1677677812
transform 1 0 4656 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6475
timestamp 1677677812
transform 1 0 4664 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6476
timestamp 1677677812
transform 1 0 4672 0 -1 2170
box -8 -3 16 105
use FILL  FILL_6477
timestamp 1677677812
transform 1 0 4680 0 -1 2170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_363
timestamp 1677677812
transform 1 0 4688 0 -1 2170
box -8 -3 104 105
use FILL  FILL_6478
timestamp 1677677812
transform 1 0 4784 0 -1 2170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_53
timestamp 1677677812
transform 1 0 4843 0 1 2070
box -10 -3 10 3
use M3_M2  M3_M2_4988
timestamp 1677677812
transform 1 0 180 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5007
timestamp 1677677812
transform 1 0 164 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5558
timestamp 1677677812
transform 1 0 108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5559
timestamp 1677677812
transform 1 0 164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5560
timestamp 1677677812
transform 1 0 172 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5648
timestamp 1677677812
transform 1 0 84 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5078
timestamp 1677677812
transform 1 0 84 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5079
timestamp 1677677812
transform 1 0 156 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5105
timestamp 1677677812
transform 1 0 100 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5106
timestamp 1677677812
transform 1 0 172 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5649
timestamp 1677677812
transform 1 0 188 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5080
timestamp 1677677812
transform 1 0 188 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5008
timestamp 1677677812
transform 1 0 204 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_4974
timestamp 1677677812
transform 1 0 220 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4989
timestamp 1677677812
transform 1 0 244 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5561
timestamp 1677677812
transform 1 0 212 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5044
timestamp 1677677812
transform 1 0 220 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5562
timestamp 1677677812
transform 1 0 228 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5045
timestamp 1677677812
transform 1 0 236 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5563
timestamp 1677677812
transform 1 0 244 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5564
timestamp 1677677812
transform 1 0 252 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5650
timestamp 1677677812
transform 1 0 204 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5065
timestamp 1677677812
transform 1 0 212 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5046
timestamp 1677677812
transform 1 0 260 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5565
timestamp 1677677812
transform 1 0 268 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5047
timestamp 1677677812
transform 1 0 276 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5651
timestamp 1677677812
transform 1 0 236 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5652
timestamp 1677677812
transform 1 0 244 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5066
timestamp 1677677812
transform 1 0 252 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5653
timestamp 1677677812
transform 1 0 276 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5654
timestamp 1677677812
transform 1 0 284 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5081
timestamp 1677677812
transform 1 0 244 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5107
timestamp 1677677812
transform 1 0 276 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5566
timestamp 1677677812
transform 1 0 300 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5567
timestamp 1677677812
transform 1 0 308 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5048
timestamp 1677677812
transform 1 0 324 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5568
timestamp 1677677812
transform 1 0 332 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5067
timestamp 1677677812
transform 1 0 308 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5655
timestamp 1677677812
transform 1 0 316 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5656
timestamp 1677677812
transform 1 0 324 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5657
timestamp 1677677812
transform 1 0 340 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5108
timestamp 1677677812
transform 1 0 340 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5049
timestamp 1677677812
transform 1 0 356 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4990
timestamp 1677677812
transform 1 0 372 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5569
timestamp 1677677812
transform 1 0 364 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5725
timestamp 1677677812
transform 1 0 356 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5658
timestamp 1677677812
transform 1 0 380 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5009
timestamp 1677677812
transform 1 0 452 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5659
timestamp 1677677812
transform 1 0 468 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5082
timestamp 1677677812
transform 1 0 460 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4991
timestamp 1677677812
transform 1 0 524 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5050
timestamp 1677677812
transform 1 0 516 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5660
timestamp 1677677812
transform 1 0 516 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5570
timestamp 1677677812
transform 1 0 524 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5010
timestamp 1677677812
transform 1 0 540 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5571
timestamp 1677677812
transform 1 0 540 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5572
timestamp 1677677812
transform 1 0 556 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5051
timestamp 1677677812
transform 1 0 564 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5661
timestamp 1677677812
transform 1 0 548 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5068
timestamp 1677677812
transform 1 0 556 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5083
timestamp 1677677812
transform 1 0 548 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5573
timestamp 1677677812
transform 1 0 580 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5662
timestamp 1677677812
transform 1 0 572 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5069
timestamp 1677677812
transform 1 0 588 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_4992
timestamp 1677677812
transform 1 0 612 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5663
timestamp 1677677812
transform 1 0 612 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4984
timestamp 1677677812
transform 1 0 692 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_4993
timestamp 1677677812
transform 1 0 676 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5574
timestamp 1677677812
transform 1 0 668 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5575
timestamp 1677677812
transform 1 0 684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5664
timestamp 1677677812
transform 1 0 668 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5665
timestamp 1677677812
transform 1 0 708 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5576
timestamp 1677677812
transform 1 0 716 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5070
timestamp 1677677812
transform 1 0 732 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5577
timestamp 1677677812
transform 1 0 796 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5578
timestamp 1677677812
transform 1 0 852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5666
timestamp 1677677812
transform 1 0 772 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5071
timestamp 1677677812
transform 1 0 836 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5084
timestamp 1677677812
transform 1 0 852 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5726
timestamp 1677677812
transform 1 0 860 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5667
timestamp 1677677812
transform 1 0 964 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5011
timestamp 1677677812
transform 1 0 980 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5727
timestamp 1677677812
transform 1 0 980 0 1 1995
box -2 -2 2 2
use M3_M2  M3_M2_5012
timestamp 1677677812
transform 1 0 996 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5579
timestamp 1677677812
transform 1 0 996 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5013
timestamp 1677677812
transform 1 0 1012 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5668
timestamp 1677677812
transform 1 0 1012 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5580
timestamp 1677677812
transform 1 0 1036 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4994
timestamp 1677677812
transform 1 0 1052 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5581
timestamp 1677677812
transform 1 0 1052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5728
timestamp 1677677812
transform 1 0 1100 0 1 1995
box -2 -2 2 2
use M2_M1  M2_M1_5669
timestamp 1677677812
transform 1 0 1132 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5670
timestamp 1677677812
transform 1 0 1140 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5014
timestamp 1677677812
transform 1 0 1260 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5582
timestamp 1677677812
transform 1 0 1260 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5671
timestamp 1677677812
transform 1 0 1268 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5109
timestamp 1677677812
transform 1 0 1276 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5672
timestamp 1677677812
transform 1 0 1332 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4995
timestamp 1677677812
transform 1 0 1372 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5583
timestamp 1677677812
transform 1 0 1364 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4970
timestamp 1677677812
transform 1 0 1396 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5015
timestamp 1677677812
transform 1 0 1436 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5110
timestamp 1677677812
transform 1 0 1436 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5673
timestamp 1677677812
transform 1 0 1508 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5016
timestamp 1677677812
transform 1 0 1572 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5584
timestamp 1677677812
transform 1 0 1564 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5585
timestamp 1677677812
transform 1 0 1572 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5674
timestamp 1677677812
transform 1 0 1588 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5085
timestamp 1677677812
transform 1 0 1588 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5017
timestamp 1677677812
transform 1 0 1604 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5675
timestamp 1677677812
transform 1 0 1604 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5086
timestamp 1677677812
transform 1 0 1620 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4975
timestamp 1677677812
transform 1 0 1684 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5586
timestamp 1677677812
transform 1 0 1676 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5587
timestamp 1677677812
transform 1 0 1684 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5588
timestamp 1677677812
transform 1 0 1708 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5676
timestamp 1677677812
transform 1 0 1700 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4976
timestamp 1677677812
transform 1 0 1732 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5677
timestamp 1677677812
transform 1 0 1740 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5052
timestamp 1677677812
transform 1 0 1788 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5678
timestamp 1677677812
transform 1 0 1788 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5589
timestamp 1677677812
transform 1 0 1804 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5018
timestamp 1677677812
transform 1 0 1836 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5590
timestamp 1677677812
transform 1 0 1828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5591
timestamp 1677677812
transform 1 0 1836 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5548
timestamp 1677677812
transform 1 0 1860 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_5019
timestamp 1677677812
transform 1 0 1868 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5549
timestamp 1677677812
transform 1 0 1924 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_5020
timestamp 1677677812
transform 1 0 1924 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5053
timestamp 1677677812
transform 1 0 1940 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5679
timestamp 1677677812
transform 1 0 1956 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4996
timestamp 1677677812
transform 1 0 1988 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5054
timestamp 1677677812
transform 1 0 1988 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5021
timestamp 1677677812
transform 1 0 2028 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5592
timestamp 1677677812
transform 1 0 2028 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5593
timestamp 1677677812
transform 1 0 2044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5680
timestamp 1677677812
transform 1 0 2020 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5681
timestamp 1677677812
transform 1 0 2036 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5682
timestamp 1677677812
transform 1 0 2052 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5683
timestamp 1677677812
transform 1 0 2060 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5087
timestamp 1677677812
transform 1 0 2052 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5594
timestamp 1677677812
transform 1 0 2148 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4971
timestamp 1677677812
transform 1 0 2244 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5595
timestamp 1677677812
transform 1 0 2212 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5684
timestamp 1677677812
transform 1 0 2164 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5111
timestamp 1677677812
transform 1 0 2180 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5596
timestamp 1677677812
transform 1 0 2252 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5022
timestamp 1677677812
transform 1 0 2332 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5597
timestamp 1677677812
transform 1 0 2332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5598
timestamp 1677677812
transform 1 0 2356 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5685
timestamp 1677677812
transform 1 0 2364 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5088
timestamp 1677677812
transform 1 0 2364 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5599
timestamp 1677677812
transform 1 0 2380 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5112
timestamp 1677677812
transform 1 0 2380 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5023
timestamp 1677677812
transform 1 0 2396 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5024
timestamp 1677677812
transform 1 0 2468 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5686
timestamp 1677677812
transform 1 0 2468 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4997
timestamp 1677677812
transform 1 0 2484 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5600
timestamp 1677677812
transform 1 0 2484 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5113
timestamp 1677677812
transform 1 0 2484 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_4972
timestamp 1677677812
transform 1 0 2508 0 1 2065
box -3 -3 3 3
use M2_M1  M2_M1_5687
timestamp 1677677812
transform 1 0 2556 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5114
timestamp 1677677812
transform 1 0 2548 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5688
timestamp 1677677812
transform 1 0 2572 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4977
timestamp 1677677812
transform 1 0 2596 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4978
timestamp 1677677812
transform 1 0 2620 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5025
timestamp 1677677812
transform 1 0 2604 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5601
timestamp 1677677812
transform 1 0 2588 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5055
timestamp 1677677812
transform 1 0 2596 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5602
timestamp 1677677812
transform 1 0 2604 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5603
timestamp 1677677812
transform 1 0 2620 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4979
timestamp 1677677812
transform 1 0 2660 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5026
timestamp 1677677812
transform 1 0 2652 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5689
timestamp 1677677812
transform 1 0 2652 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4998
timestamp 1677677812
transform 1 0 2692 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5027
timestamp 1677677812
transform 1 0 2748 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5604
timestamp 1677677812
transform 1 0 2692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5605
timestamp 1677677812
transform 1 0 2748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5690
timestamp 1677677812
transform 1 0 2668 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5072
timestamp 1677677812
transform 1 0 2732 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5606
timestamp 1677677812
transform 1 0 2820 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5691
timestamp 1677677812
transform 1 0 2860 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5028
timestamp 1677677812
transform 1 0 2900 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5552
timestamp 1677677812
transform 1 0 2908 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5607
timestamp 1677677812
transform 1 0 2924 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5056
timestamp 1677677812
transform 1 0 2940 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_4980
timestamp 1677677812
transform 1 0 2964 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_5029
timestamp 1677677812
transform 1 0 2956 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5608
timestamp 1677677812
transform 1 0 2948 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5692
timestamp 1677677812
transform 1 0 2940 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5693
timestamp 1677677812
transform 1 0 2956 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5030
timestamp 1677677812
transform 1 0 2972 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5609
timestamp 1677677812
transform 1 0 2972 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5057
timestamp 1677677812
transform 1 0 2980 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5610
timestamp 1677677812
transform 1 0 2988 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5115
timestamp 1677677812
transform 1 0 2972 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5611
timestamp 1677677812
transform 1 0 3020 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5612
timestamp 1677677812
transform 1 0 3036 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5694
timestamp 1677677812
transform 1 0 3028 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5695
timestamp 1677677812
transform 1 0 3044 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5089
timestamp 1677677812
transform 1 0 3028 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5058
timestamp 1677677812
transform 1 0 3068 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5613
timestamp 1677677812
transform 1 0 3076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5614
timestamp 1677677812
transform 1 0 3108 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5696
timestamp 1677677812
transform 1 0 3068 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5697
timestamp 1677677812
transform 1 0 3156 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5090
timestamp 1677677812
transform 1 0 3108 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5091
timestamp 1677677812
transform 1 0 3140 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5116
timestamp 1677677812
transform 1 0 3108 0 1 1985
box -3 -3 3 3
use M2_M1  M2_M1_5698
timestamp 1677677812
transform 1 0 3172 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5553
timestamp 1677677812
transform 1 0 3260 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5615
timestamp 1677677812
transform 1 0 3268 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4985
timestamp 1677677812
transform 1 0 3284 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5550
timestamp 1677677812
transform 1 0 3284 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_4999
timestamp 1677677812
transform 1 0 3292 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5554
timestamp 1677677812
transform 1 0 3300 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5616
timestamp 1677677812
transform 1 0 3292 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5092
timestamp 1677677812
transform 1 0 3308 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5699
timestamp 1677677812
transform 1 0 3332 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5093
timestamp 1677677812
transform 1 0 3332 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5117
timestamp 1677677812
transform 1 0 3324 0 1 1985
box -3 -3 3 3
use M3_M2  M3_M2_5031
timestamp 1677677812
transform 1 0 3348 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5617
timestamp 1677677812
transform 1 0 3348 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5700
timestamp 1677677812
transform 1 0 3372 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5032
timestamp 1677677812
transform 1 0 3404 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5618
timestamp 1677677812
transform 1 0 3404 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5000
timestamp 1677677812
transform 1 0 3452 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5555
timestamp 1677677812
transform 1 0 3452 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5619
timestamp 1677677812
transform 1 0 3420 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5059
timestamp 1677677812
transform 1 0 3444 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5701
timestamp 1677677812
transform 1 0 3428 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5702
timestamp 1677677812
transform 1 0 3444 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5620
timestamp 1677677812
transform 1 0 3476 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_4981
timestamp 1677677812
transform 1 0 3500 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5551
timestamp 1677677812
transform 1 0 3500 0 1 2035
box -2 -2 2 2
use M3_M2  M3_M2_5001
timestamp 1677677812
transform 1 0 3516 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5621
timestamp 1677677812
transform 1 0 3508 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5002
timestamp 1677677812
transform 1 0 3532 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5703
timestamp 1677677812
transform 1 0 3540 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5094
timestamp 1677677812
transform 1 0 3540 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5033
timestamp 1677677812
transform 1 0 3580 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5060
timestamp 1677677812
transform 1 0 3620 0 1 2015
box -3 -3 3 3
use M3_M2  M3_M2_5095
timestamp 1677677812
transform 1 0 3620 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4973
timestamp 1677677812
transform 1 0 3652 0 1 2065
box -3 -3 3 3
use M3_M2  M3_M2_5003
timestamp 1677677812
transform 1 0 3660 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5556
timestamp 1677677812
transform 1 0 3660 0 1 2025
box -2 -2 2 2
use M3_M2  M3_M2_5034
timestamp 1677677812
transform 1 0 3668 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5061
timestamp 1677677812
transform 1 0 3660 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5622
timestamp 1677677812
transform 1 0 3668 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5073
timestamp 1677677812
transform 1 0 3652 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5704
timestamp 1677677812
transform 1 0 3660 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5074
timestamp 1677677812
transform 1 0 3668 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5062
timestamp 1677677812
transform 1 0 3692 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5623
timestamp 1677677812
transform 1 0 3708 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5075
timestamp 1677677812
transform 1 0 3708 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5035
timestamp 1677677812
transform 1 0 3748 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5557
timestamp 1677677812
transform 1 0 3812 0 1 2025
box -2 -2 2 2
use M2_M1  M2_M1_5624
timestamp 1677677812
transform 1 0 3748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5625
timestamp 1677677812
transform 1 0 3804 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5705
timestamp 1677677812
transform 1 0 3724 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4986
timestamp 1677677812
transform 1 0 3860 0 1 2045
box -3 -3 3 3
use M2_M1  M2_M1_5626
timestamp 1677677812
transform 1 0 3828 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5627
timestamp 1677677812
transform 1 0 3852 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5706
timestamp 1677677812
transform 1 0 3836 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5707
timestamp 1677677812
transform 1 0 3852 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5096
timestamp 1677677812
transform 1 0 3852 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5036
timestamp 1677677812
transform 1 0 3876 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5628
timestamp 1677677812
transform 1 0 3876 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5004
timestamp 1677677812
transform 1 0 3916 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5037
timestamp 1677677812
transform 1 0 3932 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5629
timestamp 1677677812
transform 1 0 3900 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5063
timestamp 1677677812
transform 1 0 3908 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5630
timestamp 1677677812
transform 1 0 3916 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5631
timestamp 1677677812
transform 1 0 3932 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5708
timestamp 1677677812
transform 1 0 3900 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5709
timestamp 1677677812
transform 1 0 3908 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5097
timestamp 1677677812
transform 1 0 3924 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5710
timestamp 1677677812
transform 1 0 3948 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_4987
timestamp 1677677812
transform 1 0 4036 0 1 2045
box -3 -3 3 3
use M3_M2  M3_M2_5038
timestamp 1677677812
transform 1 0 4036 0 1 2025
box -3 -3 3 3
use M3_M2  M3_M2_5039
timestamp 1677677812
transform 1 0 4068 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5632
timestamp 1677677812
transform 1 0 3988 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5633
timestamp 1677677812
transform 1 0 4044 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5634
timestamp 1677677812
transform 1 0 4052 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5711
timestamp 1677677812
transform 1 0 3964 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5076
timestamp 1677677812
transform 1 0 4036 0 1 2005
box -3 -3 3 3
use M3_M2  M3_M2_5064
timestamp 1677677812
transform 1 0 4068 0 1 2015
box -3 -3 3 3
use M2_M1  M2_M1_5635
timestamp 1677677812
transform 1 0 4076 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5712
timestamp 1677677812
transform 1 0 4052 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5713
timestamp 1677677812
transform 1 0 4068 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5077
timestamp 1677677812
transform 1 0 4076 0 1 2005
box -3 -3 3 3
use M2_M1  M2_M1_5636
timestamp 1677677812
transform 1 0 4092 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5714
timestamp 1677677812
transform 1 0 4084 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5098
timestamp 1677677812
transform 1 0 4052 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5099
timestamp 1677677812
transform 1 0 4068 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_4982
timestamp 1677677812
transform 1 0 4156 0 1 2055
box -3 -3 3 3
use M3_M2  M3_M2_4983
timestamp 1677677812
transform 1 0 4212 0 1 2055
box -3 -3 3 3
use M2_M1  M2_M1_5637
timestamp 1677677812
transform 1 0 4164 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5715
timestamp 1677677812
transform 1 0 4212 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5100
timestamp 1677677812
transform 1 0 4164 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5101
timestamp 1677677812
transform 1 0 4212 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5040
timestamp 1677677812
transform 1 0 4284 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5638
timestamp 1677677812
transform 1 0 4284 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5716
timestamp 1677677812
transform 1 0 4236 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5102
timestamp 1677677812
transform 1 0 4236 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5639
timestamp 1677677812
transform 1 0 4332 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5640
timestamp 1677677812
transform 1 0 4340 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5641
timestamp 1677677812
transform 1 0 4356 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5041
timestamp 1677677812
transform 1 0 4372 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5717
timestamp 1677677812
transform 1 0 4364 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5718
timestamp 1677677812
transform 1 0 4372 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5103
timestamp 1677677812
transform 1 0 4364 0 1 1995
box -3 -3 3 3
use M3_M2  M3_M2_5104
timestamp 1677677812
transform 1 0 4396 0 1 1995
box -3 -3 3 3
use M2_M1  M2_M1_5642
timestamp 1677677812
transform 1 0 4460 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5719
timestamp 1677677812
transform 1 0 4452 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5643
timestamp 1677677812
transform 1 0 4492 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5720
timestamp 1677677812
transform 1 0 4524 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5721
timestamp 1677677812
transform 1 0 4572 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5005
timestamp 1677677812
transform 1 0 4604 0 1 2035
box -3 -3 3 3
use M2_M1  M2_M1_5644
timestamp 1677677812
transform 1 0 4596 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5645
timestamp 1677677812
transform 1 0 4620 0 1 2015
box -2 -2 2 2
use M3_M2  M3_M2_5042
timestamp 1677677812
transform 1 0 4628 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5722
timestamp 1677677812
transform 1 0 4628 0 1 2005
box -2 -2 2 2
use M3_M2  M3_M2_5006
timestamp 1677677812
transform 1 0 4692 0 1 2035
box -3 -3 3 3
use M3_M2  M3_M2_5043
timestamp 1677677812
transform 1 0 4748 0 1 2025
box -3 -3 3 3
use M2_M1  M2_M1_5646
timestamp 1677677812
transform 1 0 4692 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5647
timestamp 1677677812
transform 1 0 4748 0 1 2015
box -2 -2 2 2
use M2_M1  M2_M1_5723
timestamp 1677677812
transform 1 0 4652 0 1 2005
box -2 -2 2 2
use M2_M1  M2_M1_5724
timestamp 1677677812
transform 1 0 4668 0 1 2005
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_54
timestamp 1677677812
transform 1 0 48 0 1 1970
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_364
timestamp 1677677812
transform 1 0 72 0 1 1970
box -8 -3 104 105
use BUFX2  BUFX2_63
timestamp 1677677812
transform 1 0 168 0 1 1970
box -5 -3 28 105
use FILL  FILL_6479
timestamp 1677677812
transform 1 0 192 0 1 1970
box -8 -3 16 105
use FILL  FILL_6480
timestamp 1677677812
transform 1 0 200 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_256
timestamp 1677677812
transform -1 0 248 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_5118
timestamp 1677677812
transform 1 0 284 0 1 1975
box -3 -3 3 3
use AOI22X1  AOI22X1_257
timestamp 1677677812
transform -1 0 288 0 1 1970
box -8 -3 46 105
use FILL  FILL_6481
timestamp 1677677812
transform 1 0 288 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5119
timestamp 1677677812
transform 1 0 316 0 1 1975
box -3 -3 3 3
use INVX2  INVX2_416
timestamp 1677677812
transform -1 0 312 0 1 1970
box -9 -3 26 105
use AOI22X1  AOI22X1_258
timestamp 1677677812
transform -1 0 352 0 1 1970
box -8 -3 46 105
use FILL  FILL_6482
timestamp 1677677812
transform 1 0 352 0 1 1970
box -8 -3 16 105
use FILL  FILL_6483
timestamp 1677677812
transform 1 0 360 0 1 1970
box -8 -3 16 105
use FILL  FILL_6484
timestamp 1677677812
transform 1 0 368 0 1 1970
box -8 -3 16 105
use FILL  FILL_6485
timestamp 1677677812
transform 1 0 376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6486
timestamp 1677677812
transform 1 0 384 0 1 1970
box -8 -3 16 105
use FILL  FILL_6487
timestamp 1677677812
transform 1 0 392 0 1 1970
box -8 -3 16 105
use FILL  FILL_6488
timestamp 1677677812
transform 1 0 400 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5120
timestamp 1677677812
transform 1 0 420 0 1 1975
box -3 -3 3 3
use FILL  FILL_6489
timestamp 1677677812
transform 1 0 408 0 1 1970
box -8 -3 16 105
use FILL  FILL_6490
timestamp 1677677812
transform 1 0 416 0 1 1970
box -8 -3 16 105
use FILL  FILL_6491
timestamp 1677677812
transform 1 0 424 0 1 1970
box -8 -3 16 105
use FILL  FILL_6492
timestamp 1677677812
transform 1 0 432 0 1 1970
box -8 -3 16 105
use FILL  FILL_6493
timestamp 1677677812
transform 1 0 440 0 1 1970
box -8 -3 16 105
use FILL  FILL_6494
timestamp 1677677812
transform 1 0 448 0 1 1970
box -8 -3 16 105
use FILL  FILL_6495
timestamp 1677677812
transform 1 0 456 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_64
timestamp 1677677812
transform -1 0 488 0 1 1970
box -5 -3 28 105
use FILL  FILL_6496
timestamp 1677677812
transform 1 0 488 0 1 1970
box -8 -3 16 105
use FILL  FILL_6497
timestamp 1677677812
transform 1 0 496 0 1 1970
box -8 -3 16 105
use FILL  FILL_6498
timestamp 1677677812
transform 1 0 504 0 1 1970
box -8 -3 16 105
use FILL  FILL_6499
timestamp 1677677812
transform 1 0 512 0 1 1970
box -8 -3 16 105
use FILL  FILL_6500
timestamp 1677677812
transform 1 0 520 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_251
timestamp 1677677812
transform -1 0 568 0 1 1970
box -8 -3 46 105
use M3_M2  M3_M2_5121
timestamp 1677677812
transform 1 0 580 0 1 1975
box -3 -3 3 3
use FILL  FILL_6501
timestamp 1677677812
transform 1 0 568 0 1 1970
box -8 -3 16 105
use FILL  FILL_6502
timestamp 1677677812
transform 1 0 576 0 1 1970
box -8 -3 16 105
use FILL  FILL_6503
timestamp 1677677812
transform 1 0 584 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_65
timestamp 1677677812
transform 1 0 592 0 1 1970
box -5 -3 28 105
use FILL  FILL_6504
timestamp 1677677812
transform 1 0 616 0 1 1970
box -8 -3 16 105
use FILL  FILL_6516
timestamp 1677677812
transform 1 0 624 0 1 1970
box -8 -3 16 105
use FILL  FILL_6518
timestamp 1677677812
transform 1 0 632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6520
timestamp 1677677812
transform 1 0 640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6522
timestamp 1677677812
transform 1 0 648 0 1 1970
box -8 -3 16 105
use FILL  FILL_6523
timestamp 1677677812
transform 1 0 656 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_259
timestamp 1677677812
transform 1 0 664 0 1 1970
box -8 -3 46 105
use FILL  FILL_6524
timestamp 1677677812
transform 1 0 704 0 1 1970
box -8 -3 16 105
use FILL  FILL_6525
timestamp 1677677812
transform 1 0 712 0 1 1970
box -8 -3 16 105
use FILL  FILL_6526
timestamp 1677677812
transform 1 0 720 0 1 1970
box -8 -3 16 105
use FILL  FILL_6527
timestamp 1677677812
transform 1 0 728 0 1 1970
box -8 -3 16 105
use FILL  FILL_6528
timestamp 1677677812
transform 1 0 736 0 1 1970
box -8 -3 16 105
use FILL  FILL_6529
timestamp 1677677812
transform 1 0 744 0 1 1970
box -8 -3 16 105
use FILL  FILL_6535
timestamp 1677677812
transform 1 0 752 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_368
timestamp 1677677812
transform 1 0 760 0 1 1970
box -8 -3 104 105
use FILL  FILL_6537
timestamp 1677677812
transform 1 0 856 0 1 1970
box -8 -3 16 105
use FILL  FILL_6546
timestamp 1677677812
transform 1 0 864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6548
timestamp 1677677812
transform 1 0 872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6550
timestamp 1677677812
transform 1 0 880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6552
timestamp 1677677812
transform 1 0 888 0 1 1970
box -8 -3 16 105
use FILL  FILL_6554
timestamp 1677677812
transform 1 0 896 0 1 1970
box -8 -3 16 105
use FILL  FILL_6556
timestamp 1677677812
transform 1 0 904 0 1 1970
box -8 -3 16 105
use FILL  FILL_6558
timestamp 1677677812
transform 1 0 912 0 1 1970
box -8 -3 16 105
use FILL  FILL_6560
timestamp 1677677812
transform 1 0 920 0 1 1970
box -8 -3 16 105
use FILL  FILL_6562
timestamp 1677677812
transform 1 0 928 0 1 1970
box -8 -3 16 105
use FILL  FILL_6564
timestamp 1677677812
transform 1 0 936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6566
timestamp 1677677812
transform 1 0 944 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_62
timestamp 1677677812
transform 1 0 952 0 1 1970
box -8 -3 32 105
use FILL  FILL_6568
timestamp 1677677812
transform 1 0 976 0 1 1970
box -8 -3 16 105
use FILL  FILL_6573
timestamp 1677677812
transform 1 0 984 0 1 1970
box -8 -3 16 105
use FILL  FILL_6575
timestamp 1677677812
transform 1 0 992 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_63
timestamp 1677677812
transform 1 0 1000 0 1 1970
box -8 -3 32 105
use FILL  FILL_6577
timestamp 1677677812
transform 1 0 1024 0 1 1970
box -8 -3 16 105
use FILL  FILL_6578
timestamp 1677677812
transform 1 0 1032 0 1 1970
box -8 -3 16 105
use FILL  FILL_6579
timestamp 1677677812
transform 1 0 1040 0 1 1970
box -8 -3 16 105
use FILL  FILL_6580
timestamp 1677677812
transform 1 0 1048 0 1 1970
box -8 -3 16 105
use FILL  FILL_6581
timestamp 1677677812
transform 1 0 1056 0 1 1970
box -8 -3 16 105
use FILL  FILL_6585
timestamp 1677677812
transform 1 0 1064 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_70
timestamp 1677677812
transform 1 0 1072 0 1 1970
box -5 -3 28 105
use FILL  FILL_6587
timestamp 1677677812
transform 1 0 1096 0 1 1970
box -8 -3 16 105
use FILL  FILL_6592
timestamp 1677677812
transform 1 0 1104 0 1 1970
box -8 -3 16 105
use FILL  FILL_6594
timestamp 1677677812
transform 1 0 1112 0 1 1970
box -8 -3 16 105
use FILL  FILL_6596
timestamp 1677677812
transform 1 0 1120 0 1 1970
box -8 -3 16 105
use FILL  FILL_6598
timestamp 1677677812
transform 1 0 1128 0 1 1970
box -8 -3 16 105
use FILL  FILL_6600
timestamp 1677677812
transform 1 0 1136 0 1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_64
timestamp 1677677812
transform 1 0 1144 0 1 1970
box -8 -3 32 105
use FILL  FILL_6602
timestamp 1677677812
transform 1 0 1168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6603
timestamp 1677677812
transform 1 0 1176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6604
timestamp 1677677812
transform 1 0 1184 0 1 1970
box -8 -3 16 105
use FILL  FILL_6605
timestamp 1677677812
transform 1 0 1192 0 1 1970
box -8 -3 16 105
use FILL  FILL_6608
timestamp 1677677812
transform 1 0 1200 0 1 1970
box -8 -3 16 105
use FILL  FILL_6610
timestamp 1677677812
transform 1 0 1208 0 1 1970
box -8 -3 16 105
use FILL  FILL_6612
timestamp 1677677812
transform 1 0 1216 0 1 1970
box -8 -3 16 105
use FILL  FILL_6614
timestamp 1677677812
transform 1 0 1224 0 1 1970
box -8 -3 16 105
use FILL  FILL_6616
timestamp 1677677812
transform 1 0 1232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6618
timestamp 1677677812
transform 1 0 1240 0 1 1970
box -8 -3 16 105
use FILL  FILL_6620
timestamp 1677677812
transform 1 0 1248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6622
timestamp 1677677812
transform 1 0 1256 0 1 1970
box -8 -3 16 105
use FILL  FILL_6624
timestamp 1677677812
transform 1 0 1264 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_421
timestamp 1677677812
transform 1 0 1272 0 1 1970
box -9 -3 26 105
use FILL  FILL_6626
timestamp 1677677812
transform 1 0 1288 0 1 1970
box -8 -3 16 105
use FILL  FILL_6630
timestamp 1677677812
transform 1 0 1296 0 1 1970
box -8 -3 16 105
use FILL  FILL_6632
timestamp 1677677812
transform 1 0 1304 0 1 1970
box -8 -3 16 105
use FILL  FILL_6634
timestamp 1677677812
transform 1 0 1312 0 1 1970
box -8 -3 16 105
use FILL  FILL_6636
timestamp 1677677812
transform 1 0 1320 0 1 1970
box -8 -3 16 105
use FILL  FILL_6637
timestamp 1677677812
transform 1 0 1328 0 1 1970
box -8 -3 16 105
use FILL  FILL_6638
timestamp 1677677812
transform 1 0 1336 0 1 1970
box -8 -3 16 105
use FILL  FILL_6639
timestamp 1677677812
transform 1 0 1344 0 1 1970
box -8 -3 16 105
use FILL  FILL_6640
timestamp 1677677812
transform 1 0 1352 0 1 1970
box -8 -3 16 105
use FILL  FILL_6641
timestamp 1677677812
transform 1 0 1360 0 1 1970
box -8 -3 16 105
use FILL  FILL_6642
timestamp 1677677812
transform 1 0 1368 0 1 1970
box -8 -3 16 105
use FILL  FILL_6643
timestamp 1677677812
transform 1 0 1376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6644
timestamp 1677677812
transform 1 0 1384 0 1 1970
box -8 -3 16 105
use FILL  FILL_6645
timestamp 1677677812
transform 1 0 1392 0 1 1970
box -8 -3 16 105
use FILL  FILL_6646
timestamp 1677677812
transform 1 0 1400 0 1 1970
box -8 -3 16 105
use FILL  FILL_6647
timestamp 1677677812
transform 1 0 1408 0 1 1970
box -8 -3 16 105
use FILL  FILL_6648
timestamp 1677677812
transform 1 0 1416 0 1 1970
box -8 -3 16 105
use FILL  FILL_6650
timestamp 1677677812
transform 1 0 1424 0 1 1970
box -8 -3 16 105
use FILL  FILL_6652
timestamp 1677677812
transform 1 0 1432 0 1 1970
box -8 -3 16 105
use FILL  FILL_6654
timestamp 1677677812
transform 1 0 1440 0 1 1970
box -8 -3 16 105
use FILL  FILL_6656
timestamp 1677677812
transform 1 0 1448 0 1 1970
box -8 -3 16 105
use FILL  FILL_6657
timestamp 1677677812
transform 1 0 1456 0 1 1970
box -8 -3 16 105
use FILL  FILL_6658
timestamp 1677677812
transform 1 0 1464 0 1 1970
box -8 -3 16 105
use FILL  FILL_6659
timestamp 1677677812
transform 1 0 1472 0 1 1970
box -8 -3 16 105
use FILL  FILL_6660
timestamp 1677677812
transform 1 0 1480 0 1 1970
box -8 -3 16 105
use FILL  FILL_6661
timestamp 1677677812
transform 1 0 1488 0 1 1970
box -8 -3 16 105
use FILL  FILL_6664
timestamp 1677677812
transform 1 0 1496 0 1 1970
box -8 -3 16 105
use FILL  FILL_6666
timestamp 1677677812
transform 1 0 1504 0 1 1970
box -8 -3 16 105
use FILL  FILL_6668
timestamp 1677677812
transform 1 0 1512 0 1 1970
box -8 -3 16 105
use FILL  FILL_6670
timestamp 1677677812
transform 1 0 1520 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_71
timestamp 1677677812
transform -1 0 1552 0 1 1970
box -5 -3 28 105
use FILL  FILL_6671
timestamp 1677677812
transform 1 0 1552 0 1 1970
box -8 -3 16 105
use FILL  FILL_6672
timestamp 1677677812
transform 1 0 1560 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5122
timestamp 1677677812
transform 1 0 1604 0 1 1975
box -3 -3 3 3
use BUFX2  BUFX2_72
timestamp 1677677812
transform 1 0 1568 0 1 1970
box -5 -3 28 105
use FILL  FILL_6677
timestamp 1677677812
transform 1 0 1592 0 1 1970
box -8 -3 16 105
use FILL  FILL_6678
timestamp 1677677812
transform 1 0 1600 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_73
timestamp 1677677812
transform -1 0 1632 0 1 1970
box -5 -3 28 105
use FILL  FILL_6679
timestamp 1677677812
transform 1 0 1632 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5123
timestamp 1677677812
transform 1 0 1652 0 1 1975
box -3 -3 3 3
use FILL  FILL_6680
timestamp 1677677812
transform 1 0 1640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6681
timestamp 1677677812
transform 1 0 1648 0 1 1970
box -8 -3 16 105
use FILL  FILL_6687
timestamp 1677677812
transform 1 0 1656 0 1 1970
box -8 -3 16 105
use FILL  FILL_6689
timestamp 1677677812
transform 1 0 1664 0 1 1970
box -8 -3 16 105
use FILL  FILL_6691
timestamp 1677677812
transform 1 0 1672 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_76
timestamp 1677677812
transform 1 0 1680 0 1 1970
box -5 -3 28 105
use FILL  FILL_6692
timestamp 1677677812
transform 1 0 1704 0 1 1970
box -8 -3 16 105
use FILL  FILL_6695
timestamp 1677677812
transform 1 0 1712 0 1 1970
box -8 -3 16 105
use FILL  FILL_6697
timestamp 1677677812
transform 1 0 1720 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_423
timestamp 1677677812
transform -1 0 1744 0 1 1970
box -9 -3 26 105
use FILL  FILL_6698
timestamp 1677677812
transform 1 0 1744 0 1 1970
box -8 -3 16 105
use FILL  FILL_6699
timestamp 1677677812
transform 1 0 1752 0 1 1970
box -8 -3 16 105
use FILL  FILL_6702
timestamp 1677677812
transform 1 0 1760 0 1 1970
box -8 -3 16 105
use FILL  FILL_6704
timestamp 1677677812
transform 1 0 1768 0 1 1970
box -8 -3 16 105
use FILL  FILL_6706
timestamp 1677677812
transform 1 0 1776 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_79
timestamp 1677677812
transform -1 0 1808 0 1 1970
box -5 -3 28 105
use FILL  FILL_6707
timestamp 1677677812
transform 1 0 1808 0 1 1970
box -8 -3 16 105
use FILL  FILL_6710
timestamp 1677677812
transform 1 0 1816 0 1 1970
box -8 -3 16 105
use FILL  FILL_6711
timestamp 1677677812
transform 1 0 1824 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_81
timestamp 1677677812
transform 1 0 1832 0 1 1970
box -5 -3 28 105
use FILL  FILL_6712
timestamp 1677677812
transform 1 0 1856 0 1 1970
box -8 -3 16 105
use FILL  FILL_6716
timestamp 1677677812
transform 1 0 1864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6718
timestamp 1677677812
transform 1 0 1872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6720
timestamp 1677677812
transform 1 0 1880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6722
timestamp 1677677812
transform 1 0 1888 0 1 1970
box -8 -3 16 105
use FILL  FILL_6724
timestamp 1677677812
transform 1 0 1896 0 1 1970
box -8 -3 16 105
use FILL  FILL_6725
timestamp 1677677812
transform 1 0 1904 0 1 1970
box -8 -3 16 105
use FILL  FILL_6726
timestamp 1677677812
transform 1 0 1912 0 1 1970
box -8 -3 16 105
use FILL  FILL_6728
timestamp 1677677812
transform 1 0 1920 0 1 1970
box -8 -3 16 105
use FILL  FILL_6730
timestamp 1677677812
transform 1 0 1928 0 1 1970
box -8 -3 16 105
use FILL  FILL_6732
timestamp 1677677812
transform 1 0 1936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6734
timestamp 1677677812
transform 1 0 1944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6735
timestamp 1677677812
transform 1 0 1952 0 1 1970
box -8 -3 16 105
use FILL  FILL_6736
timestamp 1677677812
transform 1 0 1960 0 1 1970
box -8 -3 16 105
use FILL  FILL_6737
timestamp 1677677812
transform 1 0 1968 0 1 1970
box -8 -3 16 105
use FILL  FILL_6738
timestamp 1677677812
transform 1 0 1976 0 1 1970
box -8 -3 16 105
use FILL  FILL_6739
timestamp 1677677812
transform 1 0 1984 0 1 1970
box -8 -3 16 105
use FILL  FILL_6740
timestamp 1677677812
transform 1 0 1992 0 1 1970
box -8 -3 16 105
use FILL  FILL_6743
timestamp 1677677812
transform 1 0 2000 0 1 1970
box -8 -3 16 105
use FILL  FILL_6745
timestamp 1677677812
transform 1 0 2008 0 1 1970
box -8 -3 16 105
use FILL  FILL_6746
timestamp 1677677812
transform 1 0 2016 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_263
timestamp 1677677812
transform -1 0 2064 0 1 1970
box -8 -3 46 105
use FILL  FILL_6747
timestamp 1677677812
transform 1 0 2064 0 1 1970
box -8 -3 16 105
use FILL  FILL_6748
timestamp 1677677812
transform 1 0 2072 0 1 1970
box -8 -3 16 105
use FILL  FILL_6749
timestamp 1677677812
transform 1 0 2080 0 1 1970
box -8 -3 16 105
use FILL  FILL_6750
timestamp 1677677812
transform 1 0 2088 0 1 1970
box -8 -3 16 105
use FILL  FILL_6751
timestamp 1677677812
transform 1 0 2096 0 1 1970
box -8 -3 16 105
use FILL  FILL_6752
timestamp 1677677812
transform 1 0 2104 0 1 1970
box -8 -3 16 105
use FILL  FILL_6753
timestamp 1677677812
transform 1 0 2112 0 1 1970
box -8 -3 16 105
use FILL  FILL_6756
timestamp 1677677812
transform 1 0 2120 0 1 1970
box -8 -3 16 105
use FILL  FILL_6758
timestamp 1677677812
transform 1 0 2128 0 1 1970
box -8 -3 16 105
use FILL  FILL_6760
timestamp 1677677812
transform 1 0 2136 0 1 1970
box -8 -3 16 105
use FILL  FILL_6762
timestamp 1677677812
transform 1 0 2144 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_371
timestamp 1677677812
transform 1 0 2152 0 1 1970
box -8 -3 104 105
use FILL  FILL_6764
timestamp 1677677812
transform 1 0 2248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6765
timestamp 1677677812
transform 1 0 2256 0 1 1970
box -8 -3 16 105
use FILL  FILL_6766
timestamp 1677677812
transform 1 0 2264 0 1 1970
box -8 -3 16 105
use FILL  FILL_6779
timestamp 1677677812
transform 1 0 2272 0 1 1970
box -8 -3 16 105
use FILL  FILL_6781
timestamp 1677677812
transform 1 0 2280 0 1 1970
box -8 -3 16 105
use FILL  FILL_6783
timestamp 1677677812
transform 1 0 2288 0 1 1970
box -8 -3 16 105
use FILL  FILL_6785
timestamp 1677677812
transform 1 0 2296 0 1 1970
box -8 -3 16 105
use FILL  FILL_6787
timestamp 1677677812
transform 1 0 2304 0 1 1970
box -8 -3 16 105
use FILL  FILL_6789
timestamp 1677677812
transform 1 0 2312 0 1 1970
box -8 -3 16 105
use FILL  FILL_6790
timestamp 1677677812
transform 1 0 2320 0 1 1970
box -8 -3 16 105
use FILL  FILL_6791
timestamp 1677677812
transform 1 0 2328 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_264
timestamp 1677677812
transform -1 0 2376 0 1 1970
box -8 -3 46 105
use FILL  FILL_6792
timestamp 1677677812
transform 1 0 2376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6793
timestamp 1677677812
transform 1 0 2384 0 1 1970
box -8 -3 16 105
use FILL  FILL_6794
timestamp 1677677812
transform 1 0 2392 0 1 1970
box -8 -3 16 105
use FILL  FILL_6795
timestamp 1677677812
transform 1 0 2400 0 1 1970
box -8 -3 16 105
use FILL  FILL_6796
timestamp 1677677812
transform 1 0 2408 0 1 1970
box -8 -3 16 105
use FILL  FILL_6804
timestamp 1677677812
transform 1 0 2416 0 1 1970
box -8 -3 16 105
use FILL  FILL_6806
timestamp 1677677812
transform 1 0 2424 0 1 1970
box -8 -3 16 105
use FILL  FILL_6808
timestamp 1677677812
transform 1 0 2432 0 1 1970
box -8 -3 16 105
use FILL  FILL_6810
timestamp 1677677812
transform 1 0 2440 0 1 1970
box -8 -3 16 105
use FILL  FILL_6812
timestamp 1677677812
transform 1 0 2448 0 1 1970
box -8 -3 16 105
use FILL  FILL_6813
timestamp 1677677812
transform 1 0 2456 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_426
timestamp 1677677812
transform 1 0 2464 0 1 1970
box -9 -3 26 105
use FILL  FILL_6814
timestamp 1677677812
transform 1 0 2480 0 1 1970
box -8 -3 16 105
use FILL  FILL_6816
timestamp 1677677812
transform 1 0 2488 0 1 1970
box -8 -3 16 105
use FILL  FILL_6818
timestamp 1677677812
transform 1 0 2496 0 1 1970
box -8 -3 16 105
use FILL  FILL_6820
timestamp 1677677812
transform 1 0 2504 0 1 1970
box -8 -3 16 105
use FILL  FILL_6822
timestamp 1677677812
transform 1 0 2512 0 1 1970
box -8 -3 16 105
use FILL  FILL_6824
timestamp 1677677812
transform 1 0 2520 0 1 1970
box -8 -3 16 105
use FILL  FILL_6826
timestamp 1677677812
transform 1 0 2528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6828
timestamp 1677677812
transform 1 0 2536 0 1 1970
box -8 -3 16 105
use FILL  FILL_6830
timestamp 1677677812
transform 1 0 2544 0 1 1970
box -8 -3 16 105
use FILL  FILL_6831
timestamp 1677677812
transform 1 0 2552 0 1 1970
box -8 -3 16 105
use FILL  FILL_6832
timestamp 1677677812
transform 1 0 2560 0 1 1970
box -8 -3 16 105
use FILL  FILL_6833
timestamp 1677677812
transform 1 0 2568 0 1 1970
box -8 -3 16 105
use FILL  FILL_6834
timestamp 1677677812
transform 1 0 2576 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_265
timestamp 1677677812
transform 1 0 2584 0 1 1970
box -8 -3 46 105
use FILL  FILL_6835
timestamp 1677677812
transform 1 0 2624 0 1 1970
box -8 -3 16 105
use FILL  FILL_6842
timestamp 1677677812
transform 1 0 2632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6844
timestamp 1677677812
transform 1 0 2640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6846
timestamp 1677677812
transform 1 0 2648 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_372
timestamp 1677677812
transform 1 0 2656 0 1 1970
box -8 -3 104 105
use FILL  FILL_6848
timestamp 1677677812
transform 1 0 2752 0 1 1970
box -8 -3 16 105
use FILL  FILL_6858
timestamp 1677677812
transform 1 0 2760 0 1 1970
box -8 -3 16 105
use FILL  FILL_6860
timestamp 1677677812
transform 1 0 2768 0 1 1970
box -8 -3 16 105
use FILL  FILL_6862
timestamp 1677677812
transform 1 0 2776 0 1 1970
box -8 -3 16 105
use FILL  FILL_6864
timestamp 1677677812
transform 1 0 2784 0 1 1970
box -8 -3 16 105
use FILL  FILL_6865
timestamp 1677677812
transform 1 0 2792 0 1 1970
box -8 -3 16 105
use FILL  FILL_6866
timestamp 1677677812
transform 1 0 2800 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_124
timestamp 1677677812
transform 1 0 2808 0 1 1970
box -8 -3 34 105
use FILL  FILL_6867
timestamp 1677677812
transform 1 0 2840 0 1 1970
box -8 -3 16 105
use FILL  FILL_6872
timestamp 1677677812
transform 1 0 2848 0 1 1970
box -8 -3 16 105
use FILL  FILL_6874
timestamp 1677677812
transform 1 0 2856 0 1 1970
box -8 -3 16 105
use FILL  FILL_6876
timestamp 1677677812
transform 1 0 2864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6878
timestamp 1677677812
transform 1 0 2872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6880
timestamp 1677677812
transform 1 0 2880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6882
timestamp 1677677812
transform 1 0 2888 0 1 1970
box -8 -3 16 105
use FILL  FILL_6883
timestamp 1677677812
transform 1 0 2896 0 1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_126
timestamp 1677677812
transform -1 0 2936 0 1 1970
box -8 -3 34 105
use FILL  FILL_6884
timestamp 1677677812
transform 1 0 2936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6888
timestamp 1677677812
transform 1 0 2944 0 1 1970
box -8 -3 16 105
use FILL  FILL_6890
timestamp 1677677812
transform 1 0 2952 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_25
timestamp 1677677812
transform 1 0 2960 0 1 1970
box -8 -3 40 105
use FILL  FILL_6892
timestamp 1677677812
transform 1 0 2992 0 1 1970
box -8 -3 16 105
use FILL  FILL_6893
timestamp 1677677812
transform 1 0 3000 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5124
timestamp 1677677812
transform 1 0 3044 0 1 1975
box -3 -3 3 3
use OAI22X1  OAI22X1_253
timestamp 1677677812
transform -1 0 3048 0 1 1970
box -8 -3 46 105
use FILL  FILL_6894
timestamp 1677677812
transform 1 0 3048 0 1 1970
box -8 -3 16 105
use FILL  FILL_6895
timestamp 1677677812
transform 1 0 3056 0 1 1970
box -8 -3 16 105
use FILL  FILL_6896
timestamp 1677677812
transform 1 0 3064 0 1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5125
timestamp 1677677812
transform 1 0 3148 0 1 1975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_373
timestamp 1677677812
transform -1 0 3168 0 1 1970
box -8 -3 104 105
use FILL  FILL_6897
timestamp 1677677812
transform 1 0 3168 0 1 1970
box -8 -3 16 105
use FILL  FILL_6913
timestamp 1677677812
transform 1 0 3176 0 1 1970
box -8 -3 16 105
use FILL  FILL_6914
timestamp 1677677812
transform 1 0 3184 0 1 1970
box -8 -3 16 105
use BUFX2  BUFX2_85
timestamp 1677677812
transform -1 0 3216 0 1 1970
box -5 -3 28 105
use FILL  FILL_6915
timestamp 1677677812
transform 1 0 3216 0 1 1970
box -8 -3 16 105
use FILL  FILL_6916
timestamp 1677677812
transform 1 0 3224 0 1 1970
box -8 -3 16 105
use FILL  FILL_6917
timestamp 1677677812
transform 1 0 3232 0 1 1970
box -8 -3 16 105
use FILL  FILL_6918
timestamp 1677677812
transform 1 0 3240 0 1 1970
box -8 -3 16 105
use FILL  FILL_6919
timestamp 1677677812
transform 1 0 3248 0 1 1970
box -8 -3 16 105
use FILL  FILL_6920
timestamp 1677677812
transform 1 0 3256 0 1 1970
box -8 -3 16 105
use FILL  FILL_6921
timestamp 1677677812
transform 1 0 3264 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_44
timestamp 1677677812
transform -1 0 3304 0 1 1970
box -8 -3 40 105
use M3_M2  M3_M2_5126
timestamp 1677677812
transform 1 0 3316 0 1 1975
box -3 -3 3 3
use FILL  FILL_6922
timestamp 1677677812
transform 1 0 3304 0 1 1970
box -8 -3 16 105
use FILL  FILL_6923
timestamp 1677677812
transform 1 0 3312 0 1 1970
box -8 -3 16 105
use FILL  FILL_6924
timestamp 1677677812
transform 1 0 3320 0 1 1970
box -8 -3 16 105
use FILL  FILL_6925
timestamp 1677677812
transform 1 0 3328 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_26
timestamp 1677677812
transform 1 0 3336 0 1 1970
box -8 -3 40 105
use FILL  FILL_6926
timestamp 1677677812
transform 1 0 3368 0 1 1970
box -8 -3 16 105
use FILL  FILL_6937
timestamp 1677677812
transform 1 0 3376 0 1 1970
box -8 -3 16 105
use FILL  FILL_6938
timestamp 1677677812
transform 1 0 3384 0 1 1970
box -8 -3 16 105
use FILL  FILL_6939
timestamp 1677677812
transform 1 0 3392 0 1 1970
box -8 -3 16 105
use FILL  FILL_6941
timestamp 1677677812
transform 1 0 3400 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_254
timestamp 1677677812
transform -1 0 3448 0 1 1970
box -8 -3 46 105
use FILL  FILL_6942
timestamp 1677677812
transform 1 0 3448 0 1 1970
box -8 -3 16 105
use FILL  FILL_6950
timestamp 1677677812
transform 1 0 3456 0 1 1970
box -8 -3 16 105
use FILL  FILL_6952
timestamp 1677677812
transform 1 0 3464 0 1 1970
box -8 -3 16 105
use FILL  FILL_6954
timestamp 1677677812
transform 1 0 3472 0 1 1970
box -8 -3 16 105
use FILL  FILL_6956
timestamp 1677677812
transform 1 0 3480 0 1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_46
timestamp 1677677812
transform -1 0 3520 0 1 1970
box -8 -3 40 105
use FILL  FILL_6957
timestamp 1677677812
transform 1 0 3520 0 1 1970
box -8 -3 16 105
use FILL  FILL_6958
timestamp 1677677812
transform 1 0 3528 0 1 1970
box -8 -3 16 105
use FILL  FILL_6961
timestamp 1677677812
transform 1 0 3536 0 1 1970
box -8 -3 16 105
use FILL  FILL_6963
timestamp 1677677812
transform 1 0 3544 0 1 1970
box -8 -3 16 105
use FILL  FILL_6965
timestamp 1677677812
transform 1 0 3552 0 1 1970
box -8 -3 16 105
use FILL  FILL_6967
timestamp 1677677812
transform 1 0 3560 0 1 1970
box -8 -3 16 105
use FILL  FILL_6969
timestamp 1677677812
transform 1 0 3568 0 1 1970
box -8 -3 16 105
use FILL  FILL_6971
timestamp 1677677812
transform 1 0 3576 0 1 1970
box -8 -3 16 105
use FILL  FILL_6972
timestamp 1677677812
transform 1 0 3584 0 1 1970
box -8 -3 16 105
use FILL  FILL_6973
timestamp 1677677812
transform 1 0 3592 0 1 1970
box -8 -3 16 105
use FILL  FILL_6975
timestamp 1677677812
transform 1 0 3600 0 1 1970
box -8 -3 16 105
use FILL  FILL_6977
timestamp 1677677812
transform 1 0 3608 0 1 1970
box -8 -3 16 105
use FILL  FILL_6978
timestamp 1677677812
transform 1 0 3616 0 1 1970
box -8 -3 16 105
use FILL  FILL_6979
timestamp 1677677812
transform 1 0 3624 0 1 1970
box -8 -3 16 105
use FILL  FILL_6980
timestamp 1677677812
transform 1 0 3632 0 1 1970
box -8 -3 16 105
use FILL  FILL_6981
timestamp 1677677812
transform 1 0 3640 0 1 1970
box -8 -3 16 105
use FILL  FILL_6982
timestamp 1677677812
transform 1 0 3648 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_27
timestamp 1677677812
transform 1 0 3656 0 1 1970
box -8 -3 40 105
use FILL  FILL_6983
timestamp 1677677812
transform 1 0 3688 0 1 1970
box -8 -3 16 105
use FILL  FILL_6984
timestamp 1677677812
transform 1 0 3696 0 1 1970
box -8 -3 16 105
use FILL  FILL_6985
timestamp 1677677812
transform 1 0 3704 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_374
timestamp 1677677812
transform 1 0 3712 0 1 1970
box -8 -3 104 105
use FILL  FILL_6986
timestamp 1677677812
transform 1 0 3808 0 1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_255
timestamp 1677677812
transform -1 0 3856 0 1 1970
box -8 -3 46 105
use FILL  FILL_6987
timestamp 1677677812
transform 1 0 3856 0 1 1970
box -8 -3 16 105
use FILL  FILL_6988
timestamp 1677677812
transform 1 0 3864 0 1 1970
box -8 -3 16 105
use FILL  FILL_6989
timestamp 1677677812
transform 1 0 3872 0 1 1970
box -8 -3 16 105
use FILL  FILL_6990
timestamp 1677677812
transform 1 0 3880 0 1 1970
box -8 -3 16 105
use FILL  FILL_6991
timestamp 1677677812
transform 1 0 3888 0 1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_269
timestamp 1677677812
transform 1 0 3896 0 1 1970
box -8 -3 46 105
use FILL  FILL_6992
timestamp 1677677812
transform 1 0 3936 0 1 1970
box -8 -3 16 105
use FILL  FILL_6993
timestamp 1677677812
transform 1 0 3944 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_375
timestamp 1677677812
transform 1 0 3952 0 1 1970
box -8 -3 104 105
use OAI22X1  OAI22X1_256
timestamp 1677677812
transform 1 0 4048 0 1 1970
box -8 -3 46 105
use FILL  FILL_6994
timestamp 1677677812
transform 1 0 4088 0 1 1970
box -8 -3 16 105
use FILL  FILL_6995
timestamp 1677677812
transform 1 0 4096 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_430
timestamp 1677677812
transform -1 0 4120 0 1 1970
box -9 -3 26 105
use FILL  FILL_6996
timestamp 1677677812
transform 1 0 4120 0 1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_376
timestamp 1677677812
transform -1 0 4224 0 1 1970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_377
timestamp 1677677812
transform 1 0 4224 0 1 1970
box -8 -3 104 105
use INVX2  INVX2_431
timestamp 1677677812
transform 1 0 4320 0 1 1970
box -9 -3 26 105
use AND2X2  AND2X2_28
timestamp 1677677812
transform -1 0 4368 0 1 1970
box -8 -3 40 105
use FILL  FILL_6997
timestamp 1677677812
transform 1 0 4368 0 1 1970
box -8 -3 16 105
use FILL  FILL_7023
timestamp 1677677812
transform 1 0 4376 0 1 1970
box -8 -3 16 105
use FILL  FILL_7024
timestamp 1677677812
transform 1 0 4384 0 1 1970
box -8 -3 16 105
use FILL  FILL_7025
timestamp 1677677812
transform 1 0 4392 0 1 1970
box -8 -3 16 105
use FILL  FILL_7026
timestamp 1677677812
transform 1 0 4400 0 1 1970
box -8 -3 16 105
use FILL  FILL_7027
timestamp 1677677812
transform 1 0 4408 0 1 1970
box -8 -3 16 105
use FILL  FILL_7028
timestamp 1677677812
transform 1 0 4416 0 1 1970
box -8 -3 16 105
use FILL  FILL_7029
timestamp 1677677812
transform 1 0 4424 0 1 1970
box -8 -3 16 105
use FILL  FILL_7030
timestamp 1677677812
transform 1 0 4432 0 1 1970
box -8 -3 16 105
use FILL  FILL_7031
timestamp 1677677812
transform 1 0 4440 0 1 1970
box -8 -3 16 105
use AND2X2  AND2X2_29
timestamp 1677677812
transform 1 0 4448 0 1 1970
box -8 -3 40 105
use FILL  FILL_7032
timestamp 1677677812
transform 1 0 4480 0 1 1970
box -8 -3 16 105
use FILL  FILL_7033
timestamp 1677677812
transform 1 0 4488 0 1 1970
box -8 -3 16 105
use FILL  FILL_7035
timestamp 1677677812
transform 1 0 4496 0 1 1970
box -8 -3 16 105
use FILL  FILL_7036
timestamp 1677677812
transform 1 0 4504 0 1 1970
box -8 -3 16 105
use FILL  FILL_7037
timestamp 1677677812
transform 1 0 4512 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_436
timestamp 1677677812
transform 1 0 4520 0 1 1970
box -9 -3 26 105
use FILL  FILL_7038
timestamp 1677677812
transform 1 0 4536 0 1 1970
box -8 -3 16 105
use FILL  FILL_7039
timestamp 1677677812
transform 1 0 4544 0 1 1970
box -8 -3 16 105
use FILL  FILL_7040
timestamp 1677677812
transform 1 0 4552 0 1 1970
box -8 -3 16 105
use FILL  FILL_7041
timestamp 1677677812
transform 1 0 4560 0 1 1970
box -8 -3 16 105
use FILL  FILL_7042
timestamp 1677677812
transform 1 0 4568 0 1 1970
box -8 -3 16 105
use FILL  FILL_7043
timestamp 1677677812
transform 1 0 4576 0 1 1970
box -8 -3 16 105
use FILL  FILL_7044
timestamp 1677677812
transform 1 0 4584 0 1 1970
box -8 -3 16 105
use FILL  FILL_7045
timestamp 1677677812
transform 1 0 4592 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_437
timestamp 1677677812
transform -1 0 4616 0 1 1970
box -9 -3 26 105
use FILL  FILL_7046
timestamp 1677677812
transform 1 0 4616 0 1 1970
box -8 -3 16 105
use FILL  FILL_7049
timestamp 1677677812
transform 1 0 4624 0 1 1970
box -8 -3 16 105
use FILL  FILL_7050
timestamp 1677677812
transform 1 0 4632 0 1 1970
box -8 -3 16 105
use INVX2  INVX2_439
timestamp 1677677812
transform -1 0 4656 0 1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_385
timestamp 1677677812
transform 1 0 4656 0 1 1970
box -8 -3 104 105
use FILL  FILL_7051
timestamp 1677677812
transform 1 0 4752 0 1 1970
box -8 -3 16 105
use FILL  FILL_7057
timestamp 1677677812
transform 1 0 4760 0 1 1970
box -8 -3 16 105
use FILL  FILL_7059
timestamp 1677677812
transform 1 0 4768 0 1 1970
box -8 -3 16 105
use FILL  FILL_7061
timestamp 1677677812
transform 1 0 4776 0 1 1970
box -8 -3 16 105
use FILL  FILL_7063
timestamp 1677677812
transform 1 0 4784 0 1 1970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_55
timestamp 1677677812
transform 1 0 4819 0 1 1970
box -10 -3 10 3
use M2_M1  M2_M1_5733
timestamp 1677677812
transform 1 0 68 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5734
timestamp 1677677812
transform 1 0 84 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5802
timestamp 1677677812
transform 1 0 100 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5150
timestamp 1677677812
transform 1 0 124 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5151
timestamp 1677677812
transform 1 0 156 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5177
timestamp 1677677812
transform 1 0 140 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5735
timestamp 1677677812
transform 1 0 156 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5127
timestamp 1677677812
transform 1 0 340 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5128
timestamp 1677677812
transform 1 0 356 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5152
timestamp 1677677812
transform 1 0 268 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5736
timestamp 1677677812
transform 1 0 268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5737
timestamp 1677677812
transform 1 0 356 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5738
timestamp 1677677812
transform 1 0 380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5739
timestamp 1677677812
transform 1 0 468 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5803
timestamp 1677677812
transform 1 0 140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5804
timestamp 1677677812
transform 1 0 196 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5805
timestamp 1677677812
transform 1 0 236 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5806
timestamp 1677677812
transform 1 0 244 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5807
timestamp 1677677812
transform 1 0 252 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5808
timestamp 1677677812
transform 1 0 300 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5809
timestamp 1677677812
transform 1 0 348 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5810
timestamp 1677677812
transform 1 0 364 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5811
timestamp 1677677812
transform 1 0 404 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5812
timestamp 1677677812
transform 1 0 460 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5200
timestamp 1677677812
transform 1 0 364 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5201
timestamp 1677677812
transform 1 0 404 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5202
timestamp 1677677812
transform 1 0 460 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5226
timestamp 1677677812
transform 1 0 356 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5234
timestamp 1677677812
transform 1 0 268 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5227
timestamp 1677677812
transform 1 0 404 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5235
timestamp 1677677812
transform 1 0 468 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5142
timestamp 1677677812
transform 1 0 500 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5740
timestamp 1677677812
transform 1 0 500 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5741
timestamp 1677677812
transform 1 0 516 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5742
timestamp 1677677812
transform 1 0 524 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5813
timestamp 1677677812
transform 1 0 492 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5203
timestamp 1677677812
transform 1 0 516 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5814
timestamp 1677677812
transform 1 0 532 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5228
timestamp 1677677812
transform 1 0 532 0 1 1905
box -3 -3 3 3
use M3_M2  M3_M2_5178
timestamp 1677677812
transform 1 0 580 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5815
timestamp 1677677812
transform 1 0 556 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5816
timestamp 1677677812
transform 1 0 564 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5817
timestamp 1677677812
transform 1 0 580 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5204
timestamp 1677677812
transform 1 0 580 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5143
timestamp 1677677812
transform 1 0 596 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5729
timestamp 1677677812
transform 1 0 596 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5743
timestamp 1677677812
transform 1 0 620 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5205
timestamp 1677677812
transform 1 0 644 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5744
timestamp 1677677812
transform 1 0 668 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5229
timestamp 1677677812
transform 1 0 668 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5730
timestamp 1677677812
transform 1 0 700 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5818
timestamp 1677677812
transform 1 0 692 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5206
timestamp 1677677812
transform 1 0 692 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5745
timestamp 1677677812
transform 1 0 708 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5179
timestamp 1677677812
transform 1 0 724 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5819
timestamp 1677677812
transform 1 0 724 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5236
timestamp 1677677812
transform 1 0 724 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5248
timestamp 1677677812
transform 1 0 724 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5820
timestamp 1677677812
transform 1 0 740 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5249
timestamp 1677677812
transform 1 0 740 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5153
timestamp 1677677812
transform 1 0 788 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5746
timestamp 1677677812
transform 1 0 788 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5821
timestamp 1677677812
transform 1 0 796 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5129
timestamp 1677677812
transform 1 0 836 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5747
timestamp 1677677812
transform 1 0 828 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5748
timestamp 1677677812
transform 1 0 836 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5822
timestamp 1677677812
transform 1 0 860 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5823
timestamp 1677677812
transform 1 0 964 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5250
timestamp 1677677812
transform 1 0 988 0 1 1885
box -3 -3 3 3
use M2_M1  M2_M1_5749
timestamp 1677677812
transform 1 0 1028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5750
timestamp 1677677812
transform 1 0 1052 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5824
timestamp 1677677812
transform 1 0 1036 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5230
timestamp 1677677812
transform 1 0 1036 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5825
timestamp 1677677812
transform 1 0 1084 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5751
timestamp 1677677812
transform 1 0 1124 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5826
timestamp 1677677812
transform 1 0 1140 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5827
timestamp 1677677812
transform 1 0 1172 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5752
timestamp 1677677812
transform 1 0 1212 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5828
timestamp 1677677812
transform 1 0 1244 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5180
timestamp 1677677812
transform 1 0 1268 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5753
timestamp 1677677812
transform 1 0 1332 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5829
timestamp 1677677812
transform 1 0 1364 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5237
timestamp 1677677812
transform 1 0 1324 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5830
timestamp 1677677812
transform 1 0 1420 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5831
timestamp 1677677812
transform 1 0 1436 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5154
timestamp 1677677812
transform 1 0 1500 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5754
timestamp 1677677812
transform 1 0 1484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5755
timestamp 1677677812
transform 1 0 1492 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5832
timestamp 1677677812
transform 1 0 1476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5833
timestamp 1677677812
transform 1 0 1508 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5238
timestamp 1677677812
transform 1 0 1524 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5239
timestamp 1677677812
transform 1 0 1548 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5756
timestamp 1677677812
transform 1 0 1580 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5130
timestamp 1677677812
transform 1 0 1596 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5834
timestamp 1677677812
transform 1 0 1620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5757
timestamp 1677677812
transform 1 0 1644 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5758
timestamp 1677677812
transform 1 0 1676 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5759
timestamp 1677677812
transform 1 0 1684 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5187
timestamp 1677677812
transform 1 0 1676 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5144
timestamp 1677677812
transform 1 0 1724 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5155
timestamp 1677677812
transform 1 0 1724 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5835
timestamp 1677677812
transform 1 0 1724 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5836
timestamp 1677677812
transform 1 0 1732 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5207
timestamp 1677677812
transform 1 0 1724 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5760
timestamp 1677677812
transform 1 0 1748 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5156
timestamp 1677677812
transform 1 0 1812 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5761
timestamp 1677677812
transform 1 0 1804 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5762
timestamp 1677677812
transform 1 0 1812 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5208
timestamp 1677677812
transform 1 0 1804 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5240
timestamp 1677677812
transform 1 0 1828 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5837
timestamp 1677677812
transform 1 0 1844 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5209
timestamp 1677677812
transform 1 0 1844 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5188
timestamp 1677677812
transform 1 0 1884 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5131
timestamp 1677677812
transform 1 0 1900 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5763
timestamp 1677677812
transform 1 0 1900 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5764
timestamp 1677677812
transform 1 0 1916 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5145
timestamp 1677677812
transform 1 0 1980 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5838
timestamp 1677677812
transform 1 0 1948 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5839
timestamp 1677677812
transform 1 0 1956 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5840
timestamp 1677677812
transform 1 0 1972 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5841
timestamp 1677677812
transform 1 0 1988 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5210
timestamp 1677677812
transform 1 0 1948 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5189
timestamp 1677677812
transform 1 0 1996 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5157
timestamp 1677677812
transform 1 0 2012 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5765
timestamp 1677677812
transform 1 0 2012 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5132
timestamp 1677677812
transform 1 0 2044 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5158
timestamp 1677677812
transform 1 0 2052 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5766
timestamp 1677677812
transform 1 0 2100 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5842
timestamp 1677677812
transform 1 0 2020 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5843
timestamp 1677677812
transform 1 0 2052 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5190
timestamp 1677677812
transform 1 0 2100 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5211
timestamp 1677677812
transform 1 0 2052 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5191
timestamp 1677677812
transform 1 0 2164 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5241
timestamp 1677677812
transform 1 0 2164 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5159
timestamp 1677677812
transform 1 0 2188 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5146
timestamp 1677677812
transform 1 0 2212 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5133
timestamp 1677677812
transform 1 0 2244 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5767
timestamp 1677677812
transform 1 0 2244 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5147
timestamp 1677677812
transform 1 0 2268 0 1 1955
box -3 -3 3 3
use M2_M1  M2_M1_5844
timestamp 1677677812
transform 1 0 2260 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5845
timestamp 1677677812
transform 1 0 2268 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5768
timestamp 1677677812
transform 1 0 2356 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5134
timestamp 1677677812
transform 1 0 2372 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5769
timestamp 1677677812
transform 1 0 2380 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5846
timestamp 1677677812
transform 1 0 2388 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5212
timestamp 1677677812
transform 1 0 2388 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5770
timestamp 1677677812
transform 1 0 2412 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5847
timestamp 1677677812
transform 1 0 2444 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5848
timestamp 1677677812
transform 1 0 2460 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5849
timestamp 1677677812
transform 1 0 2476 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5850
timestamp 1677677812
transform 1 0 2484 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5213
timestamp 1677677812
transform 1 0 2468 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5214
timestamp 1677677812
transform 1 0 2484 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5192
timestamp 1677677812
transform 1 0 2524 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5771
timestamp 1677677812
transform 1 0 2556 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5772
timestamp 1677677812
transform 1 0 2572 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5851
timestamp 1677677812
transform 1 0 2564 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5193
timestamp 1677677812
transform 1 0 2572 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5852
timestamp 1677677812
transform 1 0 2620 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5853
timestamp 1677677812
transform 1 0 2636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5773
timestamp 1677677812
transform 1 0 2732 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5774
timestamp 1677677812
transform 1 0 2740 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5854
timestamp 1677677812
transform 1 0 2724 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5194
timestamp 1677677812
transform 1 0 2740 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5215
timestamp 1677677812
transform 1 0 2732 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5135
timestamp 1677677812
transform 1 0 2796 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5855
timestamp 1677677812
transform 1 0 2796 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5136
timestamp 1677677812
transform 1 0 2820 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5775
timestamp 1677677812
transform 1 0 2820 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5216
timestamp 1677677812
transform 1 0 2820 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5160
timestamp 1677677812
transform 1 0 2924 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5731
timestamp 1677677812
transform 1 0 2932 0 1 1945
box -2 -2 2 2
use M2_M1  M2_M1_5856
timestamp 1677677812
transform 1 0 2916 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5894
timestamp 1677677812
transform 1 0 2900 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5137
timestamp 1677677812
transform 1 0 2972 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5776
timestamp 1677677812
transform 1 0 2972 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5138
timestamp 1677677812
transform 1 0 3020 0 1 1965
box -3 -3 3 3
use M2_M1  M2_M1_5777
timestamp 1677677812
transform 1 0 3012 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5857
timestamp 1677677812
transform 1 0 2996 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5858
timestamp 1677677812
transform 1 0 3004 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5217
timestamp 1677677812
transform 1 0 2996 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5195
timestamp 1677677812
transform 1 0 3012 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5139
timestamp 1677677812
transform 1 0 3052 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5161
timestamp 1677677812
transform 1 0 3044 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5778
timestamp 1677677812
transform 1 0 3044 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5859
timestamp 1677677812
transform 1 0 3052 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5779
timestamp 1677677812
transform 1 0 3076 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5895
timestamp 1677677812
transform 1 0 3076 0 1 1915
box -2 -2 2 2
use M3_M2  M3_M2_5242
timestamp 1677677812
transform 1 0 3084 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5860
timestamp 1677677812
transform 1 0 3140 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5231
timestamp 1677677812
transform 1 0 3124 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5896
timestamp 1677677812
transform 1 0 3148 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5898
timestamp 1677677812
transform 1 0 3132 0 1 1905
box -2 -2 2 2
use M2_M1  M2_M1_5899
timestamp 1677677812
transform 1 0 3140 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5243
timestamp 1677677812
transform 1 0 3148 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5251
timestamp 1677677812
transform 1 0 3132 0 1 1885
box -3 -3 3 3
use M3_M2  M3_M2_5196
timestamp 1677677812
transform 1 0 3196 0 1 1925
box -3 -3 3 3
use M3_M2  M3_M2_5162
timestamp 1677677812
transform 1 0 3244 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5780
timestamp 1677677812
transform 1 0 3236 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5861
timestamp 1677677812
transform 1 0 3204 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5862
timestamp 1677677812
transform 1 0 3220 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5218
timestamp 1677677812
transform 1 0 3204 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5897
timestamp 1677677812
transform 1 0 3212 0 1 1915
box -2 -2 2 2
use M2_M1  M2_M1_5900
timestamp 1677677812
transform 1 0 3196 0 1 1905
box -2 -2 2 2
use M3_M2  M3_M2_5232
timestamp 1677677812
transform 1 0 3212 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5863
timestamp 1677677812
transform 1 0 3244 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5163
timestamp 1677677812
transform 1 0 3276 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5781
timestamp 1677677812
transform 1 0 3268 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5864
timestamp 1677677812
transform 1 0 3276 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5782
timestamp 1677677812
transform 1 0 3308 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5197
timestamp 1677677812
transform 1 0 3308 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5865
timestamp 1677677812
transform 1 0 3316 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5866
timestamp 1677677812
transform 1 0 3332 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5219
timestamp 1677677812
transform 1 0 3316 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5244
timestamp 1677677812
transform 1 0 3332 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5783
timestamp 1677677812
transform 1 0 3372 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5784
timestamp 1677677812
transform 1 0 3420 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5867
timestamp 1677677812
transform 1 0 3484 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5785
timestamp 1677677812
transform 1 0 3500 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5786
timestamp 1677677812
transform 1 0 3524 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5198
timestamp 1677677812
transform 1 0 3500 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5868
timestamp 1677677812
transform 1 0 3508 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5869
timestamp 1677677812
transform 1 0 3524 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5245
timestamp 1677677812
transform 1 0 3524 0 1 1895
box -3 -3 3 3
use M3_M2  M3_M2_5246
timestamp 1677677812
transform 1 0 3548 0 1 1895
box -3 -3 3 3
use M2_M1  M2_M1_5787
timestamp 1677677812
transform 1 0 3580 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5181
timestamp 1677677812
transform 1 0 3596 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5199
timestamp 1677677812
transform 1 0 3588 0 1 1925
box -3 -3 3 3
use M2_M1  M2_M1_5870
timestamp 1677677812
transform 1 0 3612 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5164
timestamp 1677677812
transform 1 0 3700 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5182
timestamp 1677677812
transform 1 0 3652 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5788
timestamp 1677677812
transform 1 0 3700 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5871
timestamp 1677677812
transform 1 0 3652 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5220
timestamp 1677677812
transform 1 0 3676 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5165
timestamp 1677677812
transform 1 0 3724 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5872
timestamp 1677677812
transform 1 0 3716 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5221
timestamp 1677677812
transform 1 0 3716 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5183
timestamp 1677677812
transform 1 0 3748 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5873
timestamp 1677677812
transform 1 0 3748 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5140
timestamp 1677677812
transform 1 0 3812 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5148
timestamp 1677677812
transform 1 0 3788 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5166
timestamp 1677677812
transform 1 0 3780 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5167
timestamp 1677677812
transform 1 0 3804 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5789
timestamp 1677677812
transform 1 0 3780 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5790
timestamp 1677677812
transform 1 0 3788 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5184
timestamp 1677677812
transform 1 0 3796 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5168
timestamp 1677677812
transform 1 0 3820 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5874
timestamp 1677677812
transform 1 0 3796 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5875
timestamp 1677677812
transform 1 0 3812 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5233
timestamp 1677677812
transform 1 0 3796 0 1 1905
box -3 -3 3 3
use M2_M1  M2_M1_5791
timestamp 1677677812
transform 1 0 3828 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5185
timestamp 1677677812
transform 1 0 3836 0 1 1935
box -3 -3 3 3
use M3_M2  M3_M2_5141
timestamp 1677677812
transform 1 0 3932 0 1 1965
box -3 -3 3 3
use M3_M2  M3_M2_5169
timestamp 1677677812
transform 1 0 3852 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5792
timestamp 1677677812
transform 1 0 3852 0 1 1935
box -2 -2 2 2
use M3_M2  M3_M2_5186
timestamp 1677677812
transform 1 0 3876 0 1 1935
box -3 -3 3 3
use M2_M1  M2_M1_5876
timestamp 1677677812
transform 1 0 3876 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5877
timestamp 1677677812
transform 1 0 3932 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5878
timestamp 1677677812
transform 1 0 3940 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5170
timestamp 1677677812
transform 1 0 3964 0 1 1945
box -3 -3 3 3
use M3_M2  M3_M2_5171
timestamp 1677677812
transform 1 0 4028 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5793
timestamp 1677677812
transform 1 0 4028 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5879
timestamp 1677677812
transform 1 0 3980 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5149
timestamp 1677677812
transform 1 0 4060 0 1 1955
box -3 -3 3 3
use M3_M2  M3_M2_5172
timestamp 1677677812
transform 1 0 4076 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5794
timestamp 1677677812
transform 1 0 4076 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5795
timestamp 1677677812
transform 1 0 4172 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5880
timestamp 1677677812
transform 1 0 4124 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5881
timestamp 1677677812
transform 1 0 4156 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5882
timestamp 1677677812
transform 1 0 4164 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5222
timestamp 1677677812
transform 1 0 4124 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5223
timestamp 1677677812
transform 1 0 4172 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5173
timestamp 1677677812
transform 1 0 4204 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5796
timestamp 1677677812
transform 1 0 4204 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5883
timestamp 1677677812
transform 1 0 4236 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5884
timestamp 1677677812
transform 1 0 4284 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5885
timestamp 1677677812
transform 1 0 4308 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5174
timestamp 1677677812
transform 1 0 4324 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5732
timestamp 1677677812
transform 1 0 4340 0 1 1945
box -2 -2 2 2
use M3_M2  M3_M2_5175
timestamp 1677677812
transform 1 0 4388 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5797
timestamp 1677677812
transform 1 0 4388 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5798
timestamp 1677677812
transform 1 0 4484 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5886
timestamp 1677677812
transform 1 0 4436 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5887
timestamp 1677677812
transform 1 0 4468 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5888
timestamp 1677677812
transform 1 0 4476 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5176
timestamp 1677677812
transform 1 0 4508 0 1 1945
box -3 -3 3 3
use M2_M1  M2_M1_5799
timestamp 1677677812
transform 1 0 4508 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5800
timestamp 1677677812
transform 1 0 4604 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5889
timestamp 1677677812
transform 1 0 4532 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5890
timestamp 1677677812
transform 1 0 4588 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5891
timestamp 1677677812
transform 1 0 4596 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5224
timestamp 1677677812
transform 1 0 4508 0 1 1915
box -3 -3 3 3
use M3_M2  M3_M2_5225
timestamp 1677677812
transform 1 0 4532 0 1 1915
box -3 -3 3 3
use M2_M1  M2_M1_5801
timestamp 1677677812
transform 1 0 4716 0 1 1935
box -2 -2 2 2
use M2_M1  M2_M1_5892
timestamp 1677677812
transform 1 0 4636 0 1 1925
box -2 -2 2 2
use M2_M1  M2_M1_5893
timestamp 1677677812
transform 1 0 4668 0 1 1925
box -2 -2 2 2
use M3_M2  M3_M2_5247
timestamp 1677677812
transform 1 0 4740 0 1 1895
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_56
timestamp 1677677812
transform 1 0 24 0 1 1870
box -10 -3 10 3
use FILL  FILL_6505
timestamp 1677677812
transform 1 0 72 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_66
timestamp 1677677812
transform -1 0 104 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6506
timestamp 1677677812
transform 1 0 104 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_67
timestamp 1677677812
transform -1 0 136 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6507
timestamp 1677677812
transform 1 0 136 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_365
timestamp 1677677812
transform 1 0 144 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_417
timestamp 1677677812
transform -1 0 256 0 -1 1970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_366
timestamp 1677677812
transform 1 0 256 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_418
timestamp 1677677812
transform 1 0 352 0 -1 1970
box -9 -3 26 105
use M3_M2  M3_M2_5252
timestamp 1677677812
transform 1 0 396 0 1 1875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_367
timestamp 1677677812
transform 1 0 368 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6508
timestamp 1677677812
transform 1 0 464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6509
timestamp 1677677812
transform 1 0 472 0 -1 1970
box -8 -3 16 105
use OAI22X1  OAI22X1_252
timestamp 1677677812
transform -1 0 520 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6510
timestamp 1677677812
transform 1 0 520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6511
timestamp 1677677812
transform 1 0 528 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5253
timestamp 1677677812
transform 1 0 564 0 1 1875
box -3 -3 3 3
use BUFX2  BUFX2_68
timestamp 1677677812
transform -1 0 560 0 -1 1970
box -5 -3 28 105
use M3_M2  M3_M2_5254
timestamp 1677677812
transform 1 0 588 0 1 1875
box -3 -3 3 3
use AND2X2  AND2X2_20
timestamp 1677677812
transform -1 0 592 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6512
timestamp 1677677812
transform 1 0 592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6513
timestamp 1677677812
transform 1 0 600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6514
timestamp 1677677812
transform 1 0 608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6515
timestamp 1677677812
transform 1 0 616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6517
timestamp 1677677812
transform 1 0 624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6519
timestamp 1677677812
transform 1 0 632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6521
timestamp 1677677812
transform 1 0 640 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_60
timestamp 1677677812
transform 1 0 648 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6530
timestamp 1677677812
transform 1 0 672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6531
timestamp 1677677812
transform 1 0 680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6532
timestamp 1677677812
transform 1 0 688 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_61
timestamp 1677677812
transform 1 0 696 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6533
timestamp 1677677812
transform 1 0 720 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_419
timestamp 1677677812
transform -1 0 744 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6534
timestamp 1677677812
transform 1 0 744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6536
timestamp 1677677812
transform 1 0 752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6538
timestamp 1677677812
transform 1 0 760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6539
timestamp 1677677812
transform 1 0 768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6540
timestamp 1677677812
transform 1 0 776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6541
timestamp 1677677812
transform 1 0 784 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_420
timestamp 1677677812
transform -1 0 808 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6542
timestamp 1677677812
transform 1 0 808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6543
timestamp 1677677812
transform 1 0 816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6544
timestamp 1677677812
transform 1 0 824 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_69
timestamp 1677677812
transform -1 0 856 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6545
timestamp 1677677812
transform 1 0 856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6547
timestamp 1677677812
transform 1 0 864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6549
timestamp 1677677812
transform 1 0 872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6551
timestamp 1677677812
transform 1 0 880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6553
timestamp 1677677812
transform 1 0 888 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6555
timestamp 1677677812
transform 1 0 896 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6557
timestamp 1677677812
transform 1 0 904 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6559
timestamp 1677677812
transform 1 0 912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6561
timestamp 1677677812
transform 1 0 920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6563
timestamp 1677677812
transform 1 0 928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6565
timestamp 1677677812
transform 1 0 936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6567
timestamp 1677677812
transform 1 0 944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6569
timestamp 1677677812
transform 1 0 952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6570
timestamp 1677677812
transform 1 0 960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6571
timestamp 1677677812
transform 1 0 968 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6572
timestamp 1677677812
transform 1 0 976 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6574
timestamp 1677677812
transform 1 0 984 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6576
timestamp 1677677812
transform 1 0 992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6582
timestamp 1677677812
transform 1 0 1000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6583
timestamp 1677677812
transform 1 0 1008 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_260
timestamp 1677677812
transform 1 0 1016 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6584
timestamp 1677677812
transform 1 0 1056 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6586
timestamp 1677677812
transform 1 0 1064 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6588
timestamp 1677677812
transform 1 0 1072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6589
timestamp 1677677812
transform 1 0 1080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6590
timestamp 1677677812
transform 1 0 1088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6591
timestamp 1677677812
transform 1 0 1096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6593
timestamp 1677677812
transform 1 0 1104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6595
timestamp 1677677812
transform 1 0 1112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6597
timestamp 1677677812
transform 1 0 1120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6599
timestamp 1677677812
transform 1 0 1128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6601
timestamp 1677677812
transform 1 0 1136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6606
timestamp 1677677812
transform 1 0 1144 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_261
timestamp 1677677812
transform 1 0 1152 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6607
timestamp 1677677812
transform 1 0 1192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6609
timestamp 1677677812
transform 1 0 1200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6611
timestamp 1677677812
transform 1 0 1208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6613
timestamp 1677677812
transform 1 0 1216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6615
timestamp 1677677812
transform 1 0 1224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6617
timestamp 1677677812
transform 1 0 1232 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6619
timestamp 1677677812
transform 1 0 1240 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6621
timestamp 1677677812
transform 1 0 1248 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6623
timestamp 1677677812
transform 1 0 1256 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6625
timestamp 1677677812
transform 1 0 1264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6627
timestamp 1677677812
transform 1 0 1272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6628
timestamp 1677677812
transform 1 0 1280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6629
timestamp 1677677812
transform 1 0 1288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6631
timestamp 1677677812
transform 1 0 1296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6633
timestamp 1677677812
transform 1 0 1304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6635
timestamp 1677677812
transform 1 0 1312 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_369
timestamp 1677677812
transform 1 0 1320 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6649
timestamp 1677677812
transform 1 0 1416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6651
timestamp 1677677812
transform 1 0 1424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6653
timestamp 1677677812
transform 1 0 1432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6655
timestamp 1677677812
transform 1 0 1440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6662
timestamp 1677677812
transform 1 0 1448 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_21
timestamp 1677677812
transform -1 0 1488 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6663
timestamp 1677677812
transform 1 0 1488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6665
timestamp 1677677812
transform 1 0 1496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6667
timestamp 1677677812
transform 1 0 1504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6669
timestamp 1677677812
transform 1 0 1512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6673
timestamp 1677677812
transform 1 0 1520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6674
timestamp 1677677812
transform 1 0 1528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6675
timestamp 1677677812
transform 1 0 1536 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5255
timestamp 1677677812
transform 1 0 1556 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_422
timestamp 1677677812
transform 1 0 1544 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6676
timestamp 1677677812
transform 1 0 1560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6682
timestamp 1677677812
transform 1 0 1568 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6683
timestamp 1677677812
transform 1 0 1576 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6684
timestamp 1677677812
transform 1 0 1584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6685
timestamp 1677677812
transform 1 0 1592 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_74
timestamp 1677677812
transform -1 0 1624 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_75
timestamp 1677677812
transform 1 0 1624 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6686
timestamp 1677677812
transform 1 0 1648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6688
timestamp 1677677812
transform 1 0 1656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6690
timestamp 1677677812
transform 1 0 1664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6693
timestamp 1677677812
transform 1 0 1672 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_77
timestamp 1677677812
transform -1 0 1704 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6694
timestamp 1677677812
transform 1 0 1704 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6696
timestamp 1677677812
transform 1 0 1712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6700
timestamp 1677677812
transform 1 0 1720 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_78
timestamp 1677677812
transform 1 0 1728 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6701
timestamp 1677677812
transform 1 0 1752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6703
timestamp 1677677812
transform 1 0 1760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6705
timestamp 1677677812
transform 1 0 1768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6708
timestamp 1677677812
transform 1 0 1776 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_80
timestamp 1677677812
transform 1 0 1784 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6709
timestamp 1677677812
transform 1 0 1808 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6713
timestamp 1677677812
transform 1 0 1816 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_82
timestamp 1677677812
transform -1 0 1848 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6714
timestamp 1677677812
transform 1 0 1848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6715
timestamp 1677677812
transform 1 0 1856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6717
timestamp 1677677812
transform 1 0 1864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6719
timestamp 1677677812
transform 1 0 1872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6721
timestamp 1677677812
transform 1 0 1880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6723
timestamp 1677677812
transform 1 0 1888 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_424
timestamp 1677677812
transform 1 0 1896 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6727
timestamp 1677677812
transform 1 0 1912 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6729
timestamp 1677677812
transform 1 0 1920 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6731
timestamp 1677677812
transform 1 0 1928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6733
timestamp 1677677812
transform 1 0 1936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6741
timestamp 1677677812
transform 1 0 1944 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_262
timestamp 1677677812
transform -1 0 1992 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6742
timestamp 1677677812
transform 1 0 1992 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6744
timestamp 1677677812
transform 1 0 2000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6754
timestamp 1677677812
transform 1 0 2008 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_370
timestamp 1677677812
transform -1 0 2112 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6755
timestamp 1677677812
transform 1 0 2112 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6757
timestamp 1677677812
transform 1 0 2120 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6759
timestamp 1677677812
transform 1 0 2128 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6761
timestamp 1677677812
transform 1 0 2136 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6763
timestamp 1677677812
transform 1 0 2144 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6767
timestamp 1677677812
transform 1 0 2152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6768
timestamp 1677677812
transform 1 0 2160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6769
timestamp 1677677812
transform 1 0 2168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6770
timestamp 1677677812
transform 1 0 2176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6771
timestamp 1677677812
transform 1 0 2184 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6772
timestamp 1677677812
transform 1 0 2192 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6773
timestamp 1677677812
transform 1 0 2200 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6774
timestamp 1677677812
transform 1 0 2208 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6775
timestamp 1677677812
transform 1 0 2216 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6776
timestamp 1677677812
transform 1 0 2224 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6777
timestamp 1677677812
transform 1 0 2232 0 -1 1970
box -8 -3 16 105
use BUFX2  BUFX2_83
timestamp 1677677812
transform -1 0 2264 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6778
timestamp 1677677812
transform 1 0 2264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6780
timestamp 1677677812
transform 1 0 2272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6782
timestamp 1677677812
transform 1 0 2280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6784
timestamp 1677677812
transform 1 0 2288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6786
timestamp 1677677812
transform 1 0 2296 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6788
timestamp 1677677812
transform 1 0 2304 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6797
timestamp 1677677812
transform 1 0 2312 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_425
timestamp 1677677812
transform -1 0 2336 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6798
timestamp 1677677812
transform 1 0 2336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6799
timestamp 1677677812
transform 1 0 2344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6800
timestamp 1677677812
transform 1 0 2352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6801
timestamp 1677677812
transform 1 0 2360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6802
timestamp 1677677812
transform 1 0 2368 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_22
timestamp 1677677812
transform 1 0 2376 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6803
timestamp 1677677812
transform 1 0 2408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6805
timestamp 1677677812
transform 1 0 2416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6807
timestamp 1677677812
transform 1 0 2424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6809
timestamp 1677677812
transform 1 0 2432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6811
timestamp 1677677812
transform 1 0 2440 0 -1 1970
box -8 -3 16 105
use AND2X2  AND2X2_23
timestamp 1677677812
transform 1 0 2448 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6815
timestamp 1677677812
transform 1 0 2480 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6817
timestamp 1677677812
transform 1 0 2488 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6819
timestamp 1677677812
transform 1 0 2496 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6821
timestamp 1677677812
transform 1 0 2504 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6823
timestamp 1677677812
transform 1 0 2512 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6825
timestamp 1677677812
transform 1 0 2520 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6827
timestamp 1677677812
transform 1 0 2528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6829
timestamp 1677677812
transform 1 0 2536 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_266
timestamp 1677677812
transform 1 0 2544 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6836
timestamp 1677677812
transform 1 0 2584 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6837
timestamp 1677677812
transform 1 0 2592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6838
timestamp 1677677812
transform 1 0 2600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6839
timestamp 1677677812
transform 1 0 2608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6840
timestamp 1677677812
transform 1 0 2616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6841
timestamp 1677677812
transform 1 0 2624 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6843
timestamp 1677677812
transform 1 0 2632 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6845
timestamp 1677677812
transform 1 0 2640 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6847
timestamp 1677677812
transform 1 0 2648 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6849
timestamp 1677677812
transform 1 0 2656 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6850
timestamp 1677677812
transform 1 0 2664 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6851
timestamp 1677677812
transform 1 0 2672 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6852
timestamp 1677677812
transform 1 0 2680 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6853
timestamp 1677677812
transform 1 0 2688 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6854
timestamp 1677677812
transform 1 0 2696 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5256
timestamp 1677677812
transform 1 0 2724 0 1 1875
box -3 -3 3 3
use AND2X2  AND2X2_24
timestamp 1677677812
transform -1 0 2736 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6855
timestamp 1677677812
transform 1 0 2736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6856
timestamp 1677677812
transform 1 0 2744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6857
timestamp 1677677812
transform 1 0 2752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6859
timestamp 1677677812
transform 1 0 2760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6861
timestamp 1677677812
transform 1 0 2768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6863
timestamp 1677677812
transform 1 0 2776 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_125
timestamp 1677677812
transform 1 0 2784 0 -1 1970
box -8 -3 34 105
use FILL  FILL_6868
timestamp 1677677812
transform 1 0 2816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6869
timestamp 1677677812
transform 1 0 2824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6870
timestamp 1677677812
transform 1 0 2832 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6871
timestamp 1677677812
transform 1 0 2840 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6873
timestamp 1677677812
transform 1 0 2848 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6875
timestamp 1677677812
transform 1 0 2856 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6877
timestamp 1677677812
transform 1 0 2864 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6879
timestamp 1677677812
transform 1 0 2872 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6881
timestamp 1677677812
transform 1 0 2880 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6885
timestamp 1677677812
transform 1 0 2888 0 -1 1970
box -8 -3 16 105
use OAI21X1  OAI21X1_127
timestamp 1677677812
transform -1 0 2928 0 -1 1970
box -8 -3 34 105
use FILL  FILL_6886
timestamp 1677677812
transform 1 0 2928 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6887
timestamp 1677677812
transform 1 0 2936 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6889
timestamp 1677677812
transform 1 0 2944 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6891
timestamp 1677677812
transform 1 0 2952 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6898
timestamp 1677677812
transform 1 0 2960 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6899
timestamp 1677677812
transform 1 0 2968 0 -1 1970
box -8 -3 16 105
use NOR2X1  NOR2X1_65
timestamp 1677677812
transform 1 0 2976 0 -1 1970
box -8 -3 32 105
use FILL  FILL_6900
timestamp 1677677812
transform 1 0 3000 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6901
timestamp 1677677812
transform 1 0 3008 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5257
timestamp 1677677812
transform 1 0 3036 0 1 1875
box -3 -3 3 3
use BUFX2  BUFX2_84
timestamp 1677677812
transform 1 0 3016 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6902
timestamp 1677677812
transform 1 0 3040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6903
timestamp 1677677812
transform 1 0 3048 0 -1 1970
box -8 -3 16 105
use M3_M2  M3_M2_5258
timestamp 1677677812
transform 1 0 3076 0 1 1875
box -3 -3 3 3
use INVX2  INVX2_427
timestamp 1677677812
transform -1 0 3072 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6904
timestamp 1677677812
transform 1 0 3072 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6905
timestamp 1677677812
transform 1 0 3080 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6906
timestamp 1677677812
transform 1 0 3088 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6907
timestamp 1677677812
transform 1 0 3096 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6908
timestamp 1677677812
transform 1 0 3104 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6909
timestamp 1677677812
transform 1 0 3112 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_43
timestamp 1677677812
transform -1 0 3152 0 -1 1970
box -8 -3 40 105
use FILL  FILL_6910
timestamp 1677677812
transform 1 0 3152 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6911
timestamp 1677677812
transform 1 0 3160 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6912
timestamp 1677677812
transform 1 0 3168 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6927
timestamp 1677677812
transform 1 0 3176 0 -1 1970
box -8 -3 16 105
use NAND3X1  NAND3X1_45
timestamp 1677677812
transform -1 0 3216 0 -1 1970
box -8 -3 40 105
use BUFX2  BUFX2_86
timestamp 1677677812
transform 1 0 3216 0 -1 1970
box -5 -3 28 105
use BUFX2  BUFX2_87
timestamp 1677677812
transform 1 0 3240 0 -1 1970
box -5 -3 28 105
use FILL  FILL_6928
timestamp 1677677812
transform 1 0 3264 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6929
timestamp 1677677812
transform 1 0 3272 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6930
timestamp 1677677812
transform 1 0 3280 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6931
timestamp 1677677812
transform 1 0 3288 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_267
timestamp 1677677812
transform 1 0 3296 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6932
timestamp 1677677812
transform 1 0 3336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6933
timestamp 1677677812
transform 1 0 3344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6934
timestamp 1677677812
transform 1 0 3352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6935
timestamp 1677677812
transform 1 0 3360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6936
timestamp 1677677812
transform 1 0 3368 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_428
timestamp 1677677812
transform 1 0 3376 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6940
timestamp 1677677812
transform 1 0 3392 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6943
timestamp 1677677812
transform 1 0 3400 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6944
timestamp 1677677812
transform 1 0 3408 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6945
timestamp 1677677812
transform 1 0 3416 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6946
timestamp 1677677812
transform 1 0 3424 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6947
timestamp 1677677812
transform 1 0 3432 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6948
timestamp 1677677812
transform 1 0 3440 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6949
timestamp 1677677812
transform 1 0 3448 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6951
timestamp 1677677812
transform 1 0 3456 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6953
timestamp 1677677812
transform 1 0 3464 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6955
timestamp 1677677812
transform 1 0 3472 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6959
timestamp 1677677812
transform 1 0 3480 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_268
timestamp 1677677812
transform 1 0 3488 0 -1 1970
box -8 -3 46 105
use FILL  FILL_6960
timestamp 1677677812
transform 1 0 3528 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6962
timestamp 1677677812
transform 1 0 3536 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6964
timestamp 1677677812
transform 1 0 3544 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6966
timestamp 1677677812
transform 1 0 3552 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6968
timestamp 1677677812
transform 1 0 3560 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6970
timestamp 1677677812
transform 1 0 3568 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_429
timestamp 1677677812
transform 1 0 3576 0 -1 1970
box -9 -3 26 105
use FILL  FILL_6974
timestamp 1677677812
transform 1 0 3592 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6976
timestamp 1677677812
transform 1 0 3600 0 -1 1970
box -8 -3 16 105
use FILL  FILL_6998
timestamp 1677677812
transform 1 0 3608 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_378
timestamp 1677677812
transform -1 0 3712 0 -1 1970
box -8 -3 104 105
use FILL  FILL_6999
timestamp 1677677812
transform 1 0 3712 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7000
timestamp 1677677812
transform 1 0 3720 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7001
timestamp 1677677812
transform 1 0 3728 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_432
timestamp 1677677812
transform -1 0 3752 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7002
timestamp 1677677812
transform 1 0 3752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7003
timestamp 1677677812
transform 1 0 3760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7004
timestamp 1677677812
transform 1 0 3768 0 -1 1970
box -8 -3 16 105
use AOI22X1  AOI22X1_270
timestamp 1677677812
transform 1 0 3776 0 -1 1970
box -8 -3 46 105
use FILL  FILL_7005
timestamp 1677677812
transform 1 0 3816 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7006
timestamp 1677677812
transform 1 0 3824 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7007
timestamp 1677677812
transform 1 0 3832 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_379
timestamp 1677677812
transform 1 0 3840 0 -1 1970
box -8 -3 104 105
use FILL  FILL_7008
timestamp 1677677812
transform 1 0 3936 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_380
timestamp 1677677812
transform -1 0 4040 0 -1 1970
box -8 -3 104 105
use FILL  FILL_7009
timestamp 1677677812
transform 1 0 4040 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7010
timestamp 1677677812
transform 1 0 4048 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7011
timestamp 1677677812
transform 1 0 4056 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_381
timestamp 1677677812
transform 1 0 4064 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_433
timestamp 1677677812
transform -1 0 4176 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7012
timestamp 1677677812
transform 1 0 4176 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7013
timestamp 1677677812
transform 1 0 4184 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_382
timestamp 1677677812
transform 1 0 4192 0 -1 1970
box -8 -3 104 105
use FILL  FILL_7014
timestamp 1677677812
transform 1 0 4288 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7015
timestamp 1677677812
transform 1 0 4296 0 -1 1970
box -8 -3 16 105
use INVX2  INVX2_434
timestamp 1677677812
transform -1 0 4320 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7016
timestamp 1677677812
transform 1 0 4320 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7017
timestamp 1677677812
transform 1 0 4328 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7018
timestamp 1677677812
transform 1 0 4336 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7019
timestamp 1677677812
transform 1 0 4344 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7020
timestamp 1677677812
transform 1 0 4352 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7021
timestamp 1677677812
transform 1 0 4360 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7022
timestamp 1677677812
transform 1 0 4368 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_383
timestamp 1677677812
transform 1 0 4376 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_435
timestamp 1677677812
transform -1 0 4488 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7034
timestamp 1677677812
transform 1 0 4488 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_384
timestamp 1677677812
transform 1 0 4496 0 -1 1970
box -8 -3 104 105
use INVX2  INVX2_438
timestamp 1677677812
transform -1 0 4608 0 -1 1970
box -9 -3 26 105
use FILL  FILL_7047
timestamp 1677677812
transform 1 0 4608 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7048
timestamp 1677677812
transform 1 0 4616 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7052
timestamp 1677677812
transform 1 0 4624 0 -1 1970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_386
timestamp 1677677812
transform -1 0 4728 0 -1 1970
box -8 -3 104 105
use FILL  FILL_7053
timestamp 1677677812
transform 1 0 4728 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7054
timestamp 1677677812
transform 1 0 4736 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7055
timestamp 1677677812
transform 1 0 4744 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7056
timestamp 1677677812
transform 1 0 4752 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7058
timestamp 1677677812
transform 1 0 4760 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7060
timestamp 1677677812
transform 1 0 4768 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7062
timestamp 1677677812
transform 1 0 4776 0 -1 1970
box -8 -3 16 105
use FILL  FILL_7064
timestamp 1677677812
transform 1 0 4784 0 -1 1970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_57
timestamp 1677677812
transform 1 0 4843 0 1 1870
box -10 -3 10 3
use M2_M1  M2_M1_6011
timestamp 1677677812
transform 1 0 84 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5371
timestamp 1677677812
transform 1 0 84 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5908
timestamp 1677677812
transform 1 0 100 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5400
timestamp 1677677812
transform 1 0 132 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5303
timestamp 1677677812
transform 1 0 204 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5304
timestamp 1677677812
transform 1 0 244 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5909
timestamp 1677677812
transform 1 0 204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5910
timestamp 1677677812
transform 1 0 236 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5911
timestamp 1677677812
transform 1 0 244 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5338
timestamp 1677677812
transform 1 0 252 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5912
timestamp 1677677812
transform 1 0 260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6012
timestamp 1677677812
transform 1 0 156 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5352
timestamp 1677677812
transform 1 0 236 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6013
timestamp 1677677812
transform 1 0 244 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5353
timestamp 1677677812
transform 1 0 260 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6014
timestamp 1677677812
transform 1 0 268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6015
timestamp 1677677812
transform 1 0 276 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5372
timestamp 1677677812
transform 1 0 156 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5373
timestamp 1677677812
transform 1 0 244 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5401
timestamp 1677677812
transform 1 0 260 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5339
timestamp 1677677812
transform 1 0 292 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5340
timestamp 1677677812
transform 1 0 308 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6016
timestamp 1677677812
transform 1 0 300 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5913
timestamp 1677677812
transform 1 0 332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5914
timestamp 1677677812
transform 1 0 348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6017
timestamp 1677677812
transform 1 0 340 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5374
timestamp 1677677812
transform 1 0 340 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5341
timestamp 1677677812
transform 1 0 380 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5915
timestamp 1677677812
transform 1 0 388 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5916
timestamp 1677677812
transform 1 0 404 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5917
timestamp 1677677812
transform 1 0 420 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6018
timestamp 1677677812
transform 1 0 372 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6019
timestamp 1677677812
transform 1 0 380 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5354
timestamp 1677677812
transform 1 0 388 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6020
timestamp 1677677812
transform 1 0 396 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5264
timestamp 1677677812
transform 1 0 436 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_6021
timestamp 1677677812
transform 1 0 436 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5265
timestamp 1677677812
transform 1 0 460 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5305
timestamp 1677677812
transform 1 0 452 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5306
timestamp 1677677812
transform 1 0 524 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5918
timestamp 1677677812
transform 1 0 492 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6022
timestamp 1677677812
transform 1 0 452 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5355
timestamp 1677677812
transform 1 0 540 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6023
timestamp 1677677812
transform 1 0 572 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5919
timestamp 1677677812
transform 1 0 596 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5375
timestamp 1677677812
transform 1 0 596 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5307
timestamp 1677677812
transform 1 0 652 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5920
timestamp 1677677812
transform 1 0 644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6024
timestamp 1677677812
transform 1 0 652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5921
timestamp 1677677812
transform 1 0 668 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5922
timestamp 1677677812
transform 1 0 684 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6025
timestamp 1677677812
transform 1 0 668 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5356
timestamp 1677677812
transform 1 0 676 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5376
timestamp 1677677812
transform 1 0 668 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5923
timestamp 1677677812
transform 1 0 724 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6026
timestamp 1677677812
transform 1 0 716 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5357
timestamp 1677677812
transform 1 0 724 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5266
timestamp 1677677812
transform 1 0 788 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5267
timestamp 1677677812
transform 1 0 820 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5276
timestamp 1677677812
transform 1 0 748 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5277
timestamp 1677677812
transform 1 0 780 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5924
timestamp 1677677812
transform 1 0 748 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5925
timestamp 1677677812
transform 1 0 804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6027
timestamp 1677677812
transform 1 0 828 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5377
timestamp 1677677812
transform 1 0 796 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5378
timestamp 1677677812
transform 1 0 812 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5926
timestamp 1677677812
transform 1 0 844 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5927
timestamp 1677677812
transform 1 0 860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5928
timestamp 1677677812
transform 1 0 956 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6028
timestamp 1677677812
transform 1 0 956 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5379
timestamp 1677677812
transform 1 0 956 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_6029
timestamp 1677677812
transform 1 0 964 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5929
timestamp 1677677812
transform 1 0 988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5930
timestamp 1677677812
transform 1 0 1012 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6030
timestamp 1677677812
transform 1 0 1012 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6031
timestamp 1677677812
transform 1 0 1028 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6106
timestamp 1677677812
transform 1 0 1020 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_6032
timestamp 1677677812
transform 1 0 1092 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5931
timestamp 1677677812
transform 1 0 1132 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5358
timestamp 1677677812
transform 1 0 1132 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5380
timestamp 1677677812
transform 1 0 1132 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5288
timestamp 1677677812
transform 1 0 1148 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5932
timestamp 1677677812
transform 1 0 1148 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5278
timestamp 1677677812
transform 1 0 1172 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5289
timestamp 1677677812
transform 1 0 1196 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5933
timestamp 1677677812
transform 1 0 1196 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6033
timestamp 1677677812
transform 1 0 1172 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5381
timestamp 1677677812
transform 1 0 1172 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5382
timestamp 1677677812
transform 1 0 1188 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5934
timestamp 1677677812
transform 1 0 1260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6034
timestamp 1677677812
transform 1 0 1260 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5279
timestamp 1677677812
transform 1 0 1292 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5280
timestamp 1677677812
transform 1 0 1340 0 1 1845
box -3 -3 3 3
use M2_M1  M2_M1_5935
timestamp 1677677812
transform 1 0 1316 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5936
timestamp 1677677812
transform 1 0 1340 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5937
timestamp 1677677812
transform 1 0 1348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6035
timestamp 1677677812
transform 1 0 1324 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5383
timestamp 1677677812
transform 1 0 1356 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5402
timestamp 1677677812
transform 1 0 1348 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6036
timestamp 1677677812
transform 1 0 1396 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5268
timestamp 1677677812
transform 1 0 1420 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5938
timestamp 1677677812
transform 1 0 1420 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5290
timestamp 1677677812
transform 1 0 1444 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5259
timestamp 1677677812
transform 1 0 1460 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5260
timestamp 1677677812
transform 1 0 1476 0 1 1865
box -3 -3 3 3
use M3_M2  M3_M2_5291
timestamp 1677677812
transform 1 0 1484 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5939
timestamp 1677677812
transform 1 0 1452 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5940
timestamp 1677677812
transform 1 0 1508 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6037
timestamp 1677677812
transform 1 0 1444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6038
timestamp 1677677812
transform 1 0 1532 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5308
timestamp 1677677812
transform 1 0 1660 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5941
timestamp 1677677812
transform 1 0 1604 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6039
timestamp 1677677812
transform 1 0 1580 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5359
timestamp 1677677812
transform 1 0 1652 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5269
timestamp 1677677812
transform 1 0 1716 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5281
timestamp 1677677812
transform 1 0 1732 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5309
timestamp 1677677812
transform 1 0 1716 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5310
timestamp 1677677812
transform 1 0 1740 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5942
timestamp 1677677812
transform 1 0 1716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5943
timestamp 1677677812
transform 1 0 1732 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5944
timestamp 1677677812
transform 1 0 1740 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6040
timestamp 1677677812
transform 1 0 1708 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6041
timestamp 1677677812
transform 1 0 1724 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5945
timestamp 1677677812
transform 1 0 1756 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5292
timestamp 1677677812
transform 1 0 1820 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5311
timestamp 1677677812
transform 1 0 1860 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5312
timestamp 1677677812
transform 1 0 1900 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5946
timestamp 1677677812
transform 1 0 1804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5947
timestamp 1677677812
transform 1 0 1860 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5948
timestamp 1677677812
transform 1 0 1900 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6042
timestamp 1677677812
transform 1 0 1780 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5360
timestamp 1677677812
transform 1 0 1788 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6043
timestamp 1677677812
transform 1 0 1796 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6044
timestamp 1677677812
transform 1 0 1884 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6045
timestamp 1677677812
transform 1 0 1900 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5384
timestamp 1677677812
transform 1 0 1780 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5385
timestamp 1677677812
transform 1 0 1804 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5386
timestamp 1677677812
transform 1 0 1836 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5313
timestamp 1677677812
transform 1 0 1948 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6046
timestamp 1677677812
transform 1 0 1948 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5314
timestamp 1677677812
transform 1 0 1972 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5949
timestamp 1677677812
transform 1 0 1964 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5950
timestamp 1677677812
transform 1 0 1980 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5315
timestamp 1677677812
transform 1 0 2052 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5951
timestamp 1677677812
transform 1 0 2052 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5342
timestamp 1677677812
transform 1 0 2060 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5952
timestamp 1677677812
transform 1 0 2068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6047
timestamp 1677677812
transform 1 0 2068 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5316
timestamp 1677677812
transform 1 0 2132 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5953
timestamp 1677677812
transform 1 0 2124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6048
timestamp 1677677812
transform 1 0 2132 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5387
timestamp 1677677812
transform 1 0 2124 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5270
timestamp 1677677812
transform 1 0 2156 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5954
timestamp 1677677812
transform 1 0 2148 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5955
timestamp 1677677812
transform 1 0 2188 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5956
timestamp 1677677812
transform 1 0 2204 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6049
timestamp 1677677812
transform 1 0 2196 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5403
timestamp 1677677812
transform 1 0 2196 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5317
timestamp 1677677812
transform 1 0 2236 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6050
timestamp 1677677812
transform 1 0 2244 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5282
timestamp 1677677812
transform 1 0 2260 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5361
timestamp 1677677812
transform 1 0 2260 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5957
timestamp 1677677812
transform 1 0 2276 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5362
timestamp 1677677812
transform 1 0 2276 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5261
timestamp 1677677812
transform 1 0 2292 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_6051
timestamp 1677677812
transform 1 0 2284 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6052
timestamp 1677677812
transform 1 0 2292 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5404
timestamp 1677677812
transform 1 0 2284 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5363
timestamp 1677677812
transform 1 0 2300 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6107
timestamp 1677677812
transform 1 0 2300 0 1 1795
box -2 -2 2 2
use M2_M1  M2_M1_5958
timestamp 1677677812
transform 1 0 2356 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6053
timestamp 1677677812
transform 1 0 2348 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5293
timestamp 1677677812
transform 1 0 2380 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5959
timestamp 1677677812
transform 1 0 2380 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6054
timestamp 1677677812
transform 1 0 2380 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5960
timestamp 1677677812
transform 1 0 2396 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5294
timestamp 1677677812
transform 1 0 2420 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5961
timestamp 1677677812
transform 1 0 2428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6055
timestamp 1677677812
transform 1 0 2420 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5962
timestamp 1677677812
transform 1 0 2468 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6056
timestamp 1677677812
transform 1 0 2460 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5388
timestamp 1677677812
transform 1 0 2468 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5262
timestamp 1677677812
transform 1 0 2524 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_5963
timestamp 1677677812
transform 1 0 2524 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5343
timestamp 1677677812
transform 1 0 2532 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6057
timestamp 1677677812
transform 1 0 2532 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5271
timestamp 1677677812
transform 1 0 2548 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5295
timestamp 1677677812
transform 1 0 2556 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5344
timestamp 1677677812
transform 1 0 2564 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5272
timestamp 1677677812
transform 1 0 2588 0 1 1855
box -3 -3 3 3
use M3_M2  M3_M2_5273
timestamp 1677677812
transform 1 0 2612 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5964
timestamp 1677677812
transform 1 0 2572 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5965
timestamp 1677677812
transform 1 0 2580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5966
timestamp 1677677812
transform 1 0 2612 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5364
timestamp 1677677812
transform 1 0 2572 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5365
timestamp 1677677812
transform 1 0 2612 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6058
timestamp 1677677812
transform 1 0 2660 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5318
timestamp 1677677812
transform 1 0 2732 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5902
timestamp 1677677812
transform 1 0 2740 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6059
timestamp 1677677812
transform 1 0 2724 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5366
timestamp 1677677812
transform 1 0 2756 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5967
timestamp 1677677812
transform 1 0 2804 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6060
timestamp 1677677812
transform 1 0 2820 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5319
timestamp 1677677812
transform 1 0 2860 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5968
timestamp 1677677812
transform 1 0 2860 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5263
timestamp 1677677812
transform 1 0 2876 0 1 1865
box -3 -3 3 3
use M2_M1  M2_M1_5969
timestamp 1677677812
transform 1 0 2884 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6061
timestamp 1677677812
transform 1 0 2876 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5367
timestamp 1677677812
transform 1 0 2884 0 1 1805
box -3 -3 3 3
use M3_M2  M3_M2_5320
timestamp 1677677812
transform 1 0 2900 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5903
timestamp 1677677812
transform 1 0 2908 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5904
timestamp 1677677812
transform 1 0 2932 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6062
timestamp 1677677812
transform 1 0 2924 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5321
timestamp 1677677812
transform 1 0 2972 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6063
timestamp 1677677812
transform 1 0 2972 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5296
timestamp 1677677812
transform 1 0 3004 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5905
timestamp 1677677812
transform 1 0 2996 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_6064
timestamp 1677677812
transform 1 0 3004 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6065
timestamp 1677677812
transform 1 0 3036 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5322
timestamp 1677677812
transform 1 0 3068 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5906
timestamp 1677677812
transform 1 0 3076 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5970
timestamp 1677677812
transform 1 0 3068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6066
timestamp 1677677812
transform 1 0 3108 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5901
timestamp 1677677812
transform 1 0 3132 0 1 1835
box -2 -2 2 2
use M2_M1  M2_M1_5907
timestamp 1677677812
transform 1 0 3148 0 1 1825
box -2 -2 2 2
use M2_M1  M2_M1_5971
timestamp 1677677812
transform 1 0 3140 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5345
timestamp 1677677812
transform 1 0 3156 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5972
timestamp 1677677812
transform 1 0 3180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6067
timestamp 1677677812
transform 1 0 3204 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5973
timestamp 1677677812
transform 1 0 3220 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5283
timestamp 1677677812
transform 1 0 3268 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5346
timestamp 1677677812
transform 1 0 3260 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6068
timestamp 1677677812
transform 1 0 3268 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6069
timestamp 1677677812
transform 1 0 3276 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5974
timestamp 1677677812
transform 1 0 3332 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6070
timestamp 1677677812
transform 1 0 3340 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5975
timestamp 1677677812
transform 1 0 3356 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5274
timestamp 1677677812
transform 1 0 3436 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5976
timestamp 1677677812
transform 1 0 3372 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5977
timestamp 1677677812
transform 1 0 3428 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6071
timestamp 1677677812
transform 1 0 3452 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5389
timestamp 1677677812
transform 1 0 3388 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5390
timestamp 1677677812
transform 1 0 3452 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5275
timestamp 1677677812
transform 1 0 3524 0 1 1855
box -3 -3 3 3
use M2_M1  M2_M1_5978
timestamp 1677677812
transform 1 0 3532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5979
timestamp 1677677812
transform 1 0 3580 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5980
timestamp 1677677812
transform 1 0 3588 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6072
timestamp 1677677812
transform 1 0 3500 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5391
timestamp 1677677812
transform 1 0 3500 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5368
timestamp 1677677812
transform 1 0 3588 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6073
timestamp 1677677812
transform 1 0 3612 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6074
timestamp 1677677812
transform 1 0 3628 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5297
timestamp 1677677812
transform 1 0 3716 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_5981
timestamp 1677677812
transform 1 0 3716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5982
timestamp 1677677812
transform 1 0 3732 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5284
timestamp 1677677812
transform 1 0 3748 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5323
timestamp 1677677812
transform 1 0 3748 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5298
timestamp 1677677812
transform 1 0 3812 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5324
timestamp 1677677812
transform 1 0 3796 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5325
timestamp 1677677812
transform 1 0 3828 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5326
timestamp 1677677812
transform 1 0 3892 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5983
timestamp 1677677812
transform 1 0 3780 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5984
timestamp 1677677812
transform 1 0 3796 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5985
timestamp 1677677812
transform 1 0 3828 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5347
timestamp 1677677812
transform 1 0 3876 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5986
timestamp 1677677812
transform 1 0 3892 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6075
timestamp 1677677812
transform 1 0 3748 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6076
timestamp 1677677812
transform 1 0 3756 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6077
timestamp 1677677812
transform 1 0 3772 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6078
timestamp 1677677812
transform 1 0 3788 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6079
timestamp 1677677812
transform 1 0 3876 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5392
timestamp 1677677812
transform 1 0 3772 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5393
timestamp 1677677812
transform 1 0 3828 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5405
timestamp 1677677812
transform 1 0 3788 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5348
timestamp 1677677812
transform 1 0 3908 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5369
timestamp 1677677812
transform 1 0 3900 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_5987
timestamp 1677677812
transform 1 0 3932 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6080
timestamp 1677677812
transform 1 0 3924 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6081
timestamp 1677677812
transform 1 0 3940 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6082
timestamp 1677677812
transform 1 0 3948 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5394
timestamp 1677677812
transform 1 0 3948 0 1 1795
box -3 -3 3 3
use M2_M1  M2_M1_5988
timestamp 1677677812
transform 1 0 3988 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6083
timestamp 1677677812
transform 1 0 3980 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6084
timestamp 1677677812
transform 1 0 3996 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5406
timestamp 1677677812
transform 1 0 3996 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5349
timestamp 1677677812
transform 1 0 4028 0 1 1815
box -3 -3 3 3
use M3_M2  M3_M2_5327
timestamp 1677677812
transform 1 0 4076 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5989
timestamp 1677677812
transform 1 0 4068 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5990
timestamp 1677677812
transform 1 0 4124 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5991
timestamp 1677677812
transform 1 0 4132 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6085
timestamp 1677677812
transform 1 0 4044 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6086
timestamp 1677677812
transform 1 0 4140 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5395
timestamp 1677677812
transform 1 0 4140 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5328
timestamp 1677677812
transform 1 0 4180 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5992
timestamp 1677677812
transform 1 0 4164 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5993
timestamp 1677677812
transform 1 0 4180 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6087
timestamp 1677677812
transform 1 0 4172 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5370
timestamp 1677677812
transform 1 0 4180 0 1 1805
box -3 -3 3 3
use M2_M1  M2_M1_6088
timestamp 1677677812
transform 1 0 4188 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6089
timestamp 1677677812
transform 1 0 4196 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5396
timestamp 1677677812
transform 1 0 4196 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5407
timestamp 1677677812
transform 1 0 4188 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5299
timestamp 1677677812
transform 1 0 4212 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5300
timestamp 1677677812
transform 1 0 4244 0 1 1835
box -3 -3 3 3
use M3_M2  M3_M2_5329
timestamp 1677677812
transform 1 0 4228 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5994
timestamp 1677677812
transform 1 0 4228 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_5995
timestamp 1677677812
transform 1 0 4244 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6090
timestamp 1677677812
transform 1 0 4236 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5330
timestamp 1677677812
transform 1 0 4260 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5996
timestamp 1677677812
transform 1 0 4260 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6091
timestamp 1677677812
transform 1 0 4268 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5408
timestamp 1677677812
transform 1 0 4268 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6092
timestamp 1677677812
transform 1 0 4284 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5350
timestamp 1677677812
transform 1 0 4324 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_5997
timestamp 1677677812
transform 1 0 4348 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6093
timestamp 1677677812
transform 1 0 4324 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_5998
timestamp 1677677812
transform 1 0 4412 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5331
timestamp 1677677812
transform 1 0 4460 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_5999
timestamp 1677677812
transform 1 0 4436 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6000
timestamp 1677677812
transform 1 0 4452 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6001
timestamp 1677677812
transform 1 0 4476 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6094
timestamp 1677677812
transform 1 0 4428 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6095
timestamp 1677677812
transform 1 0 4444 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6096
timestamp 1677677812
transform 1 0 4460 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6097
timestamp 1677677812
transform 1 0 4468 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5409
timestamp 1677677812
transform 1 0 4428 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5397
timestamp 1677677812
transform 1 0 4460 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5410
timestamp 1677677812
transform 1 0 4468 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5285
timestamp 1677677812
transform 1 0 4524 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5286
timestamp 1677677812
transform 1 0 4540 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5287
timestamp 1677677812
transform 1 0 4596 0 1 1845
box -3 -3 3 3
use M3_M2  M3_M2_5332
timestamp 1677677812
transform 1 0 4516 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5301
timestamp 1677677812
transform 1 0 4620 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6002
timestamp 1677677812
transform 1 0 4500 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6003
timestamp 1677677812
transform 1 0 4524 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6004
timestamp 1677677812
transform 1 0 4532 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6005
timestamp 1677677812
transform 1 0 4564 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5351
timestamp 1677677812
transform 1 0 4612 0 1 1815
box -3 -3 3 3
use M2_M1  M2_M1_6098
timestamp 1677677812
transform 1 0 4508 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6099
timestamp 1677677812
transform 1 0 4524 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6100
timestamp 1677677812
transform 1 0 4612 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5398
timestamp 1677677812
transform 1 0 4564 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5333
timestamp 1677677812
transform 1 0 4628 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6101
timestamp 1677677812
transform 1 0 4628 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5302
timestamp 1677677812
transform 1 0 4644 0 1 1835
box -3 -3 3 3
use M2_M1  M2_M1_6006
timestamp 1677677812
transform 1 0 4644 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6007
timestamp 1677677812
transform 1 0 4660 0 1 1815
box -2 -2 2 2
use M3_M2  M3_M2_5334
timestamp 1677677812
transform 1 0 4684 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5335
timestamp 1677677812
transform 1 0 4716 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5336
timestamp 1677677812
transform 1 0 4764 0 1 1825
box -3 -3 3 3
use M3_M2  M3_M2_5337
timestamp 1677677812
transform 1 0 4788 0 1 1825
box -3 -3 3 3
use M2_M1  M2_M1_6008
timestamp 1677677812
transform 1 0 4716 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6009
timestamp 1677677812
transform 1 0 4764 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6010
timestamp 1677677812
transform 1 0 4772 0 1 1815
box -2 -2 2 2
use M2_M1  M2_M1_6102
timestamp 1677677812
transform 1 0 4652 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6103
timestamp 1677677812
transform 1 0 4668 0 1 1805
box -2 -2 2 2
use M2_M1  M2_M1_6104
timestamp 1677677812
transform 1 0 4684 0 1 1805
box -2 -2 2 2
use M3_M2  M3_M2_5399
timestamp 1677677812
transform 1 0 4684 0 1 1795
box -3 -3 3 3
use M3_M2  M3_M2_5411
timestamp 1677677812
transform 1 0 4668 0 1 1785
box -3 -3 3 3
use M3_M2  M3_M2_5412
timestamp 1677677812
transform 1 0 4684 0 1 1785
box -3 -3 3 3
use M2_M1  M2_M1_6105
timestamp 1677677812
transform 1 0 4788 0 1 1805
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_58
timestamp 1677677812
transform 1 0 48 0 1 1770
box -10 -3 10 3
use FILL  FILL_7065
timestamp 1677677812
transform 1 0 72 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_88
timestamp 1677677812
transform -1 0 104 0 1 1770
box -5 -3 28 105
use FILL  FILL_7066
timestamp 1677677812
transform 1 0 104 0 1 1770
box -8 -3 16 105
use FILL  FILL_7067
timestamp 1677677812
transform 1 0 112 0 1 1770
box -8 -3 16 105
use FILL  FILL_7068
timestamp 1677677812
transform 1 0 120 0 1 1770
box -8 -3 16 105
use FILL  FILL_7069
timestamp 1677677812
transform 1 0 128 0 1 1770
box -8 -3 16 105
use FILL  FILL_7070
timestamp 1677677812
transform 1 0 136 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_387
timestamp 1677677812
transform 1 0 144 0 1 1770
box -8 -3 104 105
use M3_M2  M3_M2_5413
timestamp 1677677812
transform 1 0 260 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_271
timestamp 1677677812
transform 1 0 240 0 1 1770
box -8 -3 46 105
use FILL  FILL_7071
timestamp 1677677812
transform 1 0 280 0 1 1770
box -8 -3 16 105
use FILL  FILL_7072
timestamp 1677677812
transform 1 0 288 0 1 1770
box -8 -3 16 105
use FILL  FILL_7073
timestamp 1677677812
transform 1 0 296 0 1 1770
box -8 -3 16 105
use FILL  FILL_7074
timestamp 1677677812
transform 1 0 304 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5414
timestamp 1677677812
transform 1 0 332 0 1 1775
box -3 -3 3 3
use AOI22X1  AOI22X1_272
timestamp 1677677812
transform -1 0 352 0 1 1770
box -8 -3 46 105
use FILL  FILL_7075
timestamp 1677677812
transform 1 0 352 0 1 1770
box -8 -3 16 105
use FILL  FILL_7076
timestamp 1677677812
transform 1 0 360 0 1 1770
box -8 -3 16 105
use FILL  FILL_7077
timestamp 1677677812
transform 1 0 368 0 1 1770
box -8 -3 16 105
use FILL  FILL_7078
timestamp 1677677812
transform 1 0 376 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_274
timestamp 1677677812
transform 1 0 384 0 1 1770
box -8 -3 46 105
use FILL  FILL_7085
timestamp 1677677812
transform 1 0 424 0 1 1770
box -8 -3 16 105
use FILL  FILL_7087
timestamp 1677677812
transform 1 0 432 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5415
timestamp 1677677812
transform 1 0 468 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_390
timestamp 1677677812
transform 1 0 440 0 1 1770
box -8 -3 104 105
use FILL  FILL_7089
timestamp 1677677812
transform 1 0 536 0 1 1770
box -8 -3 16 105
use FILL  FILL_7090
timestamp 1677677812
transform 1 0 544 0 1 1770
box -8 -3 16 105
use FILL  FILL_7098
timestamp 1677677812
transform 1 0 552 0 1 1770
box -8 -3 16 105
use FILL  FILL_7100
timestamp 1677677812
transform 1 0 560 0 1 1770
box -8 -3 16 105
use FILL  FILL_7101
timestamp 1677677812
transform 1 0 568 0 1 1770
box -8 -3 16 105
use FILL  FILL_7102
timestamp 1677677812
transform 1 0 576 0 1 1770
box -8 -3 16 105
use FILL  FILL_7103
timestamp 1677677812
transform 1 0 584 0 1 1770
box -8 -3 16 105
use FILL  FILL_7104
timestamp 1677677812
transform 1 0 592 0 1 1770
box -8 -3 16 105
use FILL  FILL_7105
timestamp 1677677812
transform 1 0 600 0 1 1770
box -8 -3 16 105
use FILL  FILL_7107
timestamp 1677677812
transform 1 0 608 0 1 1770
box -8 -3 16 105
use FILL  FILL_7109
timestamp 1677677812
transform 1 0 616 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_30
timestamp 1677677812
transform -1 0 656 0 1 1770
box -8 -3 40 105
use FILL  FILL_7110
timestamp 1677677812
transform 1 0 656 0 1 1770
box -8 -3 16 105
use FILL  FILL_7111
timestamp 1677677812
transform 1 0 664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7112
timestamp 1677677812
transform 1 0 672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7116
timestamp 1677677812
transform 1 0 680 0 1 1770
box -8 -3 16 105
use FILL  FILL_7118
timestamp 1677677812
transform 1 0 688 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_259
timestamp 1677677812
transform 1 0 696 0 1 1770
box -8 -3 46 105
use FILL  FILL_7120
timestamp 1677677812
transform 1 0 736 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_391
timestamp 1677677812
transform -1 0 840 0 1 1770
box -8 -3 104 105
use FILL  FILL_7121
timestamp 1677677812
transform 1 0 840 0 1 1770
box -8 -3 16 105
use FILL  FILL_7122
timestamp 1677677812
transform 1 0 848 0 1 1770
box -8 -3 16 105
use FILL  FILL_7123
timestamp 1677677812
transform 1 0 856 0 1 1770
box -8 -3 16 105
use FILL  FILL_7124
timestamp 1677677812
transform 1 0 864 0 1 1770
box -8 -3 16 105
use FILL  FILL_7125
timestamp 1677677812
transform 1 0 872 0 1 1770
box -8 -3 16 105
use FILL  FILL_7126
timestamp 1677677812
transform 1 0 880 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_89
timestamp 1677677812
transform 1 0 888 0 1 1770
box -5 -3 28 105
use FILL  FILL_7127
timestamp 1677677812
transform 1 0 912 0 1 1770
box -8 -3 16 105
use FILL  FILL_7137
timestamp 1677677812
transform 1 0 920 0 1 1770
box -8 -3 16 105
use FILL  FILL_7139
timestamp 1677677812
transform 1 0 928 0 1 1770
box -8 -3 16 105
use FILL  FILL_7141
timestamp 1677677812
transform 1 0 936 0 1 1770
box -8 -3 16 105
use FILL  FILL_7142
timestamp 1677677812
transform 1 0 944 0 1 1770
box -8 -3 16 105
use FILL  FILL_7143
timestamp 1677677812
transform 1 0 952 0 1 1770
box -8 -3 16 105
use FILL  FILL_7144
timestamp 1677677812
transform 1 0 960 0 1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_278
timestamp 1677677812
transform -1 0 1008 0 1 1770
box -8 -3 46 105
use M3_M2  M3_M2_5416
timestamp 1677677812
transform 1 0 1020 0 1 1775
box -3 -3 3 3
use FILL  FILL_7145
timestamp 1677677812
transform 1 0 1008 0 1 1770
box -8 -3 16 105
use FILL  FILL_7153
timestamp 1677677812
transform 1 0 1016 0 1 1770
box -8 -3 16 105
use FILL  FILL_7155
timestamp 1677677812
transform 1 0 1024 0 1 1770
box -8 -3 16 105
use FILL  FILL_7157
timestamp 1677677812
transform 1 0 1032 0 1 1770
box -8 -3 16 105
use FILL  FILL_7159
timestamp 1677677812
transform 1 0 1040 0 1 1770
box -8 -3 16 105
use FILL  FILL_7161
timestamp 1677677812
transform 1 0 1048 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_67
timestamp 1677677812
transform 1 0 1056 0 1 1770
box -8 -3 32 105
use FILL  FILL_7163
timestamp 1677677812
transform 1 0 1080 0 1 1770
box -8 -3 16 105
use FILL  FILL_7164
timestamp 1677677812
transform 1 0 1088 0 1 1770
box -8 -3 16 105
use FILL  FILL_7165
timestamp 1677677812
transform 1 0 1096 0 1 1770
box -8 -3 16 105
use FILL  FILL_7166
timestamp 1677677812
transform 1 0 1104 0 1 1770
box -8 -3 16 105
use FILL  FILL_7167
timestamp 1677677812
transform 1 0 1112 0 1 1770
box -8 -3 16 105
use FILL  FILL_7171
timestamp 1677677812
transform 1 0 1120 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_444
timestamp 1677677812
transform 1 0 1128 0 1 1770
box -9 -3 26 105
use FILL  FILL_7173
timestamp 1677677812
transform 1 0 1144 0 1 1770
box -8 -3 16 105
use FILL  FILL_7177
timestamp 1677677812
transform 1 0 1152 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_393
timestamp 1677677812
transform 1 0 1160 0 1 1770
box -8 -3 104 105
use FILL  FILL_7179
timestamp 1677677812
transform 1 0 1256 0 1 1770
box -8 -3 16 105
use FILL  FILL_7189
timestamp 1677677812
transform 1 0 1264 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5417
timestamp 1677677812
transform 1 0 1284 0 1 1775
box -3 -3 3 3
use FILL  FILL_7191
timestamp 1677677812
transform 1 0 1272 0 1 1770
box -8 -3 16 105
use FILL  FILL_7193
timestamp 1677677812
transform 1 0 1280 0 1 1770
box -8 -3 16 105
use FILL  FILL_7194
timestamp 1677677812
transform 1 0 1288 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5418
timestamp 1677677812
transform 1 0 1308 0 1 1775
box -3 -3 3 3
use FILL  FILL_7195
timestamp 1677677812
transform 1 0 1296 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_260
timestamp 1677677812
transform -1 0 1344 0 1 1770
box -8 -3 46 105
use FILL  FILL_7196
timestamp 1677677812
transform 1 0 1344 0 1 1770
box -8 -3 16 105
use FILL  FILL_7202
timestamp 1677677812
transform 1 0 1352 0 1 1770
box -8 -3 16 105
use FILL  FILL_7204
timestamp 1677677812
transform 1 0 1360 0 1 1770
box -8 -3 16 105
use FILL  FILL_7205
timestamp 1677677812
transform 1 0 1368 0 1 1770
box -8 -3 16 105
use FILL  FILL_7206
timestamp 1677677812
transform 1 0 1376 0 1 1770
box -8 -3 16 105
use FILL  FILL_7207
timestamp 1677677812
transform 1 0 1384 0 1 1770
box -8 -3 16 105
use FILL  FILL_7208
timestamp 1677677812
transform 1 0 1392 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_33
timestamp 1677677812
transform -1 0 1432 0 1 1770
box -8 -3 40 105
use FILL  FILL_7209
timestamp 1677677812
transform 1 0 1432 0 1 1770
box -8 -3 16 105
use FILL  FILL_7216
timestamp 1677677812
transform 1 0 1440 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_394
timestamp 1677677812
transform -1 0 1544 0 1 1770
box -8 -3 104 105
use FILL  FILL_7217
timestamp 1677677812
transform 1 0 1544 0 1 1770
box -8 -3 16 105
use FILL  FILL_7218
timestamp 1677677812
transform 1 0 1552 0 1 1770
box -8 -3 16 105
use FILL  FILL_7219
timestamp 1677677812
transform 1 0 1560 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_395
timestamp 1677677812
transform 1 0 1568 0 1 1770
box -8 -3 104 105
use FILL  FILL_7227
timestamp 1677677812
transform 1 0 1664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7239
timestamp 1677677812
transform 1 0 1672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7241
timestamp 1677677812
transform 1 0 1680 0 1 1770
box -8 -3 16 105
use FILL  FILL_7243
timestamp 1677677812
transform 1 0 1688 0 1 1770
box -8 -3 16 105
use FILL  FILL_7245
timestamp 1677677812
transform 1 0 1696 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_261
timestamp 1677677812
transform -1 0 1744 0 1 1770
box -8 -3 46 105
use FILL  FILL_7246
timestamp 1677677812
transform 1 0 1744 0 1 1770
box -8 -3 16 105
use FILL  FILL_7247
timestamp 1677677812
transform 1 0 1752 0 1 1770
box -8 -3 16 105
use FILL  FILL_7251
timestamp 1677677812
transform 1 0 1760 0 1 1770
box -8 -3 16 105
use FILL  FILL_7253
timestamp 1677677812
transform 1 0 1768 0 1 1770
box -8 -3 16 105
use FILL  FILL_7255
timestamp 1677677812
transform 1 0 1776 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_446
timestamp 1677677812
transform -1 0 1800 0 1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_396
timestamp 1677677812
transform -1 0 1896 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_447
timestamp 1677677812
transform 1 0 1896 0 1 1770
box -9 -3 26 105
use FILL  FILL_7256
timestamp 1677677812
transform 1 0 1912 0 1 1770
box -8 -3 16 105
use FILL  FILL_7257
timestamp 1677677812
transform 1 0 1920 0 1 1770
box -8 -3 16 105
use FILL  FILL_7258
timestamp 1677677812
transform 1 0 1928 0 1 1770
box -8 -3 16 105
use FILL  FILL_7259
timestamp 1677677812
transform 1 0 1936 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_448
timestamp 1677677812
transform 1 0 1944 0 1 1770
box -9 -3 26 105
use FILL  FILL_7260
timestamp 1677677812
transform 1 0 1960 0 1 1770
box -8 -3 16 105
use FILL  FILL_7261
timestamp 1677677812
transform 1 0 1968 0 1 1770
box -8 -3 16 105
use FILL  FILL_7262
timestamp 1677677812
transform 1 0 1976 0 1 1770
box -8 -3 16 105
use FILL  FILL_7263
timestamp 1677677812
transform 1 0 1984 0 1 1770
box -8 -3 16 105
use FILL  FILL_7264
timestamp 1677677812
transform 1 0 1992 0 1 1770
box -8 -3 16 105
use FILL  FILL_7265
timestamp 1677677812
transform 1 0 2000 0 1 1770
box -8 -3 16 105
use FILL  FILL_7266
timestamp 1677677812
transform 1 0 2008 0 1 1770
box -8 -3 16 105
use FILL  FILL_7276
timestamp 1677677812
transform 1 0 2016 0 1 1770
box -8 -3 16 105
use FILL  FILL_7278
timestamp 1677677812
transform 1 0 2024 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_37
timestamp 1677677812
transform -1 0 2064 0 1 1770
box -8 -3 40 105
use FILL  FILL_7279
timestamp 1677677812
transform 1 0 2064 0 1 1770
box -8 -3 16 105
use FILL  FILL_7280
timestamp 1677677812
transform 1 0 2072 0 1 1770
box -8 -3 16 105
use FILL  FILL_7284
timestamp 1677677812
transform 1 0 2080 0 1 1770
box -8 -3 16 105
use FILL  FILL_7286
timestamp 1677677812
transform 1 0 2088 0 1 1770
box -8 -3 16 105
use FILL  FILL_7288
timestamp 1677677812
transform 1 0 2096 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5419
timestamp 1677677812
transform 1 0 2132 0 1 1775
box -3 -3 3 3
use AND2X2  AND2X2_39
timestamp 1677677812
transform -1 0 2136 0 1 1770
box -8 -3 40 105
use FILL  FILL_7289
timestamp 1677677812
transform 1 0 2136 0 1 1770
box -8 -3 16 105
use FILL  FILL_7290
timestamp 1677677812
transform 1 0 2144 0 1 1770
box -8 -3 16 105
use FILL  FILL_7294
timestamp 1677677812
transform 1 0 2152 0 1 1770
box -8 -3 16 105
use FILL  FILL_7296
timestamp 1677677812
transform 1 0 2160 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_41
timestamp 1677677812
transform -1 0 2200 0 1 1770
box -8 -3 40 105
use FILL  FILL_7298
timestamp 1677677812
transform 1 0 2200 0 1 1770
box -8 -3 16 105
use FILL  FILL_7300
timestamp 1677677812
transform 1 0 2208 0 1 1770
box -8 -3 16 105
use FILL  FILL_7302
timestamp 1677677812
transform 1 0 2216 0 1 1770
box -8 -3 16 105
use FILL  FILL_7304
timestamp 1677677812
transform 1 0 2224 0 1 1770
box -8 -3 16 105
use FILL  FILL_7306
timestamp 1677677812
transform 1 0 2232 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5420
timestamp 1677677812
transform 1 0 2260 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_449
timestamp 1677677812
transform 1 0 2240 0 1 1770
box -9 -3 26 105
use FILL  FILL_7308
timestamp 1677677812
transform 1 0 2256 0 1 1770
box -8 -3 16 105
use FILL  FILL_7309
timestamp 1677677812
transform 1 0 2264 0 1 1770
box -8 -3 16 105
use FILL  FILL_7310
timestamp 1677677812
transform 1 0 2272 0 1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_68
timestamp 1677677812
transform -1 0 2304 0 1 1770
box -8 -3 32 105
use FILL  FILL_7311
timestamp 1677677812
transform 1 0 2304 0 1 1770
box -8 -3 16 105
use FILL  FILL_7312
timestamp 1677677812
transform 1 0 2312 0 1 1770
box -8 -3 16 105
use FILL  FILL_7313
timestamp 1677677812
transform 1 0 2320 0 1 1770
box -8 -3 16 105
use FILL  FILL_7314
timestamp 1677677812
transform 1 0 2328 0 1 1770
box -8 -3 16 105
use FILL  FILL_7319
timestamp 1677677812
transform 1 0 2336 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_43
timestamp 1677677812
transform 1 0 2344 0 1 1770
box -8 -3 40 105
use FILL  FILL_7321
timestamp 1677677812
transform 1 0 2376 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_44
timestamp 1677677812
transform 1 0 2384 0 1 1770
box -8 -3 40 105
use FILL  FILL_7322
timestamp 1677677812
transform 1 0 2416 0 1 1770
box -8 -3 16 105
use FILL  FILL_7323
timestamp 1677677812
transform 1 0 2424 0 1 1770
box -8 -3 16 105
use FILL  FILL_7324
timestamp 1677677812
transform 1 0 2432 0 1 1770
box -8 -3 16 105
use FILL  FILL_7325
timestamp 1677677812
transform 1 0 2440 0 1 1770
box -8 -3 16 105
use FILL  FILL_7331
timestamp 1677677812
transform 1 0 2448 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_47
timestamp 1677677812
transform 1 0 2456 0 1 1770
box -8 -3 40 105
use FILL  FILL_7332
timestamp 1677677812
transform 1 0 2488 0 1 1770
box -8 -3 16 105
use FILL  FILL_7334
timestamp 1677677812
transform 1 0 2496 0 1 1770
box -8 -3 16 105
use FILL  FILL_7336
timestamp 1677677812
transform 1 0 2504 0 1 1770
box -8 -3 16 105
use FILL  FILL_7338
timestamp 1677677812
transform 1 0 2512 0 1 1770
box -8 -3 16 105
use FILL  FILL_7339
timestamp 1677677812
transform 1 0 2520 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_452
timestamp 1677677812
transform 1 0 2528 0 1 1770
box -9 -3 26 105
use FILL  FILL_7340
timestamp 1677677812
transform 1 0 2544 0 1 1770
box -8 -3 16 105
use FILL  FILL_7341
timestamp 1677677812
transform 1 0 2552 0 1 1770
box -8 -3 16 105
use FILL  FILL_7344
timestamp 1677677812
transform 1 0 2560 0 1 1770
box -8 -3 16 105
use FILL  FILL_7345
timestamp 1677677812
transform 1 0 2568 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5421
timestamp 1677677812
transform 1 0 2628 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5422
timestamp 1677677812
transform 1 0 2668 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_398
timestamp 1677677812
transform -1 0 2672 0 1 1770
box -8 -3 104 105
use FILL  FILL_7346
timestamp 1677677812
transform 1 0 2672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7350
timestamp 1677677812
transform 1 0 2680 0 1 1770
box -8 -3 16 105
use FILL  FILL_7352
timestamp 1677677812
transform 1 0 2688 0 1 1770
box -8 -3 16 105
use FILL  FILL_7354
timestamp 1677677812
transform 1 0 2696 0 1 1770
box -8 -3 16 105
use FILL  FILL_7356
timestamp 1677677812
transform 1 0 2704 0 1 1770
box -8 -3 16 105
use FILL  FILL_7358
timestamp 1677677812
transform 1 0 2712 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_455
timestamp 1677677812
transform 1 0 2720 0 1 1770
box -9 -3 26 105
use FILL  FILL_7359
timestamp 1677677812
transform 1 0 2736 0 1 1770
box -8 -3 16 105
use FILL  FILL_7360
timestamp 1677677812
transform 1 0 2744 0 1 1770
box -8 -3 16 105
use FILL  FILL_7362
timestamp 1677677812
transform 1 0 2752 0 1 1770
box -8 -3 16 105
use FILL  FILL_7364
timestamp 1677677812
transform 1 0 2760 0 1 1770
box -8 -3 16 105
use FILL  FILL_7366
timestamp 1677677812
transform 1 0 2768 0 1 1770
box -8 -3 16 105
use FILL  FILL_7368
timestamp 1677677812
transform 1 0 2776 0 1 1770
box -8 -3 16 105
use FILL  FILL_7370
timestamp 1677677812
transform 1 0 2784 0 1 1770
box -8 -3 16 105
use FILL  FILL_7371
timestamp 1677677812
transform 1 0 2792 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5423
timestamp 1677677812
transform 1 0 2812 0 1 1775
box -3 -3 3 3
use NAND2X1  NAND2X1_3
timestamp 1677677812
transform -1 0 2824 0 1 1770
box -8 -3 32 105
use FILL  FILL_7372
timestamp 1677677812
transform 1 0 2824 0 1 1770
box -8 -3 16 105
use FILL  FILL_7377
timestamp 1677677812
transform 1 0 2832 0 1 1770
box -8 -3 16 105
use FILL  FILL_7379
timestamp 1677677812
transform 1 0 2840 0 1 1770
box -8 -3 16 105
use FILL  FILL_7381
timestamp 1677677812
transform 1 0 2848 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_457
timestamp 1677677812
transform 1 0 2856 0 1 1770
box -9 -3 26 105
use FILL  FILL_7383
timestamp 1677677812
transform 1 0 2872 0 1 1770
box -8 -3 16 105
use FILL  FILL_7384
timestamp 1677677812
transform 1 0 2880 0 1 1770
box -8 -3 16 105
use FILL  FILL_7385
timestamp 1677677812
transform 1 0 2888 0 1 1770
box -8 -3 16 105
use FILL  FILL_7386
timestamp 1677677812
transform 1 0 2896 0 1 1770
box -8 -3 16 105
use NAND2X1  NAND2X1_4
timestamp 1677677812
transform 1 0 2904 0 1 1770
box -8 -3 32 105
use FILL  FILL_7387
timestamp 1677677812
transform 1 0 2928 0 1 1770
box -8 -3 16 105
use FILL  FILL_7391
timestamp 1677677812
transform 1 0 2936 0 1 1770
box -8 -3 16 105
use FILL  FILL_7393
timestamp 1677677812
transform 1 0 2944 0 1 1770
box -8 -3 16 105
use FILL  FILL_7394
timestamp 1677677812
transform 1 0 2952 0 1 1770
box -8 -3 16 105
use FILL  FILL_7395
timestamp 1677677812
transform 1 0 2960 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5424
timestamp 1677677812
transform 1 0 2996 0 1 1775
box -3 -3 3 3
use OAI21X1  OAI21X1_128
timestamp 1677677812
transform 1 0 2968 0 1 1770
box -8 -3 34 105
use FILL  FILL_7396
timestamp 1677677812
transform 1 0 3000 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5425
timestamp 1677677812
transform 1 0 3036 0 1 1775
box -3 -3 3 3
use OAI21X1  OAI21X1_129
timestamp 1677677812
transform -1 0 3040 0 1 1770
box -8 -3 34 105
use FILL  FILL_7397
timestamp 1677677812
transform 1 0 3040 0 1 1770
box -8 -3 16 105
use AND2X2  AND2X2_48
timestamp 1677677812
transform -1 0 3080 0 1 1770
box -8 -3 40 105
use FILL  FILL_7398
timestamp 1677677812
transform 1 0 3080 0 1 1770
box -8 -3 16 105
use FILL  FILL_7399
timestamp 1677677812
transform 1 0 3088 0 1 1770
box -8 -3 16 105
use FILL  FILL_7409
timestamp 1677677812
transform 1 0 3096 0 1 1770
box -8 -3 16 105
use FILL  FILL_7411
timestamp 1677677812
transform 1 0 3104 0 1 1770
box -8 -3 16 105
use FILL  FILL_7413
timestamp 1677677812
transform 1 0 3112 0 1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_51
timestamp 1677677812
transform -1 0 3152 0 1 1770
box -8 -3 40 105
use FILL  FILL_7414
timestamp 1677677812
transform 1 0 3152 0 1 1770
box -8 -3 16 105
use FILL  FILL_7417
timestamp 1677677812
transform 1 0 3160 0 1 1770
box -8 -3 16 105
use FILL  FILL_7419
timestamp 1677677812
transform 1 0 3168 0 1 1770
box -8 -3 16 105
use FILL  FILL_7420
timestamp 1677677812
transform 1 0 3176 0 1 1770
box -8 -3 16 105
use FILL  FILL_7421
timestamp 1677677812
transform 1 0 3184 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_460
timestamp 1677677812
transform -1 0 3208 0 1 1770
box -9 -3 26 105
use FILL  FILL_7422
timestamp 1677677812
transform 1 0 3208 0 1 1770
box -8 -3 16 105
use FILL  FILL_7425
timestamp 1677677812
transform 1 0 3216 0 1 1770
box -8 -3 16 105
use FILL  FILL_7427
timestamp 1677677812
transform 1 0 3224 0 1 1770
box -8 -3 16 105
use FILL  FILL_7429
timestamp 1677677812
transform 1 0 3232 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_90
timestamp 1677677812
transform 1 0 3240 0 1 1770
box -5 -3 28 105
use FILL  FILL_7430
timestamp 1677677812
transform 1 0 3264 0 1 1770
box -8 -3 16 105
use FILL  FILL_7432
timestamp 1677677812
transform 1 0 3272 0 1 1770
box -8 -3 16 105
use FILL  FILL_7434
timestamp 1677677812
transform 1 0 3280 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_461
timestamp 1677677812
transform 1 0 3288 0 1 1770
box -9 -3 26 105
use FILL  FILL_7435
timestamp 1677677812
transform 1 0 3304 0 1 1770
box -8 -3 16 105
use FILL  FILL_7436
timestamp 1677677812
transform 1 0 3312 0 1 1770
box -8 -3 16 105
use FILL  FILL_7437
timestamp 1677677812
transform 1 0 3320 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5426
timestamp 1677677812
transform 1 0 3340 0 1 1775
box -3 -3 3 3
use FILL  FILL_7438
timestamp 1677677812
transform 1 0 3328 0 1 1770
box -8 -3 16 105
use BUFX2  BUFX2_91
timestamp 1677677812
transform -1 0 3360 0 1 1770
box -5 -3 28 105
use FILL  FILL_7439
timestamp 1677677812
transform 1 0 3360 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5427
timestamp 1677677812
transform 1 0 3396 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_399
timestamp 1677677812
transform -1 0 3464 0 1 1770
box -8 -3 104 105
use FILL  FILL_7440
timestamp 1677677812
transform 1 0 3464 0 1 1770
box -8 -3 16 105
use FILL  FILL_7441
timestamp 1677677812
transform 1 0 3472 0 1 1770
box -8 -3 16 105
use FILL  FILL_7442
timestamp 1677677812
transform 1 0 3480 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_400
timestamp 1677677812
transform 1 0 3488 0 1 1770
box -8 -3 104 105
use FILL  FILL_7443
timestamp 1677677812
transform 1 0 3584 0 1 1770
box -8 -3 16 105
use FILL  FILL_7456
timestamp 1677677812
transform 1 0 3592 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_464
timestamp 1677677812
transform -1 0 3616 0 1 1770
box -9 -3 26 105
use FILL  FILL_7457
timestamp 1677677812
transform 1 0 3616 0 1 1770
box -8 -3 16 105
use FILL  FILL_7458
timestamp 1677677812
transform 1 0 3624 0 1 1770
box -8 -3 16 105
use FILL  FILL_7459
timestamp 1677677812
transform 1 0 3632 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_465
timestamp 1677677812
transform 1 0 3640 0 1 1770
box -9 -3 26 105
use FILL  FILL_7460
timestamp 1677677812
transform 1 0 3656 0 1 1770
box -8 -3 16 105
use FILL  FILL_7461
timestamp 1677677812
transform 1 0 3664 0 1 1770
box -8 -3 16 105
use FILL  FILL_7462
timestamp 1677677812
transform 1 0 3672 0 1 1770
box -8 -3 16 105
use FILL  FILL_7463
timestamp 1677677812
transform 1 0 3680 0 1 1770
box -8 -3 16 105
use FILL  FILL_7464
timestamp 1677677812
transform 1 0 3688 0 1 1770
box -8 -3 16 105
use FILL  FILL_7466
timestamp 1677677812
transform 1 0 3696 0 1 1770
box -8 -3 16 105
use FILL  FILL_7468
timestamp 1677677812
transform 1 0 3704 0 1 1770
box -8 -3 16 105
use FILL  FILL_7469
timestamp 1677677812
transform 1 0 3712 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_466
timestamp 1677677812
transform -1 0 3736 0 1 1770
box -9 -3 26 105
use FILL  FILL_7470
timestamp 1677677812
transform 1 0 3736 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5428
timestamp 1677677812
transform 1 0 3756 0 1 1775
box -3 -3 3 3
use FILL  FILL_7471
timestamp 1677677812
transform 1 0 3744 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5429
timestamp 1677677812
transform 1 0 3796 0 1 1775
box -3 -3 3 3
use OAI22X1  OAI22X1_263
timestamp 1677677812
transform 1 0 3752 0 1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_402
timestamp 1677677812
transform -1 0 3888 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_467
timestamp 1677677812
transform -1 0 3904 0 1 1770
box -9 -3 26 105
use FILL  FILL_7472
timestamp 1677677812
transform 1 0 3904 0 1 1770
box -8 -3 16 105
use FILL  FILL_7478
timestamp 1677677812
transform 1 0 3912 0 1 1770
box -8 -3 16 105
use FILL  FILL_7480
timestamp 1677677812
transform 1 0 3920 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5430
timestamp 1677677812
transform 1 0 3948 0 1 1775
box -3 -3 3 3
use INVX2  INVX2_470
timestamp 1677677812
transform -1 0 3944 0 1 1770
box -9 -3 26 105
use FILL  FILL_7481
timestamp 1677677812
transform 1 0 3944 0 1 1770
box -8 -3 16 105
use FILL  FILL_7482
timestamp 1677677812
transform 1 0 3952 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_265
timestamp 1677677812
transform 1 0 3960 0 1 1770
box -8 -3 46 105
use FILL  FILL_7483
timestamp 1677677812
transform 1 0 4000 0 1 1770
box -8 -3 16 105
use FILL  FILL_7488
timestamp 1677677812
transform 1 0 4008 0 1 1770
box -8 -3 16 105
use FILL  FILL_7489
timestamp 1677677812
transform 1 0 4016 0 1 1770
box -8 -3 16 105
use FILL  FILL_7490
timestamp 1677677812
transform 1 0 4024 0 1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5431
timestamp 1677677812
transform 1 0 4052 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5432
timestamp 1677677812
transform 1 0 4076 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5433
timestamp 1677677812
transform 1 0 4100 0 1 1775
box -3 -3 3 3
use M3_M2  M3_M2_5434
timestamp 1677677812
transform 1 0 4132 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_404
timestamp 1677677812
transform 1 0 4032 0 1 1770
box -8 -3 104 105
use FILL  FILL_7492
timestamp 1677677812
transform 1 0 4128 0 1 1770
box -8 -3 16 105
use FILL  FILL_7493
timestamp 1677677812
transform 1 0 4136 0 1 1770
box -8 -3 16 105
use FILL  FILL_7494
timestamp 1677677812
transform 1 0 4144 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_267
timestamp 1677677812
transform 1 0 4152 0 1 1770
box -8 -3 46 105
use FILL  FILL_7495
timestamp 1677677812
transform 1 0 4192 0 1 1770
box -8 -3 16 105
use FILL  FILL_7496
timestamp 1677677812
transform 1 0 4200 0 1 1770
box -8 -3 16 105
use FILL  FILL_7497
timestamp 1677677812
transform 1 0 4208 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_268
timestamp 1677677812
transform 1 0 4216 0 1 1770
box -8 -3 46 105
use FILL  FILL_7498
timestamp 1677677812
transform 1 0 4256 0 1 1770
box -8 -3 16 105
use FILL  FILL_7499
timestamp 1677677812
transform 1 0 4264 0 1 1770
box -8 -3 16 105
use INVX2  INVX2_473
timestamp 1677677812
transform -1 0 4288 0 1 1770
box -9 -3 26 105
use FILL  FILL_7500
timestamp 1677677812
transform 1 0 4288 0 1 1770
box -8 -3 16 105
use FILL  FILL_7508
timestamp 1677677812
transform 1 0 4296 0 1 1770
box -8 -3 16 105
use FILL  FILL_7510
timestamp 1677677812
transform 1 0 4304 0 1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_406
timestamp 1677677812
transform 1 0 4312 0 1 1770
box -8 -3 104 105
use FILL  FILL_7512
timestamp 1677677812
transform 1 0 4408 0 1 1770
box -8 -3 16 105
use FILL  FILL_7513
timestamp 1677677812
transform 1 0 4416 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_271
timestamp 1677677812
transform -1 0 4464 0 1 1770
box -8 -3 46 105
use FILL  FILL_7514
timestamp 1677677812
transform 1 0 4464 0 1 1770
box -8 -3 16 105
use FILL  FILL_7515
timestamp 1677677812
transform 1 0 4472 0 1 1770
box -8 -3 16 105
use FILL  FILL_7516
timestamp 1677677812
transform 1 0 4480 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_272
timestamp 1677677812
transform -1 0 4528 0 1 1770
box -8 -3 46 105
use M3_M2  M3_M2_5435
timestamp 1677677812
transform 1 0 4628 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_407
timestamp 1677677812
transform -1 0 4624 0 1 1770
box -8 -3 104 105
use FILL  FILL_7517
timestamp 1677677812
transform 1 0 4624 0 1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_276
timestamp 1677677812
transform 1 0 4632 0 1 1770
box -8 -3 46 105
use M3_M2  M3_M2_5436
timestamp 1677677812
transform 1 0 4732 0 1 1775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_408
timestamp 1677677812
transform 1 0 4672 0 1 1770
box -8 -3 104 105
use INVX2  INVX2_478
timestamp 1677677812
transform -1 0 4784 0 1 1770
box -9 -3 26 105
use FILL  FILL_7539
timestamp 1677677812
transform 1 0 4784 0 1 1770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_59
timestamp 1677677812
transform 1 0 4819 0 1 1770
box -10 -3 10 3
use M2_M1  M2_M1_6114
timestamp 1677677812
transform 1 0 92 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6219
timestamp 1677677812
transform 1 0 132 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6115
timestamp 1677677812
transform 1 0 180 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5473
timestamp 1677677812
transform 1 0 212 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5510
timestamp 1677677812
transform 1 0 204 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5474
timestamp 1677677812
transform 1 0 276 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5475
timestamp 1677677812
transform 1 0 356 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6116
timestamp 1677677812
transform 1 0 236 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6117
timestamp 1677677812
transform 1 0 244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6118
timestamp 1677677812
transform 1 0 260 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6119
timestamp 1677677812
transform 1 0 276 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5511
timestamp 1677677812
transform 1 0 300 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6220
timestamp 1677677812
transform 1 0 204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6221
timestamp 1677677812
transform 1 0 212 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6222
timestamp 1677677812
transform 1 0 228 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5536
timestamp 1677677812
transform 1 0 236 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6223
timestamp 1677677812
transform 1 0 244 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6224
timestamp 1677677812
transform 1 0 251 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5537
timestamp 1677677812
transform 1 0 260 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5538
timestamp 1677677812
transform 1 0 276 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5539
timestamp 1677677812
transform 1 0 308 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6225
timestamp 1677677812
transform 1 0 324 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6226
timestamp 1677677812
transform 1 0 356 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6227
timestamp 1677677812
transform 1 0 364 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6228
timestamp 1677677812
transform 1 0 372 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5569
timestamp 1677677812
transform 1 0 324 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5570
timestamp 1677677812
transform 1 0 364 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5646
timestamp 1677677812
transform 1 0 260 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5647
timestamp 1677677812
transform 1 0 316 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5648
timestamp 1677677812
transform 1 0 332 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5633
timestamp 1677677812
transform 1 0 372 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5476
timestamp 1677677812
transform 1 0 412 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6120
timestamp 1677677812
transform 1 0 388 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6121
timestamp 1677677812
transform 1 0 396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6122
timestamp 1677677812
transform 1 0 412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6229
timestamp 1677677812
transform 1 0 404 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6230
timestamp 1677677812
transform 1 0 420 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6231
timestamp 1677677812
transform 1 0 428 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5611
timestamp 1677677812
transform 1 0 428 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6123
timestamp 1677677812
transform 1 0 468 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5512
timestamp 1677677812
transform 1 0 476 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6124
timestamp 1677677812
transform 1 0 484 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6232
timestamp 1677677812
transform 1 0 476 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5540
timestamp 1677677812
transform 1 0 484 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6233
timestamp 1677677812
transform 1 0 492 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5541
timestamp 1677677812
transform 1 0 500 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6234
timestamp 1677677812
transform 1 0 540 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6125
timestamp 1677677812
transform 1 0 556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6126
timestamp 1677677812
transform 1 0 572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6127
timestamp 1677677812
transform 1 0 596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6235
timestamp 1677677812
transform 1 0 564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6236
timestamp 1677677812
transform 1 0 580 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5571
timestamp 1677677812
transform 1 0 556 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5634
timestamp 1677677812
transform 1 0 556 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5572
timestamp 1677677812
transform 1 0 580 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6128
timestamp 1677677812
transform 1 0 612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6237
timestamp 1677677812
transform 1 0 620 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6238
timestamp 1677677812
transform 1 0 628 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5612
timestamp 1677677812
transform 1 0 628 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5437
timestamp 1677677812
transform 1 0 644 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5448
timestamp 1677677812
transform 1 0 652 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6129
timestamp 1677677812
transform 1 0 652 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5513
timestamp 1677677812
transform 1 0 660 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5542
timestamp 1677677812
transform 1 0 644 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6239
timestamp 1677677812
transform 1 0 660 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5573
timestamp 1677677812
transform 1 0 660 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6130
timestamp 1677677812
transform 1 0 692 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5574
timestamp 1677677812
transform 1 0 692 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5477
timestamp 1677677812
transform 1 0 708 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5478
timestamp 1677677812
transform 1 0 796 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6131
timestamp 1677677812
transform 1 0 708 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5514
timestamp 1677677812
transform 1 0 772 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5515
timestamp 1677677812
transform 1 0 788 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6240
timestamp 1677677812
transform 1 0 740 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5543
timestamp 1677677812
transform 1 0 748 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6241
timestamp 1677677812
transform 1 0 788 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6242
timestamp 1677677812
transform 1 0 804 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5575
timestamp 1677677812
transform 1 0 788 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5613
timestamp 1677677812
transform 1 0 756 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5479
timestamp 1677677812
transform 1 0 828 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5576
timestamp 1677677812
transform 1 0 836 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5480
timestamp 1677677812
transform 1 0 876 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5449
timestamp 1677677812
transform 1 0 892 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6108
timestamp 1677677812
transform 1 0 892 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6132
timestamp 1677677812
transform 1 0 852 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6133
timestamp 1677677812
transform 1 0 860 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6134
timestamp 1677677812
transform 1 0 876 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6351
timestamp 1677677812
transform 1 0 844 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5516
timestamp 1677677812
transform 1 0 884 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5544
timestamp 1677677812
transform 1 0 860 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6243
timestamp 1677677812
transform 1 0 868 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6244
timestamp 1677677812
transform 1 0 892 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5614
timestamp 1677677812
transform 1 0 884 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5649
timestamp 1677677812
transform 1 0 876 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5481
timestamp 1677677812
transform 1 0 908 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6135
timestamp 1677677812
transform 1 0 964 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5545
timestamp 1677677812
transform 1 0 964 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5546
timestamp 1677677812
transform 1 0 1036 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5450
timestamp 1677677812
transform 1 0 1084 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5482
timestamp 1677677812
transform 1 0 1108 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5517
timestamp 1677677812
transform 1 0 1076 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6136
timestamp 1677677812
transform 1 0 1084 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5518
timestamp 1677677812
transform 1 0 1100 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6245
timestamp 1677677812
transform 1 0 1068 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6246
timestamp 1677677812
transform 1 0 1076 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6247
timestamp 1677677812
transform 1 0 1092 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6248
timestamp 1677677812
transform 1 0 1108 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5577
timestamp 1677677812
transform 1 0 1068 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5483
timestamp 1677677812
transform 1 0 1172 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5519
timestamp 1677677812
transform 1 0 1180 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5484
timestamp 1677677812
transform 1 0 1196 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6137
timestamp 1677677812
transform 1 0 1196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6249
timestamp 1677677812
transform 1 0 1188 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5438
timestamp 1677677812
transform 1 0 1228 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5520
timestamp 1677677812
transform 1 0 1220 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6138
timestamp 1677677812
transform 1 0 1228 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5547
timestamp 1677677812
transform 1 0 1204 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6250
timestamp 1677677812
transform 1 0 1220 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5615
timestamp 1677677812
transform 1 0 1228 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5451
timestamp 1677677812
transform 1 0 1244 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6251
timestamp 1677677812
transform 1 0 1244 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5452
timestamp 1677677812
transform 1 0 1268 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5485
timestamp 1677677812
transform 1 0 1260 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5578
timestamp 1677677812
transform 1 0 1268 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6252
timestamp 1677677812
transform 1 0 1308 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5616
timestamp 1677677812
transform 1 0 1308 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5453
timestamp 1677677812
transform 1 0 1324 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6139
timestamp 1677677812
transform 1 0 1324 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5521
timestamp 1677677812
transform 1 0 1332 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6253
timestamp 1677677812
transform 1 0 1324 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5650
timestamp 1677677812
transform 1 0 1324 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5486
timestamp 1677677812
transform 1 0 1396 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6140
timestamp 1677677812
transform 1 0 1396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6141
timestamp 1677677812
transform 1 0 1404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6254
timestamp 1677677812
transform 1 0 1388 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5617
timestamp 1677677812
transform 1 0 1388 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5651
timestamp 1677677812
transform 1 0 1372 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5652
timestamp 1677677812
transform 1 0 1388 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6255
timestamp 1677677812
transform 1 0 1404 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5487
timestamp 1677677812
transform 1 0 1420 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5488
timestamp 1677677812
transform 1 0 1436 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5439
timestamp 1677677812
transform 1 0 1460 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5489
timestamp 1677677812
transform 1 0 1476 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6142
timestamp 1677677812
transform 1 0 1452 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6143
timestamp 1677677812
transform 1 0 1476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6256
timestamp 1677677812
transform 1 0 1468 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5548
timestamp 1677677812
transform 1 0 1476 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6257
timestamp 1677677812
transform 1 0 1484 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5549
timestamp 1677677812
transform 1 0 1492 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6144
timestamp 1677677812
transform 1 0 1556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6258
timestamp 1677677812
transform 1 0 1548 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5618
timestamp 1677677812
transform 1 0 1548 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6145
timestamp 1677677812
transform 1 0 1588 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5550
timestamp 1677677812
transform 1 0 1580 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5579
timestamp 1677677812
transform 1 0 1588 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6259
timestamp 1677677812
transform 1 0 1604 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5551
timestamp 1677677812
transform 1 0 1620 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6260
timestamp 1677677812
transform 1 0 1700 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5440
timestamp 1677677812
transform 1 0 1748 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5454
timestamp 1677677812
transform 1 0 1732 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5490
timestamp 1677677812
transform 1 0 1748 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6146
timestamp 1677677812
transform 1 0 1716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6147
timestamp 1677677812
transform 1 0 1724 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6148
timestamp 1677677812
transform 1 0 1740 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6261
timestamp 1677677812
transform 1 0 1732 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6262
timestamp 1677677812
transform 1 0 1748 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5491
timestamp 1677677812
transform 1 0 1820 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5522
timestamp 1677677812
transform 1 0 1812 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6149
timestamp 1677677812
transform 1 0 1820 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6263
timestamp 1677677812
transform 1 0 1812 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6352
timestamp 1677677812
transform 1 0 1820 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6150
timestamp 1677677812
transform 1 0 1836 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6353
timestamp 1677677812
transform 1 0 1852 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5441
timestamp 1677677812
transform 1 0 1908 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5455
timestamp 1677677812
transform 1 0 1972 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6151
timestamp 1677677812
transform 1 0 1900 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6152
timestamp 1677677812
transform 1 0 1908 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6153
timestamp 1677677812
transform 1 0 1996 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6264
timestamp 1677677812
transform 1 0 1876 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6265
timestamp 1677677812
transform 1 0 1892 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6266
timestamp 1677677812
transform 1 0 1908 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6267
timestamp 1677677812
transform 1 0 1916 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6268
timestamp 1677677812
transform 1 0 1964 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5653
timestamp 1677677812
transform 1 0 1900 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5580
timestamp 1677677812
transform 1 0 1996 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5654
timestamp 1677677812
transform 1 0 1932 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5492
timestamp 1677677812
transform 1 0 2012 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6269
timestamp 1677677812
transform 1 0 2012 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5493
timestamp 1677677812
transform 1 0 2028 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5581
timestamp 1677677812
transform 1 0 2028 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5635
timestamp 1677677812
transform 1 0 2020 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5442
timestamp 1677677812
transform 1 0 2068 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6154
timestamp 1677677812
transform 1 0 2068 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6270
timestamp 1677677812
transform 1 0 2060 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5582
timestamp 1677677812
transform 1 0 2060 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6271
timestamp 1677677812
transform 1 0 2076 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5619
timestamp 1677677812
transform 1 0 2076 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5456
timestamp 1677677812
transform 1 0 2148 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6155
timestamp 1677677812
transform 1 0 2140 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6272
timestamp 1677677812
transform 1 0 2132 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5583
timestamp 1677677812
transform 1 0 2132 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5523
timestamp 1677677812
transform 1 0 2148 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6273
timestamp 1677677812
transform 1 0 2156 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6109
timestamp 1677677812
transform 1 0 2204 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6156
timestamp 1677677812
transform 1 0 2196 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6274
timestamp 1677677812
transform 1 0 2188 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6110
timestamp 1677677812
transform 1 0 2244 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_5494
timestamp 1677677812
transform 1 0 2252 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6111
timestamp 1677677812
transform 1 0 2268 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6157
timestamp 1677677812
transform 1 0 2244 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6158
timestamp 1677677812
transform 1 0 2252 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6159
timestamp 1677677812
transform 1 0 2260 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5524
timestamp 1677677812
transform 1 0 2268 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6275
timestamp 1677677812
transform 1 0 2260 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5636
timestamp 1677677812
transform 1 0 2252 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5495
timestamp 1677677812
transform 1 0 2284 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5525
timestamp 1677677812
transform 1 0 2292 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6276
timestamp 1677677812
transform 1 0 2284 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6277
timestamp 1677677812
transform 1 0 2292 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5584
timestamp 1677677812
transform 1 0 2300 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5496
timestamp 1677677812
transform 1 0 2348 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5443
timestamp 1677677812
transform 1 0 2380 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5497
timestamp 1677677812
transform 1 0 2372 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6160
timestamp 1677677812
transform 1 0 2364 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6161
timestamp 1677677812
transform 1 0 2372 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6278
timestamp 1677677812
transform 1 0 2356 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5444
timestamp 1677677812
transform 1 0 2404 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6279
timestamp 1677677812
transform 1 0 2380 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6280
timestamp 1677677812
transform 1 0 2396 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6281
timestamp 1677677812
transform 1 0 2404 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5526
timestamp 1677677812
transform 1 0 2436 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6162
timestamp 1677677812
transform 1 0 2444 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6282
timestamp 1677677812
transform 1 0 2428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6337
timestamp 1677677812
transform 1 0 2436 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5585
timestamp 1677677812
transform 1 0 2444 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6163
timestamp 1677677812
transform 1 0 2476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6283
timestamp 1677677812
transform 1 0 2484 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5586
timestamp 1677677812
transform 1 0 2484 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6338
timestamp 1677677812
transform 1 0 2492 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5457
timestamp 1677677812
transform 1 0 2508 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5552
timestamp 1677677812
transform 1 0 2532 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6284
timestamp 1677677812
transform 1 0 2540 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5587
timestamp 1677677812
transform 1 0 2540 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6354
timestamp 1677677812
transform 1 0 2532 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6164
timestamp 1677677812
transform 1 0 2564 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5527
timestamp 1677677812
transform 1 0 2604 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6165
timestamp 1677677812
transform 1 0 2612 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6285
timestamp 1677677812
transform 1 0 2572 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6286
timestamp 1677677812
transform 1 0 2596 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6339
timestamp 1677677812
transform 1 0 2580 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5637
timestamp 1677677812
transform 1 0 2564 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5588
timestamp 1677677812
transform 1 0 2596 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6355
timestamp 1677677812
transform 1 0 2588 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5553
timestamp 1677677812
transform 1 0 2612 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6287
timestamp 1677677812
transform 1 0 2628 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6288
timestamp 1677677812
transform 1 0 2652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6340
timestamp 1677677812
transform 1 0 2644 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5589
timestamp 1677677812
transform 1 0 2652 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5554
timestamp 1677677812
transform 1 0 2676 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6341
timestamp 1677677812
transform 1 0 2668 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6342
timestamp 1677677812
transform 1 0 2676 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5620
timestamp 1677677812
transform 1 0 2628 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5621
timestamp 1677677812
transform 1 0 2644 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6356
timestamp 1677677812
transform 1 0 2652 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5638
timestamp 1677677812
transform 1 0 2620 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5639
timestamp 1677677812
transform 1 0 2652 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6357
timestamp 1677677812
transform 1 0 2676 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5640
timestamp 1677677812
transform 1 0 2676 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6289
timestamp 1677677812
transform 1 0 2724 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5590
timestamp 1677677812
transform 1 0 2724 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6343
timestamp 1677677812
transform 1 0 2740 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6166
timestamp 1677677812
transform 1 0 2812 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6290
timestamp 1677677812
transform 1 0 2804 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6291
timestamp 1677677812
transform 1 0 2844 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5458
timestamp 1677677812
transform 1 0 2868 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6167
timestamp 1677677812
transform 1 0 2868 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5555
timestamp 1677677812
transform 1 0 2868 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5459
timestamp 1677677812
transform 1 0 2940 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6112
timestamp 1677677812
transform 1 0 2940 0 1 1745
box -2 -2 2 2
use M2_M1  M2_M1_6168
timestamp 1677677812
transform 1 0 2932 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5556
timestamp 1677677812
transform 1 0 2924 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5591
timestamp 1677677812
transform 1 0 2932 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6169
timestamp 1677677812
transform 1 0 2956 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6292
timestamp 1677677812
transform 1 0 2964 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6293
timestamp 1677677812
transform 1 0 2972 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5592
timestamp 1677677812
transform 1 0 2964 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6170
timestamp 1677677812
transform 1 0 3004 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6171
timestamp 1677677812
transform 1 0 3020 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5460
timestamp 1677677812
transform 1 0 3036 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6172
timestamp 1677677812
transform 1 0 3068 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6173
timestamp 1677677812
transform 1 0 3076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6294
timestamp 1677677812
transform 1 0 3060 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5557
timestamp 1677677812
transform 1 0 3068 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5593
timestamp 1677677812
transform 1 0 3068 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5461
timestamp 1677677812
transform 1 0 3100 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6295
timestamp 1677677812
transform 1 0 3084 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5558
timestamp 1677677812
transform 1 0 3092 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5594
timestamp 1677677812
transform 1 0 3084 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5641
timestamp 1677677812
transform 1 0 3076 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6358
timestamp 1677677812
transform 1 0 3092 0 1 1705
box -2 -2 2 2
use M2_M1  M2_M1_6344
timestamp 1677677812
transform 1 0 3100 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6296
timestamp 1677677812
transform 1 0 3124 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5595
timestamp 1677677812
transform 1 0 3124 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6345
timestamp 1677677812
transform 1 0 3140 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5596
timestamp 1677677812
transform 1 0 3148 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5622
timestamp 1677677812
transform 1 0 3140 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6359
timestamp 1677677812
transform 1 0 3148 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5559
timestamp 1677677812
transform 1 0 3172 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6297
timestamp 1677677812
transform 1 0 3180 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6346
timestamp 1677677812
transform 1 0 3164 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5597
timestamp 1677677812
transform 1 0 3180 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6360
timestamp 1677677812
transform 1 0 3172 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5623
timestamp 1677677812
transform 1 0 3188 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5462
timestamp 1677677812
transform 1 0 3204 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5560
timestamp 1677677812
transform 1 0 3212 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6347
timestamp 1677677812
transform 1 0 3204 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6348
timestamp 1677677812
transform 1 0 3212 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6361
timestamp 1677677812
transform 1 0 3212 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5642
timestamp 1677677812
transform 1 0 3212 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6362
timestamp 1677677812
transform 1 0 3228 0 1 1705
box -2 -2 2 2
use M3_M2  M3_M2_5463
timestamp 1677677812
transform 1 0 3260 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6298
timestamp 1677677812
transform 1 0 3244 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5598
timestamp 1677677812
transform 1 0 3244 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5561
timestamp 1677677812
transform 1 0 3284 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6349
timestamp 1677677812
transform 1 0 3284 0 1 1715
box -2 -2 2 2
use M2_M1  M2_M1_6113
timestamp 1677677812
transform 1 0 3300 0 1 1745
box -2 -2 2 2
use M3_M2  M3_M2_5498
timestamp 1677677812
transform 1 0 3404 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6174
timestamp 1677677812
transform 1 0 3404 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6175
timestamp 1677677812
transform 1 0 3412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6299
timestamp 1677677812
transform 1 0 3388 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6300
timestamp 1677677812
transform 1 0 3396 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5562
timestamp 1677677812
transform 1 0 3412 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5499
timestamp 1677677812
transform 1 0 3436 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6176
timestamp 1677677812
transform 1 0 3436 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6301
timestamp 1677677812
transform 1 0 3428 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6302
timestamp 1677677812
transform 1 0 3436 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5599
timestamp 1677677812
transform 1 0 3428 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5624
timestamp 1677677812
transform 1 0 3436 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6177
timestamp 1677677812
transform 1 0 3476 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5528
timestamp 1677677812
transform 1 0 3484 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6303
timestamp 1677677812
transform 1 0 3468 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6304
timestamp 1677677812
transform 1 0 3484 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6178
timestamp 1677677812
transform 1 0 3500 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6305
timestamp 1677677812
transform 1 0 3500 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5500
timestamp 1677677812
transform 1 0 3516 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6179
timestamp 1677677812
transform 1 0 3516 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6306
timestamp 1677677812
transform 1 0 3516 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5600
timestamp 1677677812
transform 1 0 3524 0 1 1715
box -3 -3 3 3
use M2_M1  M2_M1_6307
timestamp 1677677812
transform 1 0 3548 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6180
timestamp 1677677812
transform 1 0 3572 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6181
timestamp 1677677812
transform 1 0 3588 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5464
timestamp 1677677812
transform 1 0 3604 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5501
timestamp 1677677812
transform 1 0 3668 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6182
timestamp 1677677812
transform 1 0 3604 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5529
timestamp 1677677812
transform 1 0 3652 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5563
timestamp 1677677812
transform 1 0 3604 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6308
timestamp 1677677812
transform 1 0 3652 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6350
timestamp 1677677812
transform 1 0 3724 0 1 1715
box -2 -2 2 2
use M3_M2  M3_M2_5465
timestamp 1677677812
transform 1 0 3740 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6183
timestamp 1677677812
transform 1 0 3740 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5530
timestamp 1677677812
transform 1 0 3748 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6184
timestamp 1677677812
transform 1 0 3756 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6309
timestamp 1677677812
transform 1 0 3764 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5445
timestamp 1677677812
transform 1 0 3780 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6310
timestamp 1677677812
transform 1 0 3780 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5502
timestamp 1677677812
transform 1 0 3788 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6185
timestamp 1677677812
transform 1 0 3788 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6186
timestamp 1677677812
transform 1 0 3796 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6187
timestamp 1677677812
transform 1 0 3820 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5531
timestamp 1677677812
transform 1 0 3868 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6311
timestamp 1677677812
transform 1 0 3804 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5564
timestamp 1677677812
transform 1 0 3820 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6312
timestamp 1677677812
transform 1 0 3868 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5466
timestamp 1677677812
transform 1 0 3956 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5503
timestamp 1677677812
transform 1 0 3988 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6188
timestamp 1677677812
transform 1 0 3956 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5532
timestamp 1677677812
transform 1 0 3964 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6189
timestamp 1677677812
transform 1 0 3972 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6190
timestamp 1677677812
transform 1 0 3988 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6313
timestamp 1677677812
transform 1 0 3948 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6314
timestamp 1677677812
transform 1 0 3980 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5643
timestamp 1677677812
transform 1 0 3980 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5625
timestamp 1677677812
transform 1 0 3996 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5467
timestamp 1677677812
transform 1 0 4012 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6191
timestamp 1677677812
transform 1 0 4012 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5533
timestamp 1677677812
transform 1 0 4044 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5468
timestamp 1677677812
transform 1 0 4076 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6192
timestamp 1677677812
transform 1 0 4060 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6193
timestamp 1677677812
transform 1 0 4076 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6315
timestamp 1677677812
transform 1 0 4052 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6316
timestamp 1677677812
transform 1 0 4068 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5655
timestamp 1677677812
transform 1 0 4052 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5504
timestamp 1677677812
transform 1 0 4108 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5469
timestamp 1677677812
transform 1 0 4132 0 1 1755
box -3 -3 3 3
use M3_M2  M3_M2_5505
timestamp 1677677812
transform 1 0 4164 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6194
timestamp 1677677812
transform 1 0 4124 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6195
timestamp 1677677812
transform 1 0 4132 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6196
timestamp 1677677812
transform 1 0 4148 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5534
timestamp 1677677812
transform 1 0 4156 0 1 1735
box -3 -3 3 3
use M2_M1  M2_M1_6197
timestamp 1677677812
transform 1 0 4164 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6198
timestamp 1677677812
transform 1 0 4180 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6317
timestamp 1677677812
transform 1 0 4140 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5565
timestamp 1677677812
transform 1 0 4148 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6318
timestamp 1677677812
transform 1 0 4156 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5601
timestamp 1677677812
transform 1 0 4140 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5626
timestamp 1677677812
transform 1 0 4156 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5535
timestamp 1677677812
transform 1 0 4204 0 1 1735
box -3 -3 3 3
use M3_M2  M3_M2_5566
timestamp 1677677812
transform 1 0 4180 0 1 1725
box -3 -3 3 3
use M2_M1  M2_M1_6199
timestamp 1677677812
transform 1 0 4276 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6319
timestamp 1677677812
transform 1 0 4204 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6320
timestamp 1677677812
transform 1 0 4260 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6321
timestamp 1677677812
transform 1 0 4268 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5602
timestamp 1677677812
transform 1 0 4268 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5627
timestamp 1677677812
transform 1 0 4212 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5656
timestamp 1677677812
transform 1 0 4204 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5470
timestamp 1677677812
transform 1 0 4332 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6200
timestamp 1677677812
transform 1 0 4332 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6201
timestamp 1677677812
transform 1 0 4348 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6322
timestamp 1677677812
transform 1 0 4332 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6323
timestamp 1677677812
transform 1 0 4356 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5603
timestamp 1677677812
transform 1 0 4332 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5644
timestamp 1677677812
transform 1 0 4356 0 1 1695
box -3 -3 3 3
use M2_M1  M2_M1_6324
timestamp 1677677812
transform 1 0 4372 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5604
timestamp 1677677812
transform 1 0 4372 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5506
timestamp 1677677812
transform 1 0 4396 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6202
timestamp 1677677812
transform 1 0 4396 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6203
timestamp 1677677812
transform 1 0 4412 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6325
timestamp 1677677812
transform 1 0 4404 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5471
timestamp 1677677812
transform 1 0 4428 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6204
timestamp 1677677812
transform 1 0 4428 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5507
timestamp 1677677812
transform 1 0 4476 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6205
timestamp 1677677812
transform 1 0 4460 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6206
timestamp 1677677812
transform 1 0 4476 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6326
timestamp 1677677812
transform 1 0 4444 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6327
timestamp 1677677812
transform 1 0 4468 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5605
timestamp 1677677812
transform 1 0 4444 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5645
timestamp 1677677812
transform 1 0 4436 0 1 1695
box -3 -3 3 3
use M3_M2  M3_M2_5628
timestamp 1677677812
transform 1 0 4468 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6328
timestamp 1677677812
transform 1 0 4484 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5606
timestamp 1677677812
transform 1 0 4484 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5629
timestamp 1677677812
transform 1 0 4500 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6207
timestamp 1677677812
transform 1 0 4532 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6208
timestamp 1677677812
transform 1 0 4556 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6209
timestamp 1677677812
transform 1 0 4572 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5472
timestamp 1677677812
transform 1 0 4604 0 1 1755
box -3 -3 3 3
use M2_M1  M2_M1_6210
timestamp 1677677812
transform 1 0 4596 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6211
timestamp 1677677812
transform 1 0 4604 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6329
timestamp 1677677812
transform 1 0 4564 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6330
timestamp 1677677812
transform 1 0 4580 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6331
timestamp 1677677812
transform 1 0 4588 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5607
timestamp 1677677812
transform 1 0 4556 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5608
timestamp 1677677812
transform 1 0 4588 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5630
timestamp 1677677812
transform 1 0 4596 0 1 1705
box -3 -3 3 3
use M2_M1  M2_M1_6332
timestamp 1677677812
transform 1 0 4628 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5609
timestamp 1677677812
transform 1 0 4628 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5446
timestamp 1677677812
transform 1 0 4660 0 1 1765
box -3 -3 3 3
use M3_M2  M3_M2_5508
timestamp 1677677812
transform 1 0 4652 0 1 1745
box -3 -3 3 3
use M3_M2  M3_M2_5509
timestamp 1677677812
transform 1 0 4676 0 1 1745
box -3 -3 3 3
use M2_M1  M2_M1_6218
timestamp 1677677812
transform 1 0 4644 0 1 1733
box -2 -2 2 2
use M2_M1  M2_M1_6212
timestamp 1677677812
transform 1 0 4660 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6213
timestamp 1677677812
transform 1 0 4676 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6214
timestamp 1677677812
transform 1 0 4684 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6333
timestamp 1677677812
transform 1 0 4668 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5657
timestamp 1677677812
transform 1 0 4668 0 1 1685
box -3 -3 3 3
use M3_M2  M3_M2_5447
timestamp 1677677812
transform 1 0 4700 0 1 1765
box -3 -3 3 3
use M2_M1  M2_M1_6215
timestamp 1677677812
transform 1 0 4716 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6216
timestamp 1677677812
transform 1 0 4732 0 1 1735
box -2 -2 2 2
use M2_M1  M2_M1_6334
timestamp 1677677812
transform 1 0 4708 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6335
timestamp 1677677812
transform 1 0 4724 0 1 1725
box -2 -2 2 2
use M2_M1  M2_M1_6336
timestamp 1677677812
transform 1 0 4732 0 1 1725
box -2 -2 2 2
use M3_M2  M3_M2_5567
timestamp 1677677812
transform 1 0 4740 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5610
timestamp 1677677812
transform 1 0 4732 0 1 1715
box -3 -3 3 3
use M3_M2  M3_M2_5631
timestamp 1677677812
transform 1 0 4724 0 1 1705
box -3 -3 3 3
use M3_M2  M3_M2_5658
timestamp 1677677812
transform 1 0 4708 0 1 1685
box -3 -3 3 3
use M2_M1  M2_M1_6217
timestamp 1677677812
transform 1 0 4764 0 1 1735
box -2 -2 2 2
use M3_M2  M3_M2_5568
timestamp 1677677812
transform 1 0 4764 0 1 1725
box -3 -3 3 3
use M3_M2  M3_M2_5632
timestamp 1677677812
transform 1 0 4772 0 1 1705
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_60
timestamp 1677677812
transform 1 0 24 0 1 1670
box -10 -3 10 3
use FILL  FILL_7079
timestamp 1677677812
transform 1 0 72 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_388
timestamp 1677677812
transform 1 0 80 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7080
timestamp 1677677812
transform 1 0 176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7081
timestamp 1677677812
transform 1 0 184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7082
timestamp 1677677812
transform 1 0 192 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7083
timestamp 1677677812
transform 1 0 200 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5659
timestamp 1677677812
transform 1 0 220 0 1 1675
box -3 -3 3 3
use M3_M2  M3_M2_5660
timestamp 1677677812
transform 1 0 244 0 1 1675
box -3 -3 3 3
use AOI22X1  AOI22X1_273
timestamp 1677677812
transform -1 0 248 0 -1 1770
box -8 -3 46 105
use INVX2  INVX2_440
timestamp 1677677812
transform -1 0 264 0 -1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_389
timestamp 1677677812
transform 1 0 264 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_441
timestamp 1677677812
transform -1 0 376 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7084
timestamp 1677677812
transform 1 0 376 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_275
timestamp 1677677812
transform 1 0 384 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7086
timestamp 1677677812
transform 1 0 424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7088
timestamp 1677677812
transform 1 0 432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7091
timestamp 1677677812
transform 1 0 440 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_257
timestamp 1677677812
transform 1 0 448 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7092
timestamp 1677677812
transform 1 0 488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7093
timestamp 1677677812
transform 1 0 496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7094
timestamp 1677677812
transform 1 0 504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7095
timestamp 1677677812
transform 1 0 512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7096
timestamp 1677677812
transform 1 0 520 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_442
timestamp 1677677812
transform -1 0 544 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7097
timestamp 1677677812
transform 1 0 544 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5661
timestamp 1677677812
transform 1 0 564 0 1 1675
box -3 -3 3 3
use FILL  FILL_7099
timestamp 1677677812
transform 1 0 552 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_276
timestamp 1677677812
transform 1 0 560 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7106
timestamp 1677677812
transform 1 0 600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7108
timestamp 1677677812
transform 1 0 608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7113
timestamp 1677677812
transform 1 0 616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7114
timestamp 1677677812
transform 1 0 624 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_258
timestamp 1677677812
transform 1 0 632 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7115
timestamp 1677677812
transform 1 0 672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7117
timestamp 1677677812
transform 1 0 680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7119
timestamp 1677677812
transform 1 0 688 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_392
timestamp 1677677812
transform 1 0 696 0 -1 1770
box -8 -3 104 105
use M3_M2  M3_M2_5662
timestamp 1677677812
transform 1 0 812 0 1 1675
box -3 -3 3 3
use INVX2  INVX2_443
timestamp 1677677812
transform -1 0 808 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7128
timestamp 1677677812
transform 1 0 808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7129
timestamp 1677677812
transform 1 0 816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7130
timestamp 1677677812
transform 1 0 824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7131
timestamp 1677677812
transform 1 0 832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7132
timestamp 1677677812
transform 1 0 840 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5663
timestamp 1677677812
transform 1 0 892 0 1 1675
box -3 -3 3 3
use AOI22X1  AOI22X1_277
timestamp 1677677812
transform -1 0 888 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7133
timestamp 1677677812
transform 1 0 888 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7134
timestamp 1677677812
transform 1 0 896 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7135
timestamp 1677677812
transform 1 0 904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7136
timestamp 1677677812
transform 1 0 912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7138
timestamp 1677677812
transform 1 0 920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7140
timestamp 1677677812
transform 1 0 928 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_66
timestamp 1677677812
transform 1 0 936 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7146
timestamp 1677677812
transform 1 0 960 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7147
timestamp 1677677812
transform 1 0 968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7148
timestamp 1677677812
transform 1 0 976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7149
timestamp 1677677812
transform 1 0 984 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7150
timestamp 1677677812
transform 1 0 992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7151
timestamp 1677677812
transform 1 0 1000 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7152
timestamp 1677677812
transform 1 0 1008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7154
timestamp 1677677812
transform 1 0 1016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7156
timestamp 1677677812
transform 1 0 1024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7158
timestamp 1677677812
transform 1 0 1032 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7160
timestamp 1677677812
transform 1 0 1040 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7162
timestamp 1677677812
transform 1 0 1048 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7168
timestamp 1677677812
transform 1 0 1056 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5664
timestamp 1677677812
transform 1 0 1076 0 1 1675
box -3 -3 3 3
use FILL  FILL_7169
timestamp 1677677812
transform 1 0 1064 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_279
timestamp 1677677812
transform 1 0 1072 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7170
timestamp 1677677812
transform 1 0 1112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7172
timestamp 1677677812
transform 1 0 1120 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7174
timestamp 1677677812
transform 1 0 1128 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7175
timestamp 1677677812
transform 1 0 1136 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7176
timestamp 1677677812
transform 1 0 1144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7178
timestamp 1677677812
transform 1 0 1152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7180
timestamp 1677677812
transform 1 0 1160 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7181
timestamp 1677677812
transform 1 0 1168 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7182
timestamp 1677677812
transform 1 0 1176 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7183
timestamp 1677677812
transform 1 0 1184 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7184
timestamp 1677677812
transform 1 0 1192 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_31
timestamp 1677677812
transform -1 0 1232 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7185
timestamp 1677677812
transform 1 0 1232 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7186
timestamp 1677677812
transform 1 0 1240 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7187
timestamp 1677677812
transform 1 0 1248 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7188
timestamp 1677677812
transform 1 0 1256 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7190
timestamp 1677677812
transform 1 0 1264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7192
timestamp 1677677812
transform 1 0 1272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7197
timestamp 1677677812
transform 1 0 1280 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_32
timestamp 1677677812
transform -1 0 1320 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7198
timestamp 1677677812
transform 1 0 1320 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7199
timestamp 1677677812
transform 1 0 1328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7200
timestamp 1677677812
transform 1 0 1336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7201
timestamp 1677677812
transform 1 0 1344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7203
timestamp 1677677812
transform 1 0 1352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7210
timestamp 1677677812
transform 1 0 1360 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_34
timestamp 1677677812
transform -1 0 1400 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7211
timestamp 1677677812
transform 1 0 1400 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7212
timestamp 1677677812
transform 1 0 1408 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7213
timestamp 1677677812
transform 1 0 1416 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5665
timestamp 1677677812
transform 1 0 1436 0 1 1675
box -3 -3 3 3
use FILL  FILL_7214
timestamp 1677677812
transform 1 0 1424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7215
timestamp 1677677812
transform 1 0 1432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7220
timestamp 1677677812
transform 1 0 1440 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_280
timestamp 1677677812
transform -1 0 1488 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7221
timestamp 1677677812
transform 1 0 1488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7222
timestamp 1677677812
transform 1 0 1496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7223
timestamp 1677677812
transform 1 0 1504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7224
timestamp 1677677812
transform 1 0 1512 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7225
timestamp 1677677812
transform 1 0 1520 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_35
timestamp 1677677812
transform -1 0 1560 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7226
timestamp 1677677812
transform 1 0 1560 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7228
timestamp 1677677812
transform 1 0 1568 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7229
timestamp 1677677812
transform 1 0 1576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7230
timestamp 1677677812
transform 1 0 1584 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7231
timestamp 1677677812
transform 1 0 1592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7232
timestamp 1677677812
transform 1 0 1600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7233
timestamp 1677677812
transform 1 0 1608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7234
timestamp 1677677812
transform 1 0 1616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7235
timestamp 1677677812
transform 1 0 1624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7236
timestamp 1677677812
transform 1 0 1632 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7237
timestamp 1677677812
transform 1 0 1640 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_445
timestamp 1677677812
transform -1 0 1664 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7238
timestamp 1677677812
transform 1 0 1664 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7240
timestamp 1677677812
transform 1 0 1672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7242
timestamp 1677677812
transform 1 0 1680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7244
timestamp 1677677812
transform 1 0 1688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7248
timestamp 1677677812
transform 1 0 1696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7249
timestamp 1677677812
transform 1 0 1704 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_281
timestamp 1677677812
transform -1 0 1752 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7250
timestamp 1677677812
transform 1 0 1752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7252
timestamp 1677677812
transform 1 0 1760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7254
timestamp 1677677812
transform 1 0 1768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7267
timestamp 1677677812
transform 1 0 1776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7268
timestamp 1677677812
transform 1 0 1784 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_36
timestamp 1677677812
transform -1 0 1824 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7269
timestamp 1677677812
transform 1 0 1824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7270
timestamp 1677677812
transform 1 0 1832 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5666
timestamp 1677677812
transform 1 0 1852 0 1 1675
box -3 -3 3 3
use FILL  FILL_7271
timestamp 1677677812
transform 1 0 1840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7272
timestamp 1677677812
transform 1 0 1848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7273
timestamp 1677677812
transform 1 0 1856 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7274
timestamp 1677677812
transform 1 0 1864 0 -1 1770
box -8 -3 16 105
use AOI22X1  AOI22X1_282
timestamp 1677677812
transform -1 0 1912 0 -1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_397
timestamp 1677677812
transform -1 0 2008 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7275
timestamp 1677677812
transform 1 0 2008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7277
timestamp 1677677812
transform 1 0 2016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7281
timestamp 1677677812
transform 1 0 2024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7282
timestamp 1677677812
transform 1 0 2032 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_38
timestamp 1677677812
transform -1 0 2072 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7283
timestamp 1677677812
transform 1 0 2072 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7285
timestamp 1677677812
transform 1 0 2080 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7287
timestamp 1677677812
transform 1 0 2088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7291
timestamp 1677677812
transform 1 0 2096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7292
timestamp 1677677812
transform 1 0 2104 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_40
timestamp 1677677812
transform -1 0 2144 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7293
timestamp 1677677812
transform 1 0 2144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7295
timestamp 1677677812
transform 1 0 2152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7297
timestamp 1677677812
transform 1 0 2160 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_42
timestamp 1677677812
transform -1 0 2200 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7299
timestamp 1677677812
transform 1 0 2200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7301
timestamp 1677677812
transform 1 0 2208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7303
timestamp 1677677812
transform 1 0 2216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7305
timestamp 1677677812
transform 1 0 2224 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7307
timestamp 1677677812
transform 1 0 2232 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_69
timestamp 1677677812
transform 1 0 2240 0 -1 1770
box -8 -3 32 105
use NOR2X1  NOR2X1_70
timestamp 1677677812
transform 1 0 2264 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7315
timestamp 1677677812
transform 1 0 2288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7316
timestamp 1677677812
transform 1 0 2296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7317
timestamp 1677677812
transform 1 0 2304 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_450
timestamp 1677677812
transform -1 0 2328 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7318
timestamp 1677677812
transform 1 0 2328 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7320
timestamp 1677677812
transform 1 0 2336 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7326
timestamp 1677677812
transform 1 0 2344 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7327
timestamp 1677677812
transform 1 0 2352 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7328
timestamp 1677677812
transform 1 0 2360 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_45
timestamp 1677677812
transform 1 0 2368 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7329
timestamp 1677677812
transform 1 0 2400 0 -1 1770
box -8 -3 16 105
use AND2X2  AND2X2_46
timestamp 1677677812
transform -1 0 2440 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7330
timestamp 1677677812
transform 1 0 2440 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_451
timestamp 1677677812
transform 1 0 2448 0 -1 1770
box -9 -3 26 105
use NOR2X1  NOR2X1_71
timestamp 1677677812
transform 1 0 2464 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7333
timestamp 1677677812
transform 1 0 2488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7335
timestamp 1677677812
transform 1 0 2496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7337
timestamp 1677677812
transform 1 0 2504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7342
timestamp 1677677812
transform 1 0 2512 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_47
timestamp 1677677812
transform -1 0 2552 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7343
timestamp 1677677812
transform 1 0 2552 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_453
timestamp 1677677812
transform 1 0 2560 0 -1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_48
timestamp 1677677812
transform -1 0 2608 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7347
timestamp 1677677812
transform 1 0 2608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7348
timestamp 1677677812
transform 1 0 2616 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_454
timestamp 1677677812
transform 1 0 2624 0 -1 1770
box -9 -3 26 105
use NAND3X1  NAND3X1_49
timestamp 1677677812
transform 1 0 2640 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7349
timestamp 1677677812
transform 1 0 2672 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7351
timestamp 1677677812
transform 1 0 2680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7353
timestamp 1677677812
transform 1 0 2688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7355
timestamp 1677677812
transform 1 0 2696 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7357
timestamp 1677677812
transform 1 0 2704 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_50
timestamp 1677677812
transform 1 0 2712 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7361
timestamp 1677677812
transform 1 0 2744 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7363
timestamp 1677677812
transform 1 0 2752 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7365
timestamp 1677677812
transform 1 0 2760 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7367
timestamp 1677677812
transform 1 0 2768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7369
timestamp 1677677812
transform 1 0 2776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7373
timestamp 1677677812
transform 1 0 2784 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_456
timestamp 1677677812
transform -1 0 2808 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7374
timestamp 1677677812
transform 1 0 2808 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7375
timestamp 1677677812
transform 1 0 2816 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7376
timestamp 1677677812
transform 1 0 2824 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7378
timestamp 1677677812
transform 1 0 2832 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7380
timestamp 1677677812
transform 1 0 2840 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7382
timestamp 1677677812
transform 1 0 2848 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7388
timestamp 1677677812
transform 1 0 2856 0 -1 1770
box -8 -3 16 105
use XNOR2X1  XNOR2X1_0
timestamp 1677677812
transform -1 0 2920 0 -1 1770
box -8 -3 64 105
use FILL  FILL_7389
timestamp 1677677812
transform 1 0 2920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7390
timestamp 1677677812
transform 1 0 2928 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7392
timestamp 1677677812
transform 1 0 2936 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_72
timestamp 1677677812
transform 1 0 2944 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7400
timestamp 1677677812
transform 1 0 2968 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7401
timestamp 1677677812
transform 1 0 2976 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7402
timestamp 1677677812
transform 1 0 2984 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_458
timestamp 1677677812
transform -1 0 3008 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7403
timestamp 1677677812
transform 1 0 3008 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7404
timestamp 1677677812
transform 1 0 3016 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7405
timestamp 1677677812
transform 1 0 3024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7406
timestamp 1677677812
transform 1 0 3032 0 -1 1770
box -8 -3 16 105
use NOR2X1  NOR2X1_73
timestamp 1677677812
transform 1 0 3040 0 -1 1770
box -8 -3 32 105
use FILL  FILL_7407
timestamp 1677677812
transform 1 0 3064 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_459
timestamp 1677677812
transform 1 0 3072 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7408
timestamp 1677677812
transform 1 0 3088 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7410
timestamp 1677677812
transform 1 0 3096 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7412
timestamp 1677677812
transform 1 0 3104 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_52
timestamp 1677677812
transform 1 0 3112 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7415
timestamp 1677677812
transform 1 0 3144 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7416
timestamp 1677677812
transform 1 0 3152 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7418
timestamp 1677677812
transform 1 0 3160 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_53
timestamp 1677677812
transform 1 0 3168 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7423
timestamp 1677677812
transform 1 0 3200 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7424
timestamp 1677677812
transform 1 0 3208 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7426
timestamp 1677677812
transform 1 0 3216 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7428
timestamp 1677677812
transform 1 0 3224 0 -1 1770
box -8 -3 16 105
use NAND3X1  NAND3X1_54
timestamp 1677677812
transform 1 0 3232 0 -1 1770
box -8 -3 40 105
use FILL  FILL_7431
timestamp 1677677812
transform 1 0 3264 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7433
timestamp 1677677812
transform 1 0 3272 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7444
timestamp 1677677812
transform 1 0 3280 0 -1 1770
box -8 -3 16 105
use FAX1  FAX1_0
timestamp 1677677812
transform -1 0 3408 0 -1 1770
box -5 -3 126 105
use FILL  FILL_7445
timestamp 1677677812
transform 1 0 3408 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_462
timestamp 1677677812
transform 1 0 3416 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7446
timestamp 1677677812
transform 1 0 3432 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7447
timestamp 1677677812
transform 1 0 3440 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7448
timestamp 1677677812
transform 1 0 3448 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_262
timestamp 1677677812
transform 1 0 3456 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7449
timestamp 1677677812
transform 1 0 3496 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_463
timestamp 1677677812
transform -1 0 3520 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7450
timestamp 1677677812
transform 1 0 3520 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7451
timestamp 1677677812
transform 1 0 3528 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7452
timestamp 1677677812
transform 1 0 3536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7453
timestamp 1677677812
transform 1 0 3544 0 -1 1770
box -8 -3 16 105
use M3_M2  M3_M2_5667
timestamp 1677677812
transform 1 0 3572 0 1 1675
box -3 -3 3 3
use BUFX2  BUFX2_92
timestamp 1677677812
transform 1 0 3552 0 -1 1770
box -5 -3 28 105
use FILL  FILL_7454
timestamp 1677677812
transform 1 0 3576 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7455
timestamp 1677677812
transform 1 0 3584 0 -1 1770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_401
timestamp 1677677812
transform 1 0 3592 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7465
timestamp 1677677812
transform 1 0 3688 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7467
timestamp 1677677812
transform 1 0 3696 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_468
timestamp 1677677812
transform 1 0 3704 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7473
timestamp 1677677812
transform 1 0 3720 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7474
timestamp 1677677812
transform 1 0 3728 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_264
timestamp 1677677812
transform 1 0 3736 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7475
timestamp 1677677812
transform 1 0 3776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7476
timestamp 1677677812
transform 1 0 3784 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_469
timestamp 1677677812
transform 1 0 3792 0 -1 1770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_403
timestamp 1677677812
transform 1 0 3808 0 -1 1770
box -8 -3 104 105
use FILL  FILL_7477
timestamp 1677677812
transform 1 0 3904 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7479
timestamp 1677677812
transform 1 0 3912 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7484
timestamp 1677677812
transform 1 0 3920 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7485
timestamp 1677677812
transform 1 0 3928 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_471
timestamp 1677677812
transform 1 0 3936 0 -1 1770
box -9 -3 26 105
use OAI22X1  OAI22X1_266
timestamp 1677677812
transform 1 0 3952 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7486
timestamp 1677677812
transform 1 0 3992 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7487
timestamp 1677677812
transform 1 0 4000 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_472
timestamp 1677677812
transform 1 0 4008 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7491
timestamp 1677677812
transform 1 0 4024 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7501
timestamp 1677677812
transform 1 0 4032 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_269
timestamp 1677677812
transform -1 0 4080 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7502
timestamp 1677677812
transform 1 0 4080 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_474
timestamp 1677677812
transform -1 0 4104 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7503
timestamp 1677677812
transform 1 0 4104 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7504
timestamp 1677677812
transform 1 0 4112 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7505
timestamp 1677677812
transform 1 0 4120 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_270
timestamp 1677677812
transform 1 0 4128 0 -1 1770
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_405
timestamp 1677677812
transform 1 0 4168 0 -1 1770
box -8 -3 104 105
use INVX2  INVX2_475
timestamp 1677677812
transform -1 0 4280 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7506
timestamp 1677677812
transform 1 0 4280 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7507
timestamp 1677677812
transform 1 0 4288 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7509
timestamp 1677677812
transform 1 0 4296 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7511
timestamp 1677677812
transform 1 0 4304 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7518
timestamp 1677677812
transform 1 0 4312 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7519
timestamp 1677677812
transform 1 0 4320 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_273
timestamp 1677677812
transform 1 0 4328 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7520
timestamp 1677677812
transform 1 0 4368 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7521
timestamp 1677677812
transform 1 0 4376 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7522
timestamp 1677677812
transform 1 0 4384 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7523
timestamp 1677677812
transform 1 0 4392 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_476
timestamp 1677677812
transform -1 0 4416 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7524
timestamp 1677677812
transform 1 0 4416 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7525
timestamp 1677677812
transform 1 0 4424 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7526
timestamp 1677677812
transform 1 0 4432 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_274
timestamp 1677677812
transform 1 0 4440 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7527
timestamp 1677677812
transform 1 0 4480 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7528
timestamp 1677677812
transform 1 0 4488 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7529
timestamp 1677677812
transform 1 0 4496 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7530
timestamp 1677677812
transform 1 0 4504 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7531
timestamp 1677677812
transform 1 0 4512 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_477
timestamp 1677677812
transform -1 0 4536 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7532
timestamp 1677677812
transform 1 0 4536 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7533
timestamp 1677677812
transform 1 0 4544 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_275
timestamp 1677677812
transform -1 0 4592 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7534
timestamp 1677677812
transform 1 0 4592 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7535
timestamp 1677677812
transform 1 0 4600 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7536
timestamp 1677677812
transform 1 0 4608 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7537
timestamp 1677677812
transform 1 0 4616 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7538
timestamp 1677677812
transform 1 0 4624 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7540
timestamp 1677677812
transform 1 0 4632 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_277
timestamp 1677677812
transform 1 0 4640 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7541
timestamp 1677677812
transform 1 0 4680 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7542
timestamp 1677677812
transform 1 0 4688 0 -1 1770
box -8 -3 16 105
use OAI22X1  OAI22X1_278
timestamp 1677677812
transform -1 0 4736 0 -1 1770
box -8 -3 46 105
use FILL  FILL_7543
timestamp 1677677812
transform 1 0 4736 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7544
timestamp 1677677812
transform 1 0 4744 0 -1 1770
box -8 -3 16 105
use INVX2  INVX2_479
timestamp 1677677812
transform -1 0 4768 0 -1 1770
box -9 -3 26 105
use FILL  FILL_7545
timestamp 1677677812
transform 1 0 4768 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7546
timestamp 1677677812
transform 1 0 4776 0 -1 1770
box -8 -3 16 105
use FILL  FILL_7547
timestamp 1677677812
transform 1 0 4784 0 -1 1770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_61
timestamp 1677677812
transform 1 0 4843 0 1 1670
box -10 -3 10 3
use M3_M2  M3_M2_5743
timestamp 1677677812
transform 1 0 132 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5716
timestamp 1677677812
transform 1 0 180 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5744
timestamp 1677677812
transform 1 0 180 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6381
timestamp 1677677812
transform 1 0 132 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6382
timestamp 1677677812
transform 1 0 164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6383
timestamp 1677677812
transform 1 0 172 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6384
timestamp 1677677812
transform 1 0 180 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6490
timestamp 1677677812
transform 1 0 84 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6491
timestamp 1677677812
transform 1 0 188 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5668
timestamp 1677677812
transform 1 0 220 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5669
timestamp 1677677812
transform 1 0 276 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5678
timestamp 1677677812
transform 1 0 204 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5679
timestamp 1677677812
transform 1 0 228 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5745
timestamp 1677677812
transform 1 0 268 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5746
timestamp 1677677812
transform 1 0 308 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6385
timestamp 1677677812
transform 1 0 204 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6386
timestamp 1677677812
transform 1 0 268 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6387
timestamp 1677677812
transform 1 0 300 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6388
timestamp 1677677812
transform 1 0 308 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5795
timestamp 1677677812
transform 1 0 204 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6492
timestamp 1677677812
transform 1 0 220 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5796
timestamp 1677677812
transform 1 0 244 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5814
timestamp 1677677812
transform 1 0 180 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5815
timestamp 1677677812
transform 1 0 196 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5816
timestamp 1677677812
transform 1 0 300 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5692
timestamp 1677677812
transform 1 0 332 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6389
timestamp 1677677812
transform 1 0 332 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5717
timestamp 1677677812
transform 1 0 388 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5747
timestamp 1677677812
transform 1 0 380 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5776
timestamp 1677677812
transform 1 0 356 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6390
timestamp 1677677812
transform 1 0 364 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6391
timestamp 1677677812
transform 1 0 380 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6493
timestamp 1677677812
transform 1 0 348 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6494
timestamp 1677677812
transform 1 0 356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6495
timestamp 1677677812
transform 1 0 372 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5817
timestamp 1677677812
transform 1 0 372 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5748
timestamp 1677677812
transform 1 0 420 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5777
timestamp 1677677812
transform 1 0 396 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5693
timestamp 1677677812
transform 1 0 540 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5749
timestamp 1677677812
transform 1 0 492 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5750
timestamp 1677677812
transform 1 0 532 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6392
timestamp 1677677812
transform 1 0 404 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6393
timestamp 1677677812
transform 1 0 428 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6394
timestamp 1677677812
transform 1 0 492 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6395
timestamp 1677677812
transform 1 0 524 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6396
timestamp 1677677812
transform 1 0 532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6397
timestamp 1677677812
transform 1 0 540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6496
timestamp 1677677812
transform 1 0 388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6497
timestamp 1677677812
transform 1 0 412 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6498
timestamp 1677677812
transform 1 0 428 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6499
timestamp 1677677812
transform 1 0 444 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5797
timestamp 1677677812
transform 1 0 524 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5818
timestamp 1677677812
transform 1 0 428 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5819
timestamp 1677677812
transform 1 0 460 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5820
timestamp 1677677812
transform 1 0 516 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5859
timestamp 1677677812
transform 1 0 404 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5860
timestamp 1677677812
transform 1 0 428 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5861
timestamp 1677677812
transform 1 0 476 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5751
timestamp 1677677812
transform 1 0 572 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5752
timestamp 1677677812
transform 1 0 588 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6398
timestamp 1677677812
transform 1 0 588 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6500
timestamp 1677677812
transform 1 0 572 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6501
timestamp 1677677812
transform 1 0 580 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5798
timestamp 1677677812
transform 1 0 588 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6502
timestamp 1677677812
transform 1 0 596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6503
timestamp 1677677812
transform 1 0 612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6399
timestamp 1677677812
transform 1 0 620 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5680
timestamp 1677677812
transform 1 0 684 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6400
timestamp 1677677812
transform 1 0 740 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5753
timestamp 1677677812
transform 1 0 764 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6401
timestamp 1677677812
transform 1 0 772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6504
timestamp 1677677812
transform 1 0 764 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5718
timestamp 1677677812
transform 1 0 788 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6402
timestamp 1677677812
transform 1 0 788 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5754
timestamp 1677677812
transform 1 0 828 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6403
timestamp 1677677812
transform 1 0 828 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6404
timestamp 1677677812
transform 1 0 844 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6405
timestamp 1677677812
transform 1 0 852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6505
timestamp 1677677812
transform 1 0 812 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6506
timestamp 1677677812
transform 1 0 820 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6507
timestamp 1677677812
transform 1 0 836 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5821
timestamp 1677677812
transform 1 0 812 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5862
timestamp 1677677812
transform 1 0 820 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5822
timestamp 1677677812
transform 1 0 860 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5778
timestamp 1677677812
transform 1 0 876 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5863
timestamp 1677677812
transform 1 0 868 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6508
timestamp 1677677812
transform 1 0 892 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5823
timestamp 1677677812
transform 1 0 892 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5719
timestamp 1677677812
transform 1 0 1020 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5755
timestamp 1677677812
transform 1 0 988 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5779
timestamp 1677677812
transform 1 0 940 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5756
timestamp 1677677812
transform 1 0 1028 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6406
timestamp 1677677812
transform 1 0 988 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6407
timestamp 1677677812
transform 1 0 1020 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6408
timestamp 1677677812
transform 1 0 1028 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6509
timestamp 1677677812
transform 1 0 940 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5824
timestamp 1677677812
transform 1 0 940 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5757
timestamp 1677677812
transform 1 0 1092 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6409
timestamp 1677677812
transform 1 0 1108 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5864
timestamp 1677677812
transform 1 0 1108 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5694
timestamp 1677677812
transform 1 0 1164 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5720
timestamp 1677677812
transform 1 0 1140 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5758
timestamp 1677677812
transform 1 0 1132 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6410
timestamp 1677677812
transform 1 0 1148 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5780
timestamp 1677677812
transform 1 0 1156 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6411
timestamp 1677677812
transform 1 0 1164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6510
timestamp 1677677812
transform 1 0 1132 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6511
timestamp 1677677812
transform 1 0 1140 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5825
timestamp 1677677812
transform 1 0 1156 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5865
timestamp 1677677812
transform 1 0 1204 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6363
timestamp 1677677812
transform 1 0 1220 0 1 1645
box -2 -2 2 2
use M2_M1  M2_M1_6512
timestamp 1677677812
transform 1 0 1220 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6364
timestamp 1677677812
transform 1 0 1244 0 1 1645
box -2 -2 2 2
use M3_M2  M3_M2_5721
timestamp 1677677812
transform 1 0 1244 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6513
timestamp 1677677812
transform 1 0 1244 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6412
timestamp 1677677812
transform 1 0 1260 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5799
timestamp 1677677812
transform 1 0 1260 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6514
timestamp 1677677812
transform 1 0 1268 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5800
timestamp 1677677812
transform 1 0 1284 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6413
timestamp 1677677812
transform 1 0 1324 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5781
timestamp 1677677812
transform 1 0 1332 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5801
timestamp 1677677812
transform 1 0 1324 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6515
timestamp 1677677812
transform 1 0 1332 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5695
timestamp 1677677812
transform 1 0 1380 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5722
timestamp 1677677812
transform 1 0 1356 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5759
timestamp 1677677812
transform 1 0 1348 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6414
timestamp 1677677812
transform 1 0 1348 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6415
timestamp 1677677812
transform 1 0 1356 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5782
timestamp 1677677812
transform 1 0 1364 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6416
timestamp 1677677812
transform 1 0 1372 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6516
timestamp 1677677812
transform 1 0 1356 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6517
timestamp 1677677812
transform 1 0 1364 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6518
timestamp 1677677812
transform 1 0 1380 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5723
timestamp 1677677812
transform 1 0 1396 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6417
timestamp 1677677812
transform 1 0 1420 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5826
timestamp 1677677812
transform 1 0 1420 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5696
timestamp 1677677812
transform 1 0 1452 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5760
timestamp 1677677812
transform 1 0 1476 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6418
timestamp 1677677812
transform 1 0 1436 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5783
timestamp 1677677812
transform 1 0 1444 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6419
timestamp 1677677812
transform 1 0 1476 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6519
timestamp 1677677812
transform 1 0 1516 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5827
timestamp 1677677812
transform 1 0 1444 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5828
timestamp 1677677812
transform 1 0 1484 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5829
timestamp 1677677812
transform 1 0 1516 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5830
timestamp 1677677812
transform 1 0 1532 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5761
timestamp 1677677812
transform 1 0 1580 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6520
timestamp 1677677812
transform 1 0 1580 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5831
timestamp 1677677812
transform 1 0 1572 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5724
timestamp 1677677812
transform 1 0 1636 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6420
timestamp 1677677812
transform 1 0 1636 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6421
timestamp 1677677812
transform 1 0 1644 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6422
timestamp 1677677812
transform 1 0 1660 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6521
timestamp 1677677812
transform 1 0 1636 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5802
timestamp 1677677812
transform 1 0 1644 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6522
timestamp 1677677812
transform 1 0 1652 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5803
timestamp 1677677812
transform 1 0 1660 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5866
timestamp 1677677812
transform 1 0 1644 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5670
timestamp 1677677812
transform 1 0 1676 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5697
timestamp 1677677812
transform 1 0 1676 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5698
timestamp 1677677812
transform 1 0 1692 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6423
timestamp 1677677812
transform 1 0 1676 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5762
timestamp 1677677812
transform 1 0 1700 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6424
timestamp 1677677812
transform 1 0 1700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6425
timestamp 1677677812
transform 1 0 1716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6523
timestamp 1677677812
transform 1 0 1684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6524
timestamp 1677677812
transform 1 0 1692 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6525
timestamp 1677677812
transform 1 0 1708 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5832
timestamp 1677677812
transform 1 0 1684 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5833
timestamp 1677677812
transform 1 0 1708 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5699
timestamp 1677677812
transform 1 0 1740 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5804
timestamp 1677677812
transform 1 0 1748 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5725
timestamp 1677677812
transform 1 0 1788 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6426
timestamp 1677677812
transform 1 0 1788 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6526
timestamp 1677677812
transform 1 0 1836 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5867
timestamp 1677677812
transform 1 0 1764 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6427
timestamp 1677677812
transform 1 0 1876 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5700
timestamp 1677677812
transform 1 0 1908 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6428
timestamp 1677677812
transform 1 0 1908 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5671
timestamp 1677677812
transform 1 0 1948 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6429
timestamp 1677677812
transform 1 0 1932 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6430
timestamp 1677677812
transform 1 0 1948 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6527
timestamp 1677677812
transform 1 0 1916 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6528
timestamp 1677677812
transform 1 0 1940 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5834
timestamp 1677677812
transform 1 0 1924 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6529
timestamp 1677677812
transform 1 0 1964 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6431
timestamp 1677677812
transform 1 0 1996 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5701
timestamp 1677677812
transform 1 0 2028 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5784
timestamp 1677677812
transform 1 0 2020 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6530
timestamp 1677677812
transform 1 0 2012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6531
timestamp 1677677812
transform 1 0 2020 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5672
timestamp 1677677812
transform 1 0 2044 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6432
timestamp 1677677812
transform 1 0 2092 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5681
timestamp 1677677812
transform 1 0 2116 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5682
timestamp 1677677812
transform 1 0 2148 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6532
timestamp 1677677812
transform 1 0 2148 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5835
timestamp 1677677812
transform 1 0 2148 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5868
timestamp 1677677812
transform 1 0 2156 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6433
timestamp 1677677812
transform 1 0 2252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6434
timestamp 1677677812
transform 1 0 2292 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6533
timestamp 1677677812
transform 1 0 2212 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6534
timestamp 1677677812
transform 1 0 2300 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6596
timestamp 1677677812
transform 1 0 2340 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5673
timestamp 1677677812
transform 1 0 2372 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6597
timestamp 1677677812
transform 1 0 2364 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5763
timestamp 1677677812
transform 1 0 2444 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6435
timestamp 1677677812
transform 1 0 2444 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6535
timestamp 1677677812
transform 1 0 2396 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6436
timestamp 1677677812
transform 1 0 2484 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5764
timestamp 1677677812
transform 1 0 2532 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6437
timestamp 1677677812
transform 1 0 2540 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6438
timestamp 1677677812
transform 1 0 2556 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6536
timestamp 1677677812
transform 1 0 2548 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5683
timestamp 1677677812
transform 1 0 2652 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5765
timestamp 1677677812
transform 1 0 2660 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5726
timestamp 1677677812
transform 1 0 2716 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5766
timestamp 1677677812
transform 1 0 2708 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6439
timestamp 1677677812
transform 1 0 2604 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6440
timestamp 1677677812
transform 1 0 2660 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6441
timestamp 1677677812
transform 1 0 2700 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6537
timestamp 1677677812
transform 1 0 2596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6538
timestamp 1677677812
transform 1 0 2684 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5869
timestamp 1677677812
transform 1 0 2652 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6442
timestamp 1677677812
transform 1 0 2716 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6539
timestamp 1677677812
transform 1 0 2708 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6540
timestamp 1677677812
transform 1 0 2716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6598
timestamp 1677677812
transform 1 0 2724 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5870
timestamp 1677677812
transform 1 0 2724 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6541
timestamp 1677677812
transform 1 0 2756 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6599
timestamp 1677677812
transform 1 0 2748 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5871
timestamp 1677677812
transform 1 0 2756 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5727
timestamp 1677677812
transform 1 0 2788 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6373
timestamp 1677677812
transform 1 0 2788 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6443
timestamp 1677677812
transform 1 0 2804 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6365
timestamp 1677677812
transform 1 0 2844 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6444
timestamp 1677677812
transform 1 0 2852 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6542
timestamp 1677677812
transform 1 0 2868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6543
timestamp 1677677812
transform 1 0 2884 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6544
timestamp 1677677812
transform 1 0 2908 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6374
timestamp 1677677812
transform 1 0 2924 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5728
timestamp 1677677812
transform 1 0 2940 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6445
timestamp 1677677812
transform 1 0 2940 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6366
timestamp 1677677812
transform 1 0 2956 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6446
timestamp 1677677812
transform 1 0 2956 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6447
timestamp 1677677812
transform 1 0 3012 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5836
timestamp 1677677812
transform 1 0 3012 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6600
timestamp 1677677812
transform 1 0 3020 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5872
timestamp 1677677812
transform 1 0 3020 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6448
timestamp 1677677812
transform 1 0 3036 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5729
timestamp 1677677812
transform 1 0 3060 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6375
timestamp 1677677812
transform 1 0 3052 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6545
timestamp 1677677812
transform 1 0 3060 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5702
timestamp 1677677812
transform 1 0 3100 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6367
timestamp 1677677812
transform 1 0 3076 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5730
timestamp 1677677812
transform 1 0 3092 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6376
timestamp 1677677812
transform 1 0 3092 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6449
timestamp 1677677812
transform 1 0 3084 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5837
timestamp 1677677812
transform 1 0 3068 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6601
timestamp 1677677812
transform 1 0 3100 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5873
timestamp 1677677812
transform 1 0 3100 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5731
timestamp 1677677812
transform 1 0 3116 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5703
timestamp 1677677812
transform 1 0 3132 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6368
timestamp 1677677812
transform 1 0 3124 0 1 1635
box -2 -2 2 2
use M2_M1  M2_M1_6450
timestamp 1677677812
transform 1 0 3116 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6377
timestamp 1677677812
transform 1 0 3132 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6546
timestamp 1677677812
transform 1 0 3124 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6369
timestamp 1677677812
transform 1 0 3172 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5767
timestamp 1677677812
transform 1 0 3172 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6378
timestamp 1677677812
transform 1 0 3180 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6451
timestamp 1677677812
transform 1 0 3164 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6452
timestamp 1677677812
transform 1 0 3196 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6547
timestamp 1677677812
transform 1 0 3204 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5674
timestamp 1677677812
transform 1 0 3220 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6370
timestamp 1677677812
transform 1 0 3220 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5768
timestamp 1677677812
transform 1 0 3220 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5874
timestamp 1677677812
transform 1 0 3220 0 1 1585
box -3 -3 3 3
use M2_M1  M2_M1_6379
timestamp 1677677812
transform 1 0 3228 0 1 1625
box -2 -2 2 2
use M2_M1  M2_M1_6489
timestamp 1677677812
transform 1 0 3236 0 1 1614
box -2 -2 2 2
use M2_M1  M2_M1_6380
timestamp 1677677812
transform 1 0 3268 0 1 1625
box -2 -2 2 2
use M3_M2  M3_M2_5875
timestamp 1677677812
transform 1 0 3252 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5785
timestamp 1677677812
transform 1 0 3276 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6548
timestamp 1677677812
transform 1 0 3276 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5838
timestamp 1677677812
transform 1 0 3276 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6453
timestamp 1677677812
transform 1 0 3292 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5769
timestamp 1677677812
transform 1 0 3332 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6602
timestamp 1677677812
transform 1 0 3340 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5770
timestamp 1677677812
transform 1 0 3388 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6454
timestamp 1677677812
transform 1 0 3388 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5805
timestamp 1677677812
transform 1 0 3428 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6455
timestamp 1677677812
transform 1 0 3452 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6549
timestamp 1677677812
transform 1 0 3444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6550
timestamp 1677677812
transform 1 0 3460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6603
timestamp 1677677812
transform 1 0 3428 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5839
timestamp 1677677812
transform 1 0 3452 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5806
timestamp 1677677812
transform 1 0 3476 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6604
timestamp 1677677812
transform 1 0 3484 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5675
timestamp 1677677812
transform 1 0 3516 0 1 1665
box -3 -3 3 3
use M2_M1  M2_M1_6456
timestamp 1677677812
transform 1 0 3508 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6551
timestamp 1677677812
transform 1 0 3500 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6552
timestamp 1677677812
transform 1 0 3524 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6605
timestamp 1677677812
transform 1 0 3508 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5876
timestamp 1677677812
transform 1 0 3524 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5732
timestamp 1677677812
transform 1 0 3540 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5771
timestamp 1677677812
transform 1 0 3548 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6457
timestamp 1677677812
transform 1 0 3548 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5684
timestamp 1677677812
transform 1 0 3628 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5733
timestamp 1677677812
transform 1 0 3604 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5772
timestamp 1677677812
transform 1 0 3660 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6458
timestamp 1677677812
transform 1 0 3652 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6459
timestamp 1677677812
transform 1 0 3660 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5807
timestamp 1677677812
transform 1 0 3556 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5734
timestamp 1677677812
transform 1 0 3708 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6460
timestamp 1677677812
transform 1 0 3676 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6461
timestamp 1677677812
transform 1 0 3708 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6553
timestamp 1677677812
transform 1 0 3668 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5840
timestamp 1677677812
transform 1 0 3556 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6606
timestamp 1677677812
transform 1 0 3564 0 1 1595
box -2 -2 2 2
use M3_M2  M3_M2_5841
timestamp 1677677812
transform 1 0 3588 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5877
timestamp 1677677812
transform 1 0 3572 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_5808
timestamp 1677677812
transform 1 0 3676 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5786
timestamp 1677677812
transform 1 0 3716 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6554
timestamp 1677677812
transform 1 0 3684 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6555
timestamp 1677677812
transform 1 0 3700 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6556
timestamp 1677677812
transform 1 0 3716 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6557
timestamp 1677677812
transform 1 0 3724 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5842
timestamp 1677677812
transform 1 0 3684 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5787
timestamp 1677677812
transform 1 0 3732 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_5843
timestamp 1677677812
transform 1 0 3724 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5676
timestamp 1677677812
transform 1 0 3764 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5677
timestamp 1677677812
transform 1 0 3796 0 1 1665
box -3 -3 3 3
use M3_M2  M3_M2_5685
timestamp 1677677812
transform 1 0 3788 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5704
timestamp 1677677812
transform 1 0 3772 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6462
timestamp 1677677812
transform 1 0 3772 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6463
timestamp 1677677812
transform 1 0 3788 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5788
timestamp 1677677812
transform 1 0 3796 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6558
timestamp 1677677812
transform 1 0 3780 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6559
timestamp 1677677812
transform 1 0 3796 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5705
timestamp 1677677812
transform 1 0 3900 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5735
timestamp 1677677812
transform 1 0 3876 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6464
timestamp 1677677812
transform 1 0 3876 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6465
timestamp 1677677812
transform 1 0 3892 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6466
timestamp 1677677812
transform 1 0 3900 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6560
timestamp 1677677812
transform 1 0 3868 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6561
timestamp 1677677812
transform 1 0 3884 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5809
timestamp 1677677812
transform 1 0 3892 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5844
timestamp 1677677812
transform 1 0 3868 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5686
timestamp 1677677812
transform 1 0 3964 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6467
timestamp 1677677812
transform 1 0 3964 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5706
timestamp 1677677812
transform 1 0 3980 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6468
timestamp 1677677812
transform 1 0 3980 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6562
timestamp 1677677812
transform 1 0 3940 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6563
timestamp 1677677812
transform 1 0 3956 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6564
timestamp 1677677812
transform 1 0 3972 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5845
timestamp 1677677812
transform 1 0 3932 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5846
timestamp 1677677812
transform 1 0 3972 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5687
timestamp 1677677812
transform 1 0 4036 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6469
timestamp 1677677812
transform 1 0 4036 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5789
timestamp 1677677812
transform 1 0 4044 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6565
timestamp 1677677812
transform 1 0 4012 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6566
timestamp 1677677812
transform 1 0 4028 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6567
timestamp 1677677812
transform 1 0 4044 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6568
timestamp 1677677812
transform 1 0 4052 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5847
timestamp 1677677812
transform 1 0 4012 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6470
timestamp 1677677812
transform 1 0 4060 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5810
timestamp 1677677812
transform 1 0 4060 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5736
timestamp 1677677812
transform 1 0 4092 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6471
timestamp 1677677812
transform 1 0 4092 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5790
timestamp 1677677812
transform 1 0 4100 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6569
timestamp 1677677812
transform 1 0 4068 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6570
timestamp 1677677812
transform 1 0 4084 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6571
timestamp 1677677812
transform 1 0 4100 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5848
timestamp 1677677812
transform 1 0 4052 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5849
timestamp 1677677812
transform 1 0 4076 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5850
timestamp 1677677812
transform 1 0 4092 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6472
timestamp 1677677812
transform 1 0 4116 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5811
timestamp 1677677812
transform 1 0 4116 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5773
timestamp 1677677812
transform 1 0 4132 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5737
timestamp 1677677812
transform 1 0 4164 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5791
timestamp 1677677812
transform 1 0 4140 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6473
timestamp 1677677812
transform 1 0 4164 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5707
timestamp 1677677812
transform 1 0 4188 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5792
timestamp 1677677812
transform 1 0 4180 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6474
timestamp 1677677812
transform 1 0 4188 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6572
timestamp 1677677812
transform 1 0 4140 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6573
timestamp 1677677812
transform 1 0 4156 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6574
timestamp 1677677812
transform 1 0 4172 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6575
timestamp 1677677812
transform 1 0 4180 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5851
timestamp 1677677812
transform 1 0 4172 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5688
timestamp 1677677812
transform 1 0 4236 0 1 1655
box -3 -3 3 3
use M2_M1  M2_M1_6475
timestamp 1677677812
transform 1 0 4236 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6476
timestamp 1677677812
transform 1 0 4252 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6576
timestamp 1677677812
transform 1 0 4228 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6577
timestamp 1677677812
transform 1 0 4244 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5812
timestamp 1677677812
transform 1 0 4252 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_5852
timestamp 1677677812
transform 1 0 4244 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5708
timestamp 1677677812
transform 1 0 4308 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5738
timestamp 1677677812
transform 1 0 4316 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6477
timestamp 1677677812
transform 1 0 4316 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6578
timestamp 1677677812
transform 1 0 4292 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6579
timestamp 1677677812
transform 1 0 4308 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5853
timestamp 1677677812
transform 1 0 4292 0 1 1595
box -3 -3 3 3
use M2_M1  M2_M1_6580
timestamp 1677677812
transform 1 0 4332 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5709
timestamp 1677677812
transform 1 0 4340 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6478
timestamp 1677677812
transform 1 0 4340 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6581
timestamp 1677677812
transform 1 0 4340 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5854
timestamp 1677677812
transform 1 0 4340 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5689
timestamp 1677677812
transform 1 0 4396 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5774
timestamp 1677677812
transform 1 0 4372 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6479
timestamp 1677677812
transform 1 0 4396 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6582
timestamp 1677677812
transform 1 0 4372 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6583
timestamp 1677677812
transform 1 0 4388 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6584
timestamp 1677677812
transform 1 0 4404 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5690
timestamp 1677677812
transform 1 0 4460 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5710
timestamp 1677677812
transform 1 0 4468 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5775
timestamp 1677677812
transform 1 0 4452 0 1 1625
box -3 -3 3 3
use M2_M1  M2_M1_6480
timestamp 1677677812
transform 1 0 4452 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6481
timestamp 1677677812
transform 1 0 4468 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6585
timestamp 1677677812
transform 1 0 4444 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6586
timestamp 1677677812
transform 1 0 4460 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6587
timestamp 1677677812
transform 1 0 4476 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6588
timestamp 1677677812
transform 1 0 4484 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5855
timestamp 1677677812
transform 1 0 4476 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5739
timestamp 1677677812
transform 1 0 4516 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6482
timestamp 1677677812
transform 1 0 4516 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6483
timestamp 1677677812
transform 1 0 4532 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6589
timestamp 1677677812
transform 1 0 4524 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5813
timestamp 1677677812
transform 1 0 4532 0 1 1605
box -3 -3 3 3
use M2_M1  M2_M1_6590
timestamp 1677677812
transform 1 0 4540 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5856
timestamp 1677677812
transform 1 0 4540 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5691
timestamp 1677677812
transform 1 0 4564 0 1 1655
box -3 -3 3 3
use M3_M2  M3_M2_5711
timestamp 1677677812
transform 1 0 4556 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6371
timestamp 1677677812
transform 1 0 4564 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5712
timestamp 1677677812
transform 1 0 4580 0 1 1645
box -3 -3 3 3
use M2_M1  M2_M1_6372
timestamp 1677677812
transform 1 0 4580 0 1 1635
box -2 -2 2 2
use M3_M2  M3_M2_5740
timestamp 1677677812
transform 1 0 4620 0 1 1635
box -3 -3 3 3
use M2_M1  M2_M1_6484
timestamp 1677677812
transform 1 0 4604 0 1 1615
box -2 -2 2 2
use M3_M2  M3_M2_5793
timestamp 1677677812
transform 1 0 4612 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6485
timestamp 1677677812
transform 1 0 4620 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6591
timestamp 1677677812
transform 1 0 4596 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6592
timestamp 1677677812
transform 1 0 4612 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6593
timestamp 1677677812
transform 1 0 4628 0 1 1605
box -2 -2 2 2
use M3_M2  M3_M2_5857
timestamp 1677677812
transform 1 0 4596 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5858
timestamp 1677677812
transform 1 0 4636 0 1 1595
box -3 -3 3 3
use M3_M2  M3_M2_5713
timestamp 1677677812
transform 1 0 4684 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5714
timestamp 1677677812
transform 1 0 4732 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5715
timestamp 1677677812
transform 1 0 4756 0 1 1645
box -3 -3 3 3
use M3_M2  M3_M2_5741
timestamp 1677677812
transform 1 0 4660 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5742
timestamp 1677677812
transform 1 0 4692 0 1 1635
box -3 -3 3 3
use M3_M2  M3_M2_5794
timestamp 1677677812
transform 1 0 4668 0 1 1615
box -3 -3 3 3
use M2_M1  M2_M1_6486
timestamp 1677677812
transform 1 0 4692 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6487
timestamp 1677677812
transform 1 0 4748 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6488
timestamp 1677677812
transform 1 0 4756 0 1 1615
box -2 -2 2 2
use M2_M1  M2_M1_6594
timestamp 1677677812
transform 1 0 4668 0 1 1605
box -2 -2 2 2
use M2_M1  M2_M1_6595
timestamp 1677677812
transform 1 0 4764 0 1 1605
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_62
timestamp 1677677812
transform 1 0 48 0 1 1570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_409
timestamp 1677677812
transform 1 0 72 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_480
timestamp 1677677812
transform -1 0 184 0 1 1570
box -9 -3 26 105
use FILL  FILL_7548
timestamp 1677677812
transform 1 0 184 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_481
timestamp 1677677812
transform -1 0 208 0 1 1570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_410
timestamp 1677677812
transform 1 0 208 0 1 1570
box -8 -3 104 105
use FILL  FILL_7549
timestamp 1677677812
transform 1 0 304 0 1 1570
box -8 -3 16 105
use FILL  FILL_7550
timestamp 1677677812
transform 1 0 312 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_482
timestamp 1677677812
transform -1 0 336 0 1 1570
box -9 -3 26 105
use FILL  FILL_7551
timestamp 1677677812
transform 1 0 336 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_284
timestamp 1677677812
transform 1 0 344 0 1 1570
box -8 -3 46 105
use FILL  FILL_7555
timestamp 1677677812
transform 1 0 384 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_279
timestamp 1677677812
transform -1 0 432 0 1 1570
box -8 -3 46 105
use M3_M2  M3_M2_5878
timestamp 1677677812
transform 1 0 444 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_5879
timestamp 1677677812
transform 1 0 476 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_413
timestamp 1677677812
transform 1 0 432 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_484
timestamp 1677677812
transform -1 0 544 0 1 1570
box -9 -3 26 105
use FILL  FILL_7556
timestamp 1677677812
transform 1 0 544 0 1 1570
box -8 -3 16 105
use FILL  FILL_7557
timestamp 1677677812
transform 1 0 552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7558
timestamp 1677677812
transform 1 0 560 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_286
timestamp 1677677812
transform 1 0 568 0 1 1570
box -8 -3 46 105
use FILL  FILL_7565
timestamp 1677677812
transform 1 0 608 0 1 1570
box -8 -3 16 105
use FILL  FILL_7566
timestamp 1677677812
transform 1 0 616 0 1 1570
box -8 -3 16 105
use FILL  FILL_7567
timestamp 1677677812
transform 1 0 624 0 1 1570
box -8 -3 16 105
use FILL  FILL_7571
timestamp 1677677812
transform 1 0 632 0 1 1570
box -8 -3 16 105
use FILL  FILL_7573
timestamp 1677677812
transform 1 0 640 0 1 1570
box -8 -3 16 105
use FILL  FILL_7575
timestamp 1677677812
transform 1 0 648 0 1 1570
box -8 -3 16 105
use FILL  FILL_7577
timestamp 1677677812
transform 1 0 656 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5880
timestamp 1677677812
transform 1 0 676 0 1 1575
box -3 -3 3 3
use FILL  FILL_7578
timestamp 1677677812
transform 1 0 664 0 1 1570
box -8 -3 16 105
use FILL  FILL_7579
timestamp 1677677812
transform 1 0 672 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5881
timestamp 1677677812
transform 1 0 692 0 1 1575
box -3 -3 3 3
use FILL  FILL_7580
timestamp 1677677812
transform 1 0 680 0 1 1570
box -8 -3 16 105
use FILL  FILL_7581
timestamp 1677677812
transform 1 0 688 0 1 1570
box -8 -3 16 105
use FILL  FILL_7582
timestamp 1677677812
transform 1 0 696 0 1 1570
box -8 -3 16 105
use FILL  FILL_7584
timestamp 1677677812
transform 1 0 704 0 1 1570
box -8 -3 16 105
use FILL  FILL_7586
timestamp 1677677812
transform 1 0 712 0 1 1570
box -8 -3 16 105
use FILL  FILL_7587
timestamp 1677677812
transform 1 0 720 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_485
timestamp 1677677812
transform -1 0 744 0 1 1570
box -9 -3 26 105
use FILL  FILL_7588
timestamp 1677677812
transform 1 0 744 0 1 1570
box -8 -3 16 105
use FILL  FILL_7589
timestamp 1677677812
transform 1 0 752 0 1 1570
box -8 -3 16 105
use FILL  FILL_7590
timestamp 1677677812
transform 1 0 760 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_486
timestamp 1677677812
transform -1 0 784 0 1 1570
box -9 -3 26 105
use FILL  FILL_7591
timestamp 1677677812
transform 1 0 784 0 1 1570
box -8 -3 16 105
use FILL  FILL_7592
timestamp 1677677812
transform 1 0 792 0 1 1570
box -8 -3 16 105
use FILL  FILL_7593
timestamp 1677677812
transform 1 0 800 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_288
timestamp 1677677812
transform 1 0 808 0 1 1570
box -8 -3 46 105
use FILL  FILL_7594
timestamp 1677677812
transform 1 0 848 0 1 1570
box -8 -3 16 105
use FILL  FILL_7595
timestamp 1677677812
transform 1 0 856 0 1 1570
box -8 -3 16 105
use FILL  FILL_7596
timestamp 1677677812
transform 1 0 864 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_93
timestamp 1677677812
transform 1 0 872 0 1 1570
box -5 -3 28 105
use FILL  FILL_7597
timestamp 1677677812
transform 1 0 896 0 1 1570
box -8 -3 16 105
use FILL  FILL_7605
timestamp 1677677812
transform 1 0 904 0 1 1570
box -8 -3 16 105
use FILL  FILL_7607
timestamp 1677677812
transform 1 0 912 0 1 1570
box -8 -3 16 105
use FILL  FILL_7608
timestamp 1677677812
transform 1 0 920 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_416
timestamp 1677677812
transform 1 0 928 0 1 1570
box -8 -3 104 105
use FILL  FILL_7609
timestamp 1677677812
transform 1 0 1024 0 1 1570
box -8 -3 16 105
use FILL  FILL_7619
timestamp 1677677812
transform 1 0 1032 0 1 1570
box -8 -3 16 105
use FILL  FILL_7621
timestamp 1677677812
transform 1 0 1040 0 1 1570
box -8 -3 16 105
use FILL  FILL_7623
timestamp 1677677812
transform 1 0 1048 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_487
timestamp 1677677812
transform -1 0 1072 0 1 1570
box -9 -3 26 105
use FILL  FILL_7624
timestamp 1677677812
transform 1 0 1072 0 1 1570
box -8 -3 16 105
use FILL  FILL_7629
timestamp 1677677812
transform 1 0 1080 0 1 1570
box -8 -3 16 105
use FILL  FILL_7630
timestamp 1677677812
transform 1 0 1088 0 1 1570
box -8 -3 16 105
use FILL  FILL_7631
timestamp 1677677812
transform 1 0 1096 0 1 1570
box -8 -3 16 105
use FILL  FILL_7632
timestamp 1677677812
transform 1 0 1104 0 1 1570
box -8 -3 16 105
use FILL  FILL_7633
timestamp 1677677812
transform 1 0 1112 0 1 1570
box -8 -3 16 105
use FILL  FILL_7634
timestamp 1677677812
transform 1 0 1120 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_290
timestamp 1677677812
transform -1 0 1168 0 1 1570
box -8 -3 46 105
use FILL  FILL_7635
timestamp 1677677812
transform 1 0 1168 0 1 1570
box -8 -3 16 105
use FILL  FILL_7636
timestamp 1677677812
transform 1 0 1176 0 1 1570
box -8 -3 16 105
use FILL  FILL_7638
timestamp 1677677812
transform 1 0 1184 0 1 1570
box -8 -3 16 105
use FILL  FILL_7640
timestamp 1677677812
transform 1 0 1192 0 1 1570
box -8 -3 16 105
use FILL  FILL_7642
timestamp 1677677812
transform 1 0 1200 0 1 1570
box -8 -3 16 105
use FILL  FILL_7644
timestamp 1677677812
transform 1 0 1208 0 1 1570
box -8 -3 16 105
use FILL  FILL_7646
timestamp 1677677812
transform 1 0 1216 0 1 1570
box -8 -3 16 105
use FILL  FILL_7647
timestamp 1677677812
transform 1 0 1224 0 1 1570
box -8 -3 16 105
use FILL  FILL_7648
timestamp 1677677812
transform 1 0 1232 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5882
timestamp 1677677812
transform 1 0 1252 0 1 1575
box -3 -3 3 3
use FILL  FILL_7649
timestamp 1677677812
transform 1 0 1240 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_282
timestamp 1677677812
transform -1 0 1288 0 1 1570
box -8 -3 46 105
use FILL  FILL_7650
timestamp 1677677812
transform 1 0 1288 0 1 1570
box -8 -3 16 105
use FILL  FILL_7656
timestamp 1677677812
transform 1 0 1296 0 1 1570
box -8 -3 16 105
use FILL  FILL_7657
timestamp 1677677812
transform 1 0 1304 0 1 1570
box -8 -3 16 105
use FILL  FILL_7658
timestamp 1677677812
transform 1 0 1312 0 1 1570
box -8 -3 16 105
use FILL  FILL_7659
timestamp 1677677812
transform 1 0 1320 0 1 1570
box -8 -3 16 105
use FILL  FILL_7660
timestamp 1677677812
transform 1 0 1328 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5883
timestamp 1677677812
transform 1 0 1356 0 1 1575
box -3 -3 3 3
use INVX2  INVX2_488
timestamp 1677677812
transform -1 0 1352 0 1 1570
box -9 -3 26 105
use AOI22X1  AOI22X1_292
timestamp 1677677812
transform -1 0 1392 0 1 1570
box -8 -3 46 105
use FILL  FILL_7661
timestamp 1677677812
transform 1 0 1392 0 1 1570
box -8 -3 16 105
use FILL  FILL_7662
timestamp 1677677812
transform 1 0 1400 0 1 1570
box -8 -3 16 105
use FILL  FILL_7663
timestamp 1677677812
transform 1 0 1408 0 1 1570
box -8 -3 16 105
use FILL  FILL_7664
timestamp 1677677812
transform 1 0 1416 0 1 1570
box -8 -3 16 105
use FILL  FILL_7665
timestamp 1677677812
transform 1 0 1424 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_418
timestamp 1677677812
transform -1 0 1528 0 1 1570
box -8 -3 104 105
use FILL  FILL_7666
timestamp 1677677812
transform 1 0 1528 0 1 1570
box -8 -3 16 105
use FILL  FILL_7667
timestamp 1677677812
transform 1 0 1536 0 1 1570
box -8 -3 16 105
use FILL  FILL_7668
timestamp 1677677812
transform 1 0 1544 0 1 1570
box -8 -3 16 105
use FILL  FILL_7669
timestamp 1677677812
transform 1 0 1552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7670
timestamp 1677677812
transform 1 0 1560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7671
timestamp 1677677812
transform 1 0 1568 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_489
timestamp 1677677812
transform 1 0 1576 0 1 1570
box -9 -3 26 105
use FILL  FILL_7672
timestamp 1677677812
transform 1 0 1592 0 1 1570
box -8 -3 16 105
use FILL  FILL_7687
timestamp 1677677812
transform 1 0 1600 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5884
timestamp 1677677812
transform 1 0 1620 0 1 1575
box -3 -3 3 3
use FILL  FILL_7689
timestamp 1677677812
transform 1 0 1608 0 1 1570
box -8 -3 16 105
use FILL  FILL_7690
timestamp 1677677812
transform 1 0 1616 0 1 1570
box -8 -3 16 105
use FILL  FILL_7691
timestamp 1677677812
transform 1 0 1624 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_284
timestamp 1677677812
transform 1 0 1632 0 1 1570
box -8 -3 46 105
use M3_M2  M3_M2_5885
timestamp 1677677812
transform 1 0 1684 0 1 1575
box -3 -3 3 3
use FILL  FILL_7692
timestamp 1677677812
transform 1 0 1672 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_294
timestamp 1677677812
transform 1 0 1680 0 1 1570
box -8 -3 46 105
use FILL  FILL_7693
timestamp 1677677812
transform 1 0 1720 0 1 1570
box -8 -3 16 105
use FILL  FILL_7697
timestamp 1677677812
transform 1 0 1728 0 1 1570
box -8 -3 16 105
use FILL  FILL_7698
timestamp 1677677812
transform 1 0 1736 0 1 1570
box -8 -3 16 105
use FILL  FILL_7699
timestamp 1677677812
transform 1 0 1744 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5886
timestamp 1677677812
transform 1 0 1836 0 1 1575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_421
timestamp 1677677812
transform -1 0 1848 0 1 1570
box -8 -3 104 105
use FILL  FILL_7700
timestamp 1677677812
transform 1 0 1848 0 1 1570
box -8 -3 16 105
use FILL  FILL_7701
timestamp 1677677812
transform 1 0 1856 0 1 1570
box -8 -3 16 105
use FILL  FILL_7702
timestamp 1677677812
transform 1 0 1864 0 1 1570
box -8 -3 16 105
use FILL  FILL_7703
timestamp 1677677812
transform 1 0 1872 0 1 1570
box -8 -3 16 105
use FILL  FILL_7704
timestamp 1677677812
transform 1 0 1880 0 1 1570
box -8 -3 16 105
use FILL  FILL_7705
timestamp 1677677812
transform 1 0 1888 0 1 1570
box -8 -3 16 105
use FILL  FILL_7706
timestamp 1677677812
transform 1 0 1896 0 1 1570
box -8 -3 16 105
use FILL  FILL_7707
timestamp 1677677812
transform 1 0 1904 0 1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_295
timestamp 1677677812
transform -1 0 1952 0 1 1570
box -8 -3 46 105
use FILL  FILL_7708
timestamp 1677677812
transform 1 0 1952 0 1 1570
box -8 -3 16 105
use FILL  FILL_7709
timestamp 1677677812
transform 1 0 1960 0 1 1570
box -8 -3 16 105
use FILL  FILL_7721
timestamp 1677677812
transform 1 0 1968 0 1 1570
box -8 -3 16 105
use AND2X2  AND2X2_49
timestamp 1677677812
transform -1 0 2008 0 1 1570
box -8 -3 40 105
use FILL  FILL_7722
timestamp 1677677812
transform 1 0 2008 0 1 1570
box -8 -3 16 105
use FILL  FILL_7726
timestamp 1677677812
transform 1 0 2016 0 1 1570
box -8 -3 16 105
use FILL  FILL_7728
timestamp 1677677812
transform 1 0 2024 0 1 1570
box -8 -3 16 105
use FILL  FILL_7730
timestamp 1677677812
transform 1 0 2032 0 1 1570
box -8 -3 16 105
use FILL  FILL_7731
timestamp 1677677812
transform 1 0 2040 0 1 1570
box -8 -3 16 105
use FILL  FILL_7732
timestamp 1677677812
transform 1 0 2048 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_95
timestamp 1677677812
transform -1 0 2080 0 1 1570
box -5 -3 28 105
use FILL  FILL_7733
timestamp 1677677812
transform 1 0 2080 0 1 1570
box -8 -3 16 105
use FILL  FILL_7734
timestamp 1677677812
transform 1 0 2088 0 1 1570
box -8 -3 16 105
use FILL  FILL_7735
timestamp 1677677812
transform 1 0 2096 0 1 1570
box -8 -3 16 105
use FILL  FILL_7736
timestamp 1677677812
transform 1 0 2104 0 1 1570
box -8 -3 16 105
use FILL  FILL_7737
timestamp 1677677812
transform 1 0 2112 0 1 1570
box -8 -3 16 105
use FILL  FILL_7738
timestamp 1677677812
transform 1 0 2120 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_96
timestamp 1677677812
transform 1 0 2128 0 1 1570
box -5 -3 28 105
use FILL  FILL_7739
timestamp 1677677812
transform 1 0 2152 0 1 1570
box -8 -3 16 105
use FILL  FILL_7740
timestamp 1677677812
transform 1 0 2160 0 1 1570
box -8 -3 16 105
use FILL  FILL_7743
timestamp 1677677812
transform 1 0 2168 0 1 1570
box -8 -3 16 105
use FILL  FILL_7745
timestamp 1677677812
transform 1 0 2176 0 1 1570
box -8 -3 16 105
use FILL  FILL_7747
timestamp 1677677812
transform 1 0 2184 0 1 1570
box -8 -3 16 105
use FILL  FILL_7749
timestamp 1677677812
transform 1 0 2192 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_424
timestamp 1677677812
transform 1 0 2200 0 1 1570
box -8 -3 104 105
use FILL  FILL_7750
timestamp 1677677812
transform 1 0 2296 0 1 1570
box -8 -3 16 105
use FILL  FILL_7761
timestamp 1677677812
transform 1 0 2304 0 1 1570
box -8 -3 16 105
use FILL  FILL_7763
timestamp 1677677812
transform 1 0 2312 0 1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_76
timestamp 1677677812
transform -1 0 2344 0 1 1570
box -8 -3 32 105
use FILL  FILL_7764
timestamp 1677677812
transform 1 0 2344 0 1 1570
box -8 -3 16 105
use FILL  FILL_7765
timestamp 1677677812
transform 1 0 2352 0 1 1570
box -8 -3 16 105
use FILL  FILL_7766
timestamp 1677677812
transform 1 0 2360 0 1 1570
box -8 -3 16 105
use FILL  FILL_7767
timestamp 1677677812
transform 1 0 2368 0 1 1570
box -8 -3 16 105
use FILL  FILL_7768
timestamp 1677677812
transform 1 0 2376 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_425
timestamp 1677677812
transform 1 0 2384 0 1 1570
box -8 -3 104 105
use FILL  FILL_7769
timestamp 1677677812
transform 1 0 2480 0 1 1570
box -8 -3 16 105
use FILL  FILL_7770
timestamp 1677677812
transform 1 0 2488 0 1 1570
box -8 -3 16 105
use FILL  FILL_7771
timestamp 1677677812
transform 1 0 2496 0 1 1570
box -8 -3 16 105
use FILL  FILL_7772
timestamp 1677677812
transform 1 0 2504 0 1 1570
box -8 -3 16 105
use FILL  FILL_7773
timestamp 1677677812
transform 1 0 2512 0 1 1570
box -8 -3 16 105
use FILL  FILL_7774
timestamp 1677677812
transform 1 0 2520 0 1 1570
box -8 -3 16 105
use FILL  FILL_7775
timestamp 1677677812
transform 1 0 2528 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_492
timestamp 1677677812
transform -1 0 2552 0 1 1570
box -9 -3 26 105
use FILL  FILL_7776
timestamp 1677677812
transform 1 0 2552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7777
timestamp 1677677812
transform 1 0 2560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7778
timestamp 1677677812
transform 1 0 2568 0 1 1570
box -8 -3 16 105
use BUFX2  BUFX2_98
timestamp 1677677812
transform 1 0 2576 0 1 1570
box -5 -3 28 105
use DFFNEGX1  DFFNEGX1_426
timestamp 1677677812
transform -1 0 2696 0 1 1570
box -8 -3 104 105
use NOR2X1  NOR2X1_77
timestamp 1677677812
transform -1 0 2720 0 1 1570
box -8 -3 32 105
use NOR2X1  NOR2X1_78
timestamp 1677677812
transform -1 0 2744 0 1 1570
box -8 -3 32 105
use FILL  FILL_7779
timestamp 1677677812
transform 1 0 2744 0 1 1570
box -8 -3 16 105
use FILL  FILL_7780
timestamp 1677677812
transform 1 0 2752 0 1 1570
box -8 -3 16 105
use FILL  FILL_7781
timestamp 1677677812
transform 1 0 2760 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_493
timestamp 1677677812
transform 1 0 2768 0 1 1570
box -9 -3 26 105
use NAND3X1  NAND3X1_56
timestamp 1677677812
transform -1 0 2816 0 1 1570
box -8 -3 40 105
use FILL  FILL_7782
timestamp 1677677812
transform 1 0 2816 0 1 1570
box -8 -3 16 105
use FILL  FILL_7811
timestamp 1677677812
transform 1 0 2824 0 1 1570
box -8 -3 16 105
use FILL  FILL_7813
timestamp 1677677812
transform 1 0 2832 0 1 1570
box -8 -3 16 105
use FILL  FILL_7814
timestamp 1677677812
transform 1 0 2840 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_494
timestamp 1677677812
transform -1 0 2864 0 1 1570
box -9 -3 26 105
use FILL  FILL_7815
timestamp 1677677812
transform 1 0 2864 0 1 1570
box -8 -3 16 105
use FILL  FILL_7817
timestamp 1677677812
transform 1 0 2872 0 1 1570
box -8 -3 16 105
use FILL  FILL_7819
timestamp 1677677812
transform 1 0 2880 0 1 1570
box -8 -3 16 105
use FILL  FILL_7821
timestamp 1677677812
transform 1 0 2888 0 1 1570
box -8 -3 16 105
use FILL  FILL_7822
timestamp 1677677812
transform 1 0 2896 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_495
timestamp 1677677812
transform 1 0 2904 0 1 1570
box -9 -3 26 105
use FILL  FILL_7823
timestamp 1677677812
transform 1 0 2920 0 1 1570
box -8 -3 16 105
use FILL  FILL_7824
timestamp 1677677812
transform 1 0 2928 0 1 1570
box -8 -3 16 105
use FILL  FILL_7825
timestamp 1677677812
transform 1 0 2936 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_58
timestamp 1677677812
transform 1 0 2944 0 1 1570
box -8 -3 40 105
use FILL  FILL_7826
timestamp 1677677812
transform 1 0 2976 0 1 1570
box -8 -3 16 105
use FILL  FILL_7827
timestamp 1677677812
transform 1 0 2984 0 1 1570
box -8 -3 16 105
use FILL  FILL_7828
timestamp 1677677812
transform 1 0 2992 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_496
timestamp 1677677812
transform 1 0 3000 0 1 1570
box -9 -3 26 105
use NOR2X1  NOR2X1_79
timestamp 1677677812
transform 1 0 3016 0 1 1570
box -8 -3 32 105
use FILL  FILL_7829
timestamp 1677677812
transform 1 0 3040 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5887
timestamp 1677677812
transform 1 0 3060 0 1 1575
box -3 -3 3 3
use FILL  FILL_7830
timestamp 1677677812
transform 1 0 3048 0 1 1570
box -8 -3 16 105
use FILL  FILL_7831
timestamp 1677677812
transform 1 0 3056 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_59
timestamp 1677677812
transform -1 0 3096 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_5888
timestamp 1677677812
transform 1 0 3108 0 1 1575
box -3 -3 3 3
use NOR2X1  NOR2X1_80
timestamp 1677677812
transform 1 0 3096 0 1 1570
box -8 -3 32 105
use FILL  FILL_7832
timestamp 1677677812
transform 1 0 3120 0 1 1570
box -8 -3 16 105
use FILL  FILL_7833
timestamp 1677677812
transform 1 0 3128 0 1 1570
box -8 -3 16 105
use FILL  FILL_7834
timestamp 1677677812
transform 1 0 3136 0 1 1570
box -8 -3 16 105
use FILL  FILL_7840
timestamp 1677677812
transform 1 0 3144 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_60
timestamp 1677677812
transform 1 0 3152 0 1 1570
box -8 -3 40 105
use M3_M2  M3_M2_5889
timestamp 1677677812
transform 1 0 3196 0 1 1575
box -3 -3 3 3
use FILL  FILL_7841
timestamp 1677677812
transform 1 0 3184 0 1 1570
box -8 -3 16 105
use FILL  FILL_7844
timestamp 1677677812
transform 1 0 3192 0 1 1570
box -8 -3 16 105
use INVX2  INVX2_499
timestamp 1677677812
transform 1 0 3200 0 1 1570
box -9 -3 26 105
use FILL  FILL_7845
timestamp 1677677812
transform 1 0 3216 0 1 1570
box -8 -3 16 105
use FILL  FILL_7846
timestamp 1677677812
transform 1 0 3224 0 1 1570
box -8 -3 16 105
use FILL  FILL_7847
timestamp 1677677812
transform 1 0 3232 0 1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_61
timestamp 1677677812
transform 1 0 3240 0 1 1570
box -8 -3 40 105
use FILL  FILL_7848
timestamp 1677677812
transform 1 0 3272 0 1 1570
box -8 -3 16 105
use FILL  FILL_7849
timestamp 1677677812
transform 1 0 3280 0 1 1570
box -8 -3 16 105
use FILL  FILL_7850
timestamp 1677677812
transform 1 0 3288 0 1 1570
box -8 -3 16 105
use FILL  FILL_7851
timestamp 1677677812
transform 1 0 3296 0 1 1570
box -8 -3 16 105
use FILL  FILL_7852
timestamp 1677677812
transform 1 0 3304 0 1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1677677812
transform 1 0 3312 0 1 1570
box -7 -3 39 105
use FILL  FILL_7853
timestamp 1677677812
transform 1 0 3344 0 1 1570
box -8 -3 16 105
use FILL  FILL_7854
timestamp 1677677812
transform 1 0 3352 0 1 1570
box -8 -3 16 105
use FILL  FILL_7855
timestamp 1677677812
transform 1 0 3360 0 1 1570
box -8 -3 16 105
use FILL  FILL_7856
timestamp 1677677812
transform 1 0 3368 0 1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_6
timestamp 1677677812
transform 1 0 3376 0 1 1570
box -8 -3 32 105
use FILL  FILL_7860
timestamp 1677677812
transform 1 0 3400 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5890
timestamp 1677677812
transform 1 0 3420 0 1 1575
box -3 -3 3 3
use FILL  FILL_7861
timestamp 1677677812
transform 1 0 3408 0 1 1570
box -8 -3 16 105
use FILL  FILL_7862
timestamp 1677677812
transform 1 0 3416 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5891
timestamp 1677677812
transform 1 0 3444 0 1 1575
box -3 -3 3 3
use AOI21X1  AOI21X1_1
timestamp 1677677812
transform -1 0 3456 0 1 1570
box -7 -3 39 105
use INVX2  INVX2_501
timestamp 1677677812
transform 1 0 3456 0 1 1570
box -9 -3 26 105
use FILL  FILL_7863
timestamp 1677677812
transform 1 0 3472 0 1 1570
box -8 -3 16 105
use FILL  FILL_7864
timestamp 1677677812
transform 1 0 3480 0 1 1570
box -8 -3 16 105
use FILL  FILL_7865
timestamp 1677677812
transform 1 0 3488 0 1 1570
box -8 -3 16 105
use FILL  FILL_7866
timestamp 1677677812
transform 1 0 3496 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5892
timestamp 1677677812
transform 1 0 3532 0 1 1575
box -3 -3 3 3
use AOI21X1  AOI21X1_2
timestamp 1677677812
transform -1 0 3536 0 1 1570
box -7 -3 39 105
use FILL  FILL_7867
timestamp 1677677812
transform 1 0 3536 0 1 1570
box -8 -3 16 105
use FILL  FILL_7880
timestamp 1677677812
transform 1 0 3544 0 1 1570
box -8 -3 16 105
use M3_M2  M3_M2_5893
timestamp 1677677812
transform 1 0 3612 0 1 1575
box -3 -3 3 3
use FAX1  FAX1_3
timestamp 1677677812
transform -1 0 3672 0 1 1570
box -5 -3 126 105
use FILL  FILL_7881
timestamp 1677677812
transform 1 0 3672 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_287
timestamp 1677677812
transform 1 0 3680 0 1 1570
box -8 -3 46 105
use FILL  FILL_7882
timestamp 1677677812
transform 1 0 3720 0 1 1570
box -8 -3 16 105
use FILL  FILL_7883
timestamp 1677677812
transform 1 0 3728 0 1 1570
box -8 -3 16 105
use FILL  FILL_7884
timestamp 1677677812
transform 1 0 3736 0 1 1570
box -8 -3 16 105
use FILL  FILL_7885
timestamp 1677677812
transform 1 0 3744 0 1 1570
box -8 -3 16 105
use FILL  FILL_7896
timestamp 1677677812
transform 1 0 3752 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_288
timestamp 1677677812
transform 1 0 3760 0 1 1570
box -8 -3 46 105
use FILL  FILL_7898
timestamp 1677677812
transform 1 0 3800 0 1 1570
box -8 -3 16 105
use FILL  FILL_7899
timestamp 1677677812
transform 1 0 3808 0 1 1570
box -8 -3 16 105
use FILL  FILL_7900
timestamp 1677677812
transform 1 0 3816 0 1 1570
box -8 -3 16 105
use FILL  FILL_7901
timestamp 1677677812
transform 1 0 3824 0 1 1570
box -8 -3 16 105
use FILL  FILL_7902
timestamp 1677677812
transform 1 0 3832 0 1 1570
box -8 -3 16 105
use FILL  FILL_7903
timestamp 1677677812
transform 1 0 3840 0 1 1570
box -8 -3 16 105
use FILL  FILL_7904
timestamp 1677677812
transform 1 0 3848 0 1 1570
box -8 -3 16 105
use FILL  FILL_7905
timestamp 1677677812
transform 1 0 3856 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_289
timestamp 1677677812
transform -1 0 3904 0 1 1570
box -8 -3 46 105
use FILL  FILL_7906
timestamp 1677677812
transform 1 0 3904 0 1 1570
box -8 -3 16 105
use FILL  FILL_7916
timestamp 1677677812
transform 1 0 3912 0 1 1570
box -8 -3 16 105
use FILL  FILL_7918
timestamp 1677677812
transform 1 0 3920 0 1 1570
box -8 -3 16 105
use FILL  FILL_7920
timestamp 1677677812
transform 1 0 3928 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_290
timestamp 1677677812
transform 1 0 3936 0 1 1570
box -8 -3 46 105
use FILL  FILL_7921
timestamp 1677677812
transform 1 0 3976 0 1 1570
box -8 -3 16 105
use FILL  FILL_7926
timestamp 1677677812
transform 1 0 3984 0 1 1570
box -8 -3 16 105
use FILL  FILL_7928
timestamp 1677677812
transform 1 0 3992 0 1 1570
box -8 -3 16 105
use FILL  FILL_7930
timestamp 1677677812
transform 1 0 4000 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_291
timestamp 1677677812
transform 1 0 4008 0 1 1570
box -8 -3 46 105
use FILL  FILL_7932
timestamp 1677677812
transform 1 0 4048 0 1 1570
box -8 -3 16 105
use FILL  FILL_7933
timestamp 1677677812
transform 1 0 4056 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_292
timestamp 1677677812
transform 1 0 4064 0 1 1570
box -8 -3 46 105
use FILL  FILL_7934
timestamp 1677677812
transform 1 0 4104 0 1 1570
box -8 -3 16 105
use FILL  FILL_7935
timestamp 1677677812
transform 1 0 4112 0 1 1570
box -8 -3 16 105
use FILL  FILL_7936
timestamp 1677677812
transform 1 0 4120 0 1 1570
box -8 -3 16 105
use FILL  FILL_7937
timestamp 1677677812
transform 1 0 4128 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_293
timestamp 1677677812
transform 1 0 4136 0 1 1570
box -8 -3 46 105
use FILL  FILL_7938
timestamp 1677677812
transform 1 0 4176 0 1 1570
box -8 -3 16 105
use FILL  FILL_7950
timestamp 1677677812
transform 1 0 4184 0 1 1570
box -8 -3 16 105
use FILL  FILL_7952
timestamp 1677677812
transform 1 0 4192 0 1 1570
box -8 -3 16 105
use FILL  FILL_7954
timestamp 1677677812
transform 1 0 4200 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_294
timestamp 1677677812
transform 1 0 4208 0 1 1570
box -8 -3 46 105
use FILL  FILL_7956
timestamp 1677677812
transform 1 0 4248 0 1 1570
box -8 -3 16 105
use FILL  FILL_7960
timestamp 1677677812
transform 1 0 4256 0 1 1570
box -8 -3 16 105
use FILL  FILL_7962
timestamp 1677677812
transform 1 0 4264 0 1 1570
box -8 -3 16 105
use FILL  FILL_7964
timestamp 1677677812
transform 1 0 4272 0 1 1570
box -8 -3 16 105
use FILL  FILL_7966
timestamp 1677677812
transform 1 0 4280 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_295
timestamp 1677677812
transform 1 0 4288 0 1 1570
box -8 -3 46 105
use FILL  FILL_7968
timestamp 1677677812
transform 1 0 4328 0 1 1570
box -8 -3 16 105
use FILL  FILL_7971
timestamp 1677677812
transform 1 0 4336 0 1 1570
box -8 -3 16 105
use FILL  FILL_7973
timestamp 1677677812
transform 1 0 4344 0 1 1570
box -8 -3 16 105
use FILL  FILL_7975
timestamp 1677677812
transform 1 0 4352 0 1 1570
box -8 -3 16 105
use FILL  FILL_7977
timestamp 1677677812
transform 1 0 4360 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_296
timestamp 1677677812
transform 1 0 4368 0 1 1570
box -8 -3 46 105
use FILL  FILL_7978
timestamp 1677677812
transform 1 0 4408 0 1 1570
box -8 -3 16 105
use FILL  FILL_7982
timestamp 1677677812
transform 1 0 4416 0 1 1570
box -8 -3 16 105
use FILL  FILL_7984
timestamp 1677677812
transform 1 0 4424 0 1 1570
box -8 -3 16 105
use FILL  FILL_7986
timestamp 1677677812
transform 1 0 4432 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_297
timestamp 1677677812
transform -1 0 4480 0 1 1570
box -8 -3 46 105
use FILL  FILL_7987
timestamp 1677677812
transform 1 0 4480 0 1 1570
box -8 -3 16 105
use FILL  FILL_7988
timestamp 1677677812
transform 1 0 4488 0 1 1570
box -8 -3 16 105
use FILL  FILL_7989
timestamp 1677677812
transform 1 0 4496 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_298
timestamp 1677677812
transform -1 0 4544 0 1 1570
box -8 -3 46 105
use FILL  FILL_7990
timestamp 1677677812
transform 1 0 4544 0 1 1570
box -8 -3 16 105
use FILL  FILL_7991
timestamp 1677677812
transform 1 0 4552 0 1 1570
box -8 -3 16 105
use FILL  FILL_7992
timestamp 1677677812
transform 1 0 4560 0 1 1570
box -8 -3 16 105
use FILL  FILL_7993
timestamp 1677677812
transform 1 0 4568 0 1 1570
box -8 -3 16 105
use FILL  FILL_7994
timestamp 1677677812
transform 1 0 4576 0 1 1570
box -8 -3 16 105
use FILL  FILL_7995
timestamp 1677677812
transform 1 0 4584 0 1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_300
timestamp 1677677812
transform 1 0 4592 0 1 1570
box -8 -3 46 105
use FILL  FILL_8003
timestamp 1677677812
transform 1 0 4632 0 1 1570
box -8 -3 16 105
use FILL  FILL_8005
timestamp 1677677812
transform 1 0 4640 0 1 1570
box -8 -3 16 105
use FILL  FILL_8006
timestamp 1677677812
transform 1 0 4648 0 1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_430
timestamp 1677677812
transform 1 0 4656 0 1 1570
box -8 -3 104 105
use INVX2  INVX2_504
timestamp 1677677812
transform -1 0 4768 0 1 1570
box -9 -3 26 105
use FILL  FILL_8007
timestamp 1677677812
transform 1 0 4768 0 1 1570
box -8 -3 16 105
use FILL  FILL_8008
timestamp 1677677812
transform 1 0 4776 0 1 1570
box -8 -3 16 105
use FILL  FILL_8009
timestamp 1677677812
transform 1 0 4784 0 1 1570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_63
timestamp 1677677812
transform 1 0 4819 0 1 1570
box -10 -3 10 3
use M2_M1  M2_M1_6614
timestamp 1677677812
transform 1 0 84 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5964
timestamp 1677677812
transform 1 0 132 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5965
timestamp 1677677812
transform 1 0 172 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6706
timestamp 1677677812
transform 1 0 132 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6077
timestamp 1677677812
transform 1 0 156 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5909
timestamp 1677677812
transform 1 0 188 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6615
timestamp 1677677812
transform 1 0 188 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6616
timestamp 1677677812
transform 1 0 204 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5928
timestamp 1677677812
transform 1 0 308 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6617
timestamp 1677677812
transform 1 0 228 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5966
timestamp 1677677812
transform 1 0 324 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6707
timestamp 1677677812
transform 1 0 180 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6708
timestamp 1677677812
transform 1 0 196 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6709
timestamp 1677677812
transform 1 0 212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6710
timestamp 1677677812
transform 1 0 276 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6711
timestamp 1677677812
transform 1 0 308 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6712
timestamp 1677677812
transform 1 0 316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6713
timestamp 1677677812
transform 1 0 324 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6026
timestamp 1677677812
transform 1 0 212 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6027
timestamp 1677677812
transform 1 0 276 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6028
timestamp 1677677812
transform 1 0 316 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6054
timestamp 1677677812
transform 1 0 276 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6078
timestamp 1677677812
transform 1 0 236 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5996
timestamp 1677677812
transform 1 0 340 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6055
timestamp 1677677812
transform 1 0 340 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5910
timestamp 1677677812
transform 1 0 388 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5929
timestamp 1677677812
transform 1 0 380 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6618
timestamp 1677677812
transform 1 0 356 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6619
timestamp 1677677812
transform 1 0 364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6620
timestamp 1677677812
transform 1 0 380 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6621
timestamp 1677677812
transform 1 0 388 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6714
timestamp 1677677812
transform 1 0 356 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5997
timestamp 1677677812
transform 1 0 364 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6715
timestamp 1677677812
transform 1 0 372 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6716
timestamp 1677677812
transform 1 0 388 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6029
timestamp 1677677812
transform 1 0 356 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5894
timestamp 1677677812
transform 1 0 412 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5930
timestamp 1677677812
transform 1 0 452 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6622
timestamp 1677677812
transform 1 0 436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6623
timestamp 1677677812
transform 1 0 452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6717
timestamp 1677677812
transform 1 0 428 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6718
timestamp 1677677812
transform 1 0 444 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6624
timestamp 1677677812
transform 1 0 476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6719
timestamp 1677677812
transform 1 0 516 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6079
timestamp 1677677812
transform 1 0 516 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6080
timestamp 1677677812
transform 1 0 532 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5967
timestamp 1677677812
transform 1 0 564 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5931
timestamp 1677677812
transform 1 0 580 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6625
timestamp 1677677812
transform 1 0 572 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5932
timestamp 1677677812
transform 1 0 612 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6626
timestamp 1677677812
transform 1 0 588 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5968
timestamp 1677677812
transform 1 0 604 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6627
timestamp 1677677812
transform 1 0 612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6720
timestamp 1677677812
transform 1 0 580 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6721
timestamp 1677677812
transform 1 0 588 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6722
timestamp 1677677812
transform 1 0 604 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6723
timestamp 1677677812
transform 1 0 620 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6030
timestamp 1677677812
transform 1 0 588 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5911
timestamp 1677677812
transform 1 0 676 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6628
timestamp 1677677812
transform 1 0 676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6724
timestamp 1677677812
transform 1 0 668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6725
timestamp 1677677812
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6629
timestamp 1677677812
transform 1 0 804 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6726
timestamp 1677677812
transform 1 0 724 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6727
timestamp 1677677812
transform 1 0 772 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6031
timestamp 1677677812
transform 1 0 724 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6630
timestamp 1677677812
transform 1 0 820 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6032
timestamp 1677677812
transform 1 0 820 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6631
timestamp 1677677812
transform 1 0 868 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5969
timestamp 1677677812
transform 1 0 876 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6728
timestamp 1677677812
transform 1 0 844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6729
timestamp 1677677812
transform 1 0 860 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6730
timestamp 1677677812
transform 1 0 876 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6033
timestamp 1677677812
transform 1 0 876 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6056
timestamp 1677677812
transform 1 0 876 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5912
timestamp 1677677812
transform 1 0 892 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6607
timestamp 1677677812
transform 1 0 892 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6632
timestamp 1677677812
transform 1 0 916 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5998
timestamp 1677677812
transform 1 0 916 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5895
timestamp 1677677812
transform 1 0 932 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6608
timestamp 1677677812
transform 1 0 932 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_6057
timestamp 1677677812
transform 1 0 972 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5913
timestamp 1677677812
transform 1 0 988 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6731
timestamp 1677677812
transform 1 0 988 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6633
timestamp 1677677812
transform 1 0 1012 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6732
timestamp 1677677812
transform 1 0 1068 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6034
timestamp 1677677812
transform 1 0 1068 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6634
timestamp 1677677812
transform 1 0 1092 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6733
timestamp 1677677812
transform 1 0 1124 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6058
timestamp 1677677812
transform 1 0 1084 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6081
timestamp 1677677812
transform 1 0 1148 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_6082
timestamp 1677677812
transform 1 0 1180 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6734
timestamp 1677677812
transform 1 0 1204 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6059
timestamp 1677677812
transform 1 0 1212 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5896
timestamp 1677677812
transform 1 0 1236 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5897
timestamp 1677677812
transform 1 0 1268 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5933
timestamp 1677677812
transform 1 0 1236 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5934
timestamp 1677677812
transform 1 0 1260 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5970
timestamp 1677677812
transform 1 0 1228 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6635
timestamp 1677677812
transform 1 0 1236 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5971
timestamp 1677677812
transform 1 0 1244 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6636
timestamp 1677677812
transform 1 0 1252 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6637
timestamp 1677677812
transform 1 0 1260 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6735
timestamp 1677677812
transform 1 0 1220 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6736
timestamp 1677677812
transform 1 0 1244 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5999
timestamp 1677677812
transform 1 0 1252 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6737
timestamp 1677677812
transform 1 0 1260 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6060
timestamp 1677677812
transform 1 0 1228 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5935
timestamp 1677677812
transform 1 0 1292 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6000
timestamp 1677677812
transform 1 0 1284 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6738
timestamp 1677677812
transform 1 0 1292 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5914
timestamp 1677677812
transform 1 0 1324 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6638
timestamp 1677677812
transform 1 0 1324 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6001
timestamp 1677677812
transform 1 0 1308 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6739
timestamp 1677677812
transform 1 0 1316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6740
timestamp 1677677812
transform 1 0 1340 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5915
timestamp 1677677812
transform 1 0 1420 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5936
timestamp 1677677812
transform 1 0 1404 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6639
timestamp 1677677812
transform 1 0 1404 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5972
timestamp 1677677812
transform 1 0 1412 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6640
timestamp 1677677812
transform 1 0 1420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6741
timestamp 1677677812
transform 1 0 1396 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6002
timestamp 1677677812
transform 1 0 1404 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6742
timestamp 1677677812
transform 1 0 1412 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6003
timestamp 1677677812
transform 1 0 1420 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6641
timestamp 1677677812
transform 1 0 1436 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6004
timestamp 1677677812
transform 1 0 1436 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6743
timestamp 1677677812
transform 1 0 1444 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5916
timestamp 1677677812
transform 1 0 1540 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5937
timestamp 1677677812
transform 1 0 1492 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5973
timestamp 1677677812
transform 1 0 1484 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5974
timestamp 1677677812
transform 1 0 1524 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6642
timestamp 1677677812
transform 1 0 1572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6744
timestamp 1677677812
transform 1 0 1484 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6745
timestamp 1677677812
transform 1 0 1492 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6746
timestamp 1677677812
transform 1 0 1524 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6005
timestamp 1677677812
transform 1 0 1572 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6006
timestamp 1677677812
transform 1 0 1596 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5898
timestamp 1677677812
transform 1 0 1636 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6643
timestamp 1677677812
transform 1 0 1620 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6747
timestamp 1677677812
transform 1 0 1652 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6007
timestamp 1677677812
transform 1 0 1692 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6083
timestamp 1677677812
transform 1 0 1628 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6748
timestamp 1677677812
transform 1 0 1724 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5899
timestamp 1677677812
transform 1 0 1780 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6644
timestamp 1677677812
transform 1 0 1756 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6645
timestamp 1677677812
transform 1 0 1772 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6749
timestamp 1677677812
transform 1 0 1748 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6750
timestamp 1677677812
transform 1 0 1764 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6035
timestamp 1677677812
transform 1 0 1756 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6751
timestamp 1677677812
transform 1 0 1780 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5917
timestamp 1677677812
transform 1 0 1828 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5918
timestamp 1677677812
transform 1 0 1852 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6646
timestamp 1677677812
transform 1 0 1900 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6752
timestamp 1677677812
transform 1 0 1876 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6036
timestamp 1677677812
transform 1 0 1876 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5900
timestamp 1677677812
transform 1 0 1916 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6753
timestamp 1677677812
transform 1 0 1916 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6037
timestamp 1677677812
transform 1 0 1916 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6647
timestamp 1677677812
transform 1 0 1932 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6008
timestamp 1677677812
transform 1 0 1932 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6009
timestamp 1677677812
transform 1 0 1956 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5919
timestamp 1677677812
transform 1 0 1972 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6648
timestamp 1677677812
transform 1 0 1972 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6754
timestamp 1677677812
transform 1 0 2004 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6084
timestamp 1677677812
transform 1 0 2004 0 1 1485
box -3 -3 3 3
use M3_M2  M3_M2_5975
timestamp 1677677812
transform 1 0 2020 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6755
timestamp 1677677812
transform 1 0 2020 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6756
timestamp 1677677812
transform 1 0 2028 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5938
timestamp 1677677812
transform 1 0 2124 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6649
timestamp 1677677812
transform 1 0 2124 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5976
timestamp 1677677812
transform 1 0 2140 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6757
timestamp 1677677812
transform 1 0 2084 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6758
timestamp 1677677812
transform 1 0 2140 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6038
timestamp 1677677812
transform 1 0 2044 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6650
timestamp 1677677812
transform 1 0 2156 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6010
timestamp 1677677812
transform 1 0 2156 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6821
timestamp 1677677812
transform 1 0 2172 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_5939
timestamp 1677677812
transform 1 0 2212 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6759
timestamp 1677677812
transform 1 0 2204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6802
timestamp 1677677812
transform 1 0 2196 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6822
timestamp 1677677812
transform 1 0 2212 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_6085
timestamp 1677677812
transform 1 0 2212 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6803
timestamp 1677677812
transform 1 0 2236 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5901
timestamp 1677677812
transform 1 0 2260 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5940
timestamp 1677677812
transform 1 0 2300 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_6011
timestamp 1677677812
transform 1 0 2316 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6760
timestamp 1677677812
transform 1 0 2340 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5941
timestamp 1677677812
transform 1 0 2396 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5942
timestamp 1677677812
transform 1 0 2428 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6651
timestamp 1677677812
transform 1 0 2428 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6761
timestamp 1677677812
transform 1 0 2380 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6086
timestamp 1677677812
transform 1 0 2380 0 1 1485
box -3 -3 3 3
use M2_M1  M2_M1_6762
timestamp 1677677812
transform 1 0 2444 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5902
timestamp 1677677812
transform 1 0 2556 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5943
timestamp 1677677812
transform 1 0 2572 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6652
timestamp 1677677812
transform 1 0 2572 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6763
timestamp 1677677812
transform 1 0 2548 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6072
timestamp 1677677812
transform 1 0 2532 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_6073
timestamp 1677677812
transform 1 0 2556 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6764
timestamp 1677677812
transform 1 0 2588 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6039
timestamp 1677677812
transform 1 0 2596 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5944
timestamp 1677677812
transform 1 0 2684 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5945
timestamp 1677677812
transform 1 0 2732 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5946
timestamp 1677677812
transform 1 0 2780 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5977
timestamp 1677677812
transform 1 0 2740 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6653
timestamp 1677677812
transform 1 0 2780 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6012
timestamp 1677677812
transform 1 0 2748 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6765
timestamp 1677677812
transform 1 0 2756 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6040
timestamp 1677677812
transform 1 0 2756 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6013
timestamp 1677677812
transform 1 0 2796 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5947
timestamp 1677677812
transform 1 0 2812 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6804
timestamp 1677677812
transform 1 0 2796 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6041
timestamp 1677677812
transform 1 0 2804 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6823
timestamp 1677677812
transform 1 0 2812 0 1 1505
box -2 -2 2 2
use M2_M1  M2_M1_6766
timestamp 1677677812
transform 1 0 2844 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5948
timestamp 1677677812
transform 1 0 2868 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6654
timestamp 1677677812
transform 1 0 2868 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6767
timestamp 1677677812
transform 1 0 2868 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6805
timestamp 1677677812
transform 1 0 2884 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6061
timestamp 1677677812
transform 1 0 2884 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6609
timestamp 1677677812
transform 1 0 3028 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_5949
timestamp 1677677812
transform 1 0 3052 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6655
timestamp 1677677812
transform 1 0 2916 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6656
timestamp 1677677812
transform 1 0 2924 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5978
timestamp 1677677812
transform 1 0 2932 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6657
timestamp 1677677812
transform 1 0 3036 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5979
timestamp 1677677812
transform 1 0 3044 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6658
timestamp 1677677812
transform 1 0 3052 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6659
timestamp 1677677812
transform 1 0 3060 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6014
timestamp 1677677812
transform 1 0 2916 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6768
timestamp 1677677812
transform 1 0 2924 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6769
timestamp 1677677812
transform 1 0 2940 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6770
timestamp 1677677812
transform 1 0 3044 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6806
timestamp 1677677812
transform 1 0 2916 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6042
timestamp 1677677812
transform 1 0 2924 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6062
timestamp 1677677812
transform 1 0 2916 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6063
timestamp 1677677812
transform 1 0 3020 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6064
timestamp 1677677812
transform 1 0 3044 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6015
timestamp 1677677812
transform 1 0 3076 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5950
timestamp 1677677812
transform 1 0 3100 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6660
timestamp 1677677812
transform 1 0 3100 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5951
timestamp 1677677812
transform 1 0 3148 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6661
timestamp 1677677812
transform 1 0 3148 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6807
timestamp 1677677812
transform 1 0 3140 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6610
timestamp 1677677812
transform 1 0 3180 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6662
timestamp 1677677812
transform 1 0 3172 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6043
timestamp 1677677812
transform 1 0 3172 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6663
timestamp 1677677812
transform 1 0 3188 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5903
timestamp 1677677812
transform 1 0 3212 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5920
timestamp 1677677812
transform 1 0 3260 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6611
timestamp 1677677812
transform 1 0 3316 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_5952
timestamp 1677677812
transform 1 0 3324 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6664
timestamp 1677677812
transform 1 0 3212 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5980
timestamp 1677677812
transform 1 0 3228 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5981
timestamp 1677677812
transform 1 0 3268 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6771
timestamp 1677677812
transform 1 0 3204 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6772
timestamp 1677677812
transform 1 0 3212 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6773
timestamp 1677677812
transform 1 0 3228 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6016
timestamp 1677677812
transform 1 0 3316 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6044
timestamp 1677677812
transform 1 0 3212 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6065
timestamp 1677677812
transform 1 0 3260 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_6066
timestamp 1677677812
transform 1 0 3284 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6665
timestamp 1677677812
transform 1 0 3332 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5953
timestamp 1677677812
transform 1 0 3340 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6666
timestamp 1677677812
transform 1 0 3340 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6017
timestamp 1677677812
transform 1 0 3332 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6774
timestamp 1677677812
transform 1 0 3372 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5921
timestamp 1677677812
transform 1 0 3404 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6612
timestamp 1677677812
transform 1 0 3404 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6667
timestamp 1677677812
transform 1 0 3420 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6775
timestamp 1677677812
transform 1 0 3444 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5904
timestamp 1677677812
transform 1 0 3460 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6668
timestamp 1677677812
transform 1 0 3460 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6776
timestamp 1677677812
transform 1 0 3468 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6067
timestamp 1677677812
transform 1 0 3460 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5922
timestamp 1677677812
transform 1 0 3492 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6669
timestamp 1677677812
transform 1 0 3492 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6018
timestamp 1677677812
transform 1 0 3484 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6777
timestamp 1677677812
transform 1 0 3500 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6613
timestamp 1677677812
transform 1 0 3516 0 1 1545
box -2 -2 2 2
use M2_M1  M2_M1_6670
timestamp 1677677812
transform 1 0 3572 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6045
timestamp 1677677812
transform 1 0 3556 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6068
timestamp 1677677812
transform 1 0 3548 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6671
timestamp 1677677812
transform 1 0 3588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6778
timestamp 1677677812
transform 1 0 3580 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6046
timestamp 1677677812
transform 1 0 3580 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6779
timestamp 1677677812
transform 1 0 3612 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5954
timestamp 1677677812
transform 1 0 3668 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6780
timestamp 1677677812
transform 1 0 3668 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6781
timestamp 1677677812
transform 1 0 3676 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6672
timestamp 1677677812
transform 1 0 3692 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6074
timestamp 1677677812
transform 1 0 3692 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5982
timestamp 1677677812
transform 1 0 3700 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6673
timestamp 1677677812
transform 1 0 3708 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5983
timestamp 1677677812
transform 1 0 3732 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6674
timestamp 1677677812
transform 1 0 3740 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6019
timestamp 1677677812
transform 1 0 3716 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6782
timestamp 1677677812
transform 1 0 3732 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6808
timestamp 1677677812
transform 1 0 3716 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6675
timestamp 1677677812
transform 1 0 3796 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5984
timestamp 1677677812
transform 1 0 3812 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6783
timestamp 1677677812
transform 1 0 3812 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6020
timestamp 1677677812
transform 1 0 3828 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6784
timestamp 1677677812
transform 1 0 3844 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6809
timestamp 1677677812
transform 1 0 3828 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6047
timestamp 1677677812
transform 1 0 3844 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5905
timestamp 1677677812
transform 1 0 3876 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6676
timestamp 1677677812
transform 1 0 3876 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5985
timestamp 1677677812
transform 1 0 3884 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6785
timestamp 1677677812
transform 1 0 3876 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6677
timestamp 1677677812
transform 1 0 3908 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6786
timestamp 1677677812
transform 1 0 3908 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6069
timestamp 1677677812
transform 1 0 3908 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_5923
timestamp 1677677812
transform 1 0 3932 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6678
timestamp 1677677812
transform 1 0 3924 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6679
timestamp 1677677812
transform 1 0 3932 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6810
timestamp 1677677812
transform 1 0 3964 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6680
timestamp 1677677812
transform 1 0 4036 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6048
timestamp 1677677812
transform 1 0 4028 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_5986
timestamp 1677677812
transform 1 0 4052 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6787
timestamp 1677677812
transform 1 0 4052 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6021
timestamp 1677677812
transform 1 0 4068 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_6049
timestamp 1677677812
transform 1 0 4052 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_6811
timestamp 1677677812
transform 1 0 4068 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6681
timestamp 1677677812
transform 1 0 4076 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5987
timestamp 1677677812
transform 1 0 4084 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6682
timestamp 1677677812
transform 1 0 4100 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5988
timestamp 1677677812
transform 1 0 4116 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6683
timestamp 1677677812
transform 1 0 4124 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6684
timestamp 1677677812
transform 1 0 4132 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_6022
timestamp 1677677812
transform 1 0 4100 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6788
timestamp 1677677812
transform 1 0 4116 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6023
timestamp 1677677812
transform 1 0 4132 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6812
timestamp 1677677812
transform 1 0 4132 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5955
timestamp 1677677812
transform 1 0 4148 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5989
timestamp 1677677812
transform 1 0 4156 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6789
timestamp 1677677812
transform 1 0 4148 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5956
timestamp 1677677812
transform 1 0 4196 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6685
timestamp 1677677812
transform 1 0 4196 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5906
timestamp 1677677812
transform 1 0 4244 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_6686
timestamp 1677677812
transform 1 0 4228 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5990
timestamp 1677677812
transform 1 0 4236 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6687
timestamp 1677677812
transform 1 0 4244 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6813
timestamp 1677677812
transform 1 0 4260 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6814
timestamp 1677677812
transform 1 0 4268 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6075
timestamp 1677677812
transform 1 0 4268 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_5924
timestamp 1677677812
transform 1 0 4332 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6688
timestamp 1677677812
transform 1 0 4324 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6689
timestamp 1677677812
transform 1 0 4332 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6790
timestamp 1677677812
transform 1 0 4316 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6815
timestamp 1677677812
transform 1 0 4300 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6690
timestamp 1677677812
transform 1 0 4396 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6791
timestamp 1677677812
transform 1 0 4388 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6816
timestamp 1677677812
transform 1 0 4372 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6070
timestamp 1677677812
transform 1 0 4372 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6817
timestamp 1677677812
transform 1 0 4404 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6071
timestamp 1677677812
transform 1 0 4404 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_6818
timestamp 1677677812
transform 1 0 4420 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_5957
timestamp 1677677812
transform 1 0 4476 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6691
timestamp 1677677812
transform 1 0 4444 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5991
timestamp 1677677812
transform 1 0 4452 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6692
timestamp 1677677812
transform 1 0 4476 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6792
timestamp 1677677812
transform 1 0 4460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6793
timestamp 1677677812
transform 1 0 4476 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6819
timestamp 1677677812
transform 1 0 4444 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_6820
timestamp 1677677812
transform 1 0 4484 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_6076
timestamp 1677677812
transform 1 0 4484 0 1 1495
box -3 -3 3 3
use M2_M1  M2_M1_6693
timestamp 1677677812
transform 1 0 4508 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5992
timestamp 1677677812
transform 1 0 4516 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6694
timestamp 1677677812
transform 1 0 4524 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5958
timestamp 1677677812
transform 1 0 4548 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6695
timestamp 1677677812
transform 1 0 4548 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6696
timestamp 1677677812
transform 1 0 4564 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5993
timestamp 1677677812
transform 1 0 4572 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_6794
timestamp 1677677812
transform 1 0 4556 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6795
timestamp 1677677812
transform 1 0 4572 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_5925
timestamp 1677677812
transform 1 0 4588 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5926
timestamp 1677677812
transform 1 0 4628 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_5959
timestamp 1677677812
transform 1 0 4596 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5960
timestamp 1677677812
transform 1 0 4612 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5961
timestamp 1677677812
transform 1 0 4636 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_5962
timestamp 1677677812
transform 1 0 4668 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6697
timestamp 1677677812
transform 1 0 4588 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6698
timestamp 1677677812
transform 1 0 4596 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6699
timestamp 1677677812
transform 1 0 4612 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6700
timestamp 1677677812
transform 1 0 4628 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6796
timestamp 1677677812
transform 1 0 4604 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6797
timestamp 1677677812
transform 1 0 4620 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6701
timestamp 1677677812
transform 1 0 4644 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6702
timestamp 1677677812
transform 1 0 4660 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5994
timestamp 1677677812
transform 1 0 4668 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_5907
timestamp 1677677812
transform 1 0 4700 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5908
timestamp 1677677812
transform 1 0 4724 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_5963
timestamp 1677677812
transform 1 0 4692 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6703
timestamp 1677677812
transform 1 0 4676 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6704
timestamp 1677677812
transform 1 0 4692 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_5995
timestamp 1677677812
transform 1 0 4716 0 1 1535
box -3 -3 3 3
use M3_M2  M3_M2_6024
timestamp 1677677812
transform 1 0 4652 0 1 1525
box -3 -3 3 3
use M2_M1  M2_M1_6798
timestamp 1677677812
transform 1 0 4668 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6025
timestamp 1677677812
transform 1 0 4676 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_5927
timestamp 1677677812
transform 1 0 4796 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_6705
timestamp 1677677812
transform 1 0 4788 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_6799
timestamp 1677677812
transform 1 0 4716 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6800
timestamp 1677677812
transform 1 0 4772 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_6801
timestamp 1677677812
transform 1 0 4796 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_6050
timestamp 1677677812
transform 1 0 4668 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6051
timestamp 1677677812
transform 1 0 4724 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6052
timestamp 1677677812
transform 1 0 4772 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_6053
timestamp 1677677812
transform 1 0 4788 0 1 1515
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_64
timestamp 1677677812
transform 1 0 24 0 1 1470
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_411
timestamp 1677677812
transform 1 0 72 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7552
timestamp 1677677812
transform 1 0 168 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_283
timestamp 1677677812
transform -1 0 216 0 -1 1570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_412
timestamp 1677677812
transform 1 0 216 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_483
timestamp 1677677812
transform -1 0 328 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7553
timestamp 1677677812
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7554
timestamp 1677677812
transform 1 0 336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7559
timestamp 1677677812
transform 1 0 344 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_285
timestamp 1677677812
transform 1 0 352 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7560
timestamp 1677677812
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7561
timestamp 1677677812
transform 1 0 400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7562
timestamp 1677677812
transform 1 0 408 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_280
timestamp 1677677812
transform -1 0 456 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7563
timestamp 1677677812
transform 1 0 456 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6087
timestamp 1677677812
transform 1 0 484 0 1 1475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_414
timestamp 1677677812
transform 1 0 464 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7564
timestamp 1677677812
transform 1 0 560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7568
timestamp 1677677812
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7569
timestamp 1677677812
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_287
timestamp 1677677812
transform 1 0 584 0 -1 1570
box -8 -3 46 105
use M3_M2  M3_M2_6088
timestamp 1677677812
transform 1 0 636 0 1 1475
box -3 -3 3 3
use FILL  FILL_7570
timestamp 1677677812
transform 1 0 624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7572
timestamp 1677677812
transform 1 0 632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7574
timestamp 1677677812
transform 1 0 640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7576
timestamp 1677677812
transform 1 0 648 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_281
timestamp 1677677812
transform 1 0 656 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7583
timestamp 1677677812
transform 1 0 696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7585
timestamp 1677677812
transform 1 0 704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7598
timestamp 1677677812
transform 1 0 712 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_415
timestamp 1677677812
transform -1 0 816 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7599
timestamp 1677677812
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7600
timestamp 1677677812
transform 1 0 824 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7601
timestamp 1677677812
transform 1 0 832 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_289
timestamp 1677677812
transform -1 0 880 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7602
timestamp 1677677812
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7603
timestamp 1677677812
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7604
timestamp 1677677812
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7606
timestamp 1677677812
transform 1 0 904 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_74
timestamp 1677677812
transform 1 0 912 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7610
timestamp 1677677812
transform 1 0 936 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7611
timestamp 1677677812
transform 1 0 944 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7612
timestamp 1677677812
transform 1 0 952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7613
timestamp 1677677812
transform 1 0 960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7614
timestamp 1677677812
transform 1 0 968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7615
timestamp 1677677812
transform 1 0 976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7616
timestamp 1677677812
transform 1 0 984 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_75
timestamp 1677677812
transform 1 0 992 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7617
timestamp 1677677812
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7618
timestamp 1677677812
transform 1 0 1024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7620
timestamp 1677677812
transform 1 0 1032 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7622
timestamp 1677677812
transform 1 0 1040 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7625
timestamp 1677677812
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7626
timestamp 1677677812
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7627
timestamp 1677677812
transform 1 0 1064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7628
timestamp 1677677812
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_417
timestamp 1677677812
transform 1 0 1080 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7637
timestamp 1677677812
transform 1 0 1176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7639
timestamp 1677677812
transform 1 0 1184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7641
timestamp 1677677812
transform 1 0 1192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7643
timestamp 1677677812
transform 1 0 1200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7645
timestamp 1677677812
transform 1 0 1208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7651
timestamp 1677677812
transform 1 0 1216 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_291
timestamp 1677677812
transform -1 0 1264 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7652
timestamp 1677677812
transform 1 0 1264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7653
timestamp 1677677812
transform 1 0 1272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7654
timestamp 1677677812
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7655
timestamp 1677677812
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7673
timestamp 1677677812
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_283
timestamp 1677677812
transform -1 0 1344 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7674
timestamp 1677677812
transform 1 0 1344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7675
timestamp 1677677812
transform 1 0 1352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7676
timestamp 1677677812
transform 1 0 1360 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6089
timestamp 1677677812
transform 1 0 1380 0 1 1475
box -3 -3 3 3
use FILL  FILL_7677
timestamp 1677677812
transform 1 0 1368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7678
timestamp 1677677812
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7679
timestamp 1677677812
transform 1 0 1384 0 -1 1570
box -8 -3 16 105
use AOI22X1  AOI22X1_293
timestamp 1677677812
transform -1 0 1432 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7680
timestamp 1677677812
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7681
timestamp 1677677812
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_490
timestamp 1677677812
transform 1 0 1448 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7682
timestamp 1677677812
transform 1 0 1464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7683
timestamp 1677677812
transform 1 0 1472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7684
timestamp 1677677812
transform 1 0 1480 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_419
timestamp 1677677812
transform -1 0 1584 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7685
timestamp 1677677812
transform 1 0 1584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7686
timestamp 1677677812
transform 1 0 1592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7688
timestamp 1677677812
transform 1 0 1600 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6090
timestamp 1677677812
transform 1 0 1676 0 1 1475
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_420
timestamp 1677677812
transform 1 0 1608 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7694
timestamp 1677677812
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7695
timestamp 1677677812
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7696
timestamp 1677677812
transform 1 0 1720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7710
timestamp 1677677812
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_285
timestamp 1677677812
transform -1 0 1776 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7711
timestamp 1677677812
transform 1 0 1776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7712
timestamp 1677677812
transform 1 0 1784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7713
timestamp 1677677812
transform 1 0 1792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7714
timestamp 1677677812
transform 1 0 1800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7715
timestamp 1677677812
transform 1 0 1808 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_422
timestamp 1677677812
transform -1 0 1912 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7716
timestamp 1677677812
transform 1 0 1912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7717
timestamp 1677677812
transform 1 0 1920 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7718
timestamp 1677677812
transform 1 0 1928 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7719
timestamp 1677677812
transform 1 0 1936 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_491
timestamp 1677677812
transform 1 0 1944 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7720
timestamp 1677677812
transform 1 0 1960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7723
timestamp 1677677812
transform 1 0 1968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7724
timestamp 1677677812
transform 1 0 1976 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6091
timestamp 1677677812
transform 1 0 2004 0 1 1475
box -3 -3 3 3
use BUFX2  BUFX2_94
timestamp 1677677812
transform -1 0 2008 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7725
timestamp 1677677812
transform 1 0 2008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7727
timestamp 1677677812
transform 1 0 2016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7729
timestamp 1677677812
transform 1 0 2024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7741
timestamp 1677677812
transform 1 0 2032 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_423
timestamp 1677677812
transform -1 0 2136 0 -1 1570
box -8 -3 104 105
use BUFX2  BUFX2_97
timestamp 1677677812
transform 1 0 2136 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7742
timestamp 1677677812
transform 1 0 2160 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6092
timestamp 1677677812
transform 1 0 2180 0 1 1475
box -3 -3 3 3
use FILL  FILL_7744
timestamp 1677677812
transform 1 0 2168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7746
timestamp 1677677812
transform 1 0 2176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7748
timestamp 1677677812
transform 1 0 2184 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_55
timestamp 1677677812
transform 1 0 2192 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7751
timestamp 1677677812
transform 1 0 2224 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7752
timestamp 1677677812
transform 1 0 2232 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7753
timestamp 1677677812
transform 1 0 2240 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7754
timestamp 1677677812
transform 1 0 2248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7755
timestamp 1677677812
transform 1 0 2256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7756
timestamp 1677677812
transform 1 0 2264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7757
timestamp 1677677812
transform 1 0 2272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7758
timestamp 1677677812
transform 1 0 2280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7759
timestamp 1677677812
transform 1 0 2288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7760
timestamp 1677677812
transform 1 0 2296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7762
timestamp 1677677812
transform 1 0 2304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7783
timestamp 1677677812
transform 1 0 2312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7784
timestamp 1677677812
transform 1 0 2320 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6093
timestamp 1677677812
transform 1 0 2340 0 1 1475
box -3 -3 3 3
use FILL  FILL_7785
timestamp 1677677812
transform 1 0 2328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7786
timestamp 1677677812
transform 1 0 2336 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_427
timestamp 1677677812
transform -1 0 2440 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7787
timestamp 1677677812
transform 1 0 2440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7788
timestamp 1677677812
transform 1 0 2448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7789
timestamp 1677677812
transform 1 0 2456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7790
timestamp 1677677812
transform 1 0 2464 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7791
timestamp 1677677812
transform 1 0 2472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7792
timestamp 1677677812
transform 1 0 2480 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_428
timestamp 1677677812
transform -1 0 2584 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7793
timestamp 1677677812
transform 1 0 2584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7794
timestamp 1677677812
transform 1 0 2592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7795
timestamp 1677677812
transform 1 0 2600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7796
timestamp 1677677812
transform 1 0 2608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7797
timestamp 1677677812
transform 1 0 2616 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7798
timestamp 1677677812
transform 1 0 2624 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7799
timestamp 1677677812
transform 1 0 2632 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7800
timestamp 1677677812
transform 1 0 2640 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7801
timestamp 1677677812
transform 1 0 2648 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7802
timestamp 1677677812
transform 1 0 2656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7803
timestamp 1677677812
transform 1 0 2664 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7804
timestamp 1677677812
transform 1 0 2672 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7805
timestamp 1677677812
transform 1 0 2680 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7806
timestamp 1677677812
transform 1 0 2688 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_429
timestamp 1677677812
transform -1 0 2792 0 -1 1570
box -8 -3 104 105
use FILL  FILL_7807
timestamp 1677677812
transform 1 0 2792 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7808
timestamp 1677677812
transform 1 0 2800 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7809
timestamp 1677677812
transform 1 0 2808 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7810
timestamp 1677677812
transform 1 0 2816 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7812
timestamp 1677677812
transform 1 0 2824 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_57
timestamp 1677677812
transform 1 0 2832 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7816
timestamp 1677677812
transform 1 0 2864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7818
timestamp 1677677812
transform 1 0 2872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7820
timestamp 1677677812
transform 1 0 2880 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_130
timestamp 1677677812
transform 1 0 2888 0 -1 1570
box -8 -3 34 105
use FAX1  FAX1_1
timestamp 1677677812
transform 1 0 2920 0 -1 1570
box -5 -3 126 105
use INVX2  INVX2_497
timestamp 1677677812
transform -1 0 3056 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7835
timestamp 1677677812
transform 1 0 3056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7836
timestamp 1677677812
transform 1 0 3064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7837
timestamp 1677677812
transform 1 0 3072 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_498
timestamp 1677677812
transform 1 0 3080 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7838
timestamp 1677677812
transform 1 0 3096 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_131
timestamp 1677677812
transform 1 0 3104 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7839
timestamp 1677677812
transform 1 0 3136 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7842
timestamp 1677677812
transform 1 0 3144 0 -1 1570
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1677677812
transform -1 0 3184 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7843
timestamp 1677677812
transform 1 0 3184 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_500
timestamp 1677677812
transform 1 0 3192 0 -1 1570
box -9 -3 26 105
use FAX1  FAX1_2
timestamp 1677677812
transform 1 0 3208 0 -1 1570
box -5 -3 126 105
use FILL  FILL_7857
timestamp 1677677812
transform 1 0 3328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7858
timestamp 1677677812
transform 1 0 3336 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1677677812
transform 1 0 3344 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7859
timestamp 1677677812
transform 1 0 3368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7868
timestamp 1677677812
transform 1 0 3376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7869
timestamp 1677677812
transform 1 0 3384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7870
timestamp 1677677812
transform 1 0 3392 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_3
timestamp 1677677812
transform -1 0 3432 0 -1 1570
box -7 -3 39 105
use FILL  FILL_7871
timestamp 1677677812
transform 1 0 3432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7872
timestamp 1677677812
transform 1 0 3440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7873
timestamp 1677677812
transform 1 0 3448 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7874
timestamp 1677677812
transform 1 0 3456 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7875
timestamp 1677677812
transform 1 0 3464 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_286
timestamp 1677677812
transform 1 0 3472 0 -1 1570
box -8 -3 46 105
use FILL  FILL_7876
timestamp 1677677812
transform 1 0 3512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7877
timestamp 1677677812
transform 1 0 3520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7878
timestamp 1677677812
transform 1 0 3528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7879
timestamp 1677677812
transform 1 0 3536 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7886
timestamp 1677677812
transform 1 0 3544 0 -1 1570
box -8 -3 16 105
use AOI21X1  AOI21X1_4
timestamp 1677677812
transform -1 0 3584 0 -1 1570
box -7 -3 39 105
use FILL  FILL_7887
timestamp 1677677812
transform 1 0 3584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7888
timestamp 1677677812
transform 1 0 3592 0 -1 1570
box -8 -3 16 105
use AND2X2  AND2X2_50
timestamp 1677677812
transform 1 0 3600 0 -1 1570
box -8 -3 40 105
use FILL  FILL_7889
timestamp 1677677812
transform 1 0 3632 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_502
timestamp 1677677812
transform 1 0 3640 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7890
timestamp 1677677812
transform 1 0 3656 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7891
timestamp 1677677812
transform 1 0 3664 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_503
timestamp 1677677812
transform -1 0 3688 0 -1 1570
box -9 -3 26 105
use FILL  FILL_7892
timestamp 1677677812
transform 1 0 3688 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7893
timestamp 1677677812
transform 1 0 3696 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7894
timestamp 1677677812
transform 1 0 3704 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_132
timestamp 1677677812
transform -1 0 3744 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7895
timestamp 1677677812
transform 1 0 3744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7897
timestamp 1677677812
transform 1 0 3752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7907
timestamp 1677677812
transform 1 0 3760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7908
timestamp 1677677812
transform 1 0 3768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7909
timestamp 1677677812
transform 1 0 3776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7910
timestamp 1677677812
transform 1 0 3784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7911
timestamp 1677677812
transform 1 0 3792 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_133
timestamp 1677677812
transform 1 0 3800 0 -1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_7
timestamp 1677677812
transform -1 0 3856 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7912
timestamp 1677677812
transform 1 0 3856 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7913
timestamp 1677677812
transform 1 0 3864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7914
timestamp 1677677812
transform 1 0 3872 0 -1 1570
box -8 -3 16 105
use BUFX2  BUFX2_99
timestamp 1677677812
transform 1 0 3880 0 -1 1570
box -5 -3 28 105
use FILL  FILL_7915
timestamp 1677677812
transform 1 0 3904 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7917
timestamp 1677677812
transform 1 0 3912 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7919
timestamp 1677677812
transform 1 0 3920 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_8
timestamp 1677677812
transform 1 0 3928 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7922
timestamp 1677677812
transform 1 0 3952 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7923
timestamp 1677677812
transform 1 0 3960 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7924
timestamp 1677677812
transform 1 0 3968 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7925
timestamp 1677677812
transform 1 0 3976 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7927
timestamp 1677677812
transform 1 0 3984 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7929
timestamp 1677677812
transform 1 0 3992 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7931
timestamp 1677677812
transform 1 0 4000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7939
timestamp 1677677812
transform 1 0 4008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7940
timestamp 1677677812
transform 1 0 4016 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7941
timestamp 1677677812
transform 1 0 4024 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7942
timestamp 1677677812
transform 1 0 4032 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_134
timestamp 1677677812
transform 1 0 4040 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7943
timestamp 1677677812
transform 1 0 4072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7944
timestamp 1677677812
transform 1 0 4080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7945
timestamp 1677677812
transform 1 0 4088 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_135
timestamp 1677677812
transform -1 0 4128 0 -1 1570
box -8 -3 34 105
use NAND2X1  NAND2X1_9
timestamp 1677677812
transform -1 0 4152 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7946
timestamp 1677677812
transform 1 0 4152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7947
timestamp 1677677812
transform 1 0 4160 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7948
timestamp 1677677812
transform 1 0 4168 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7949
timestamp 1677677812
transform 1 0 4176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7951
timestamp 1677677812
transform 1 0 4184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7953
timestamp 1677677812
transform 1 0 4192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7955
timestamp 1677677812
transform 1 0 4200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7957
timestamp 1677677812
transform 1 0 4208 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7958
timestamp 1677677812
transform 1 0 4216 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_10
timestamp 1677677812
transform 1 0 4224 0 -1 1570
box -8 -3 32 105
use FILL  FILL_7959
timestamp 1677677812
transform 1 0 4248 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7961
timestamp 1677677812
transform 1 0 4256 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7963
timestamp 1677677812
transform 1 0 4264 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7965
timestamp 1677677812
transform 1 0 4272 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7967
timestamp 1677677812
transform 1 0 4280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7969
timestamp 1677677812
transform 1 0 4288 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_136
timestamp 1677677812
transform -1 0 4328 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7970
timestamp 1677677812
transform 1 0 4328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7972
timestamp 1677677812
transform 1 0 4336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7974
timestamp 1677677812
transform 1 0 4344 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7976
timestamp 1677677812
transform 1 0 4352 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7979
timestamp 1677677812
transform 1 0 4360 0 -1 1570
box -8 -3 16 105
use M3_M2  M3_M2_6094
timestamp 1677677812
transform 1 0 4380 0 1 1475
box -3 -3 3 3
use OAI21X1  OAI21X1_137
timestamp 1677677812
transform -1 0 4400 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7980
timestamp 1677677812
transform 1 0 4400 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7981
timestamp 1677677812
transform 1 0 4408 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7983
timestamp 1677677812
transform 1 0 4416 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7985
timestamp 1677677812
transform 1 0 4424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7996
timestamp 1677677812
transform 1 0 4432 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_138
timestamp 1677677812
transform -1 0 4472 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7997
timestamp 1677677812
transform 1 0 4472 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_139
timestamp 1677677812
transform -1 0 4512 0 -1 1570
box -8 -3 34 105
use FILL  FILL_7998
timestamp 1677677812
transform 1 0 4512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7999
timestamp 1677677812
transform 1 0 4520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8000
timestamp 1677677812
transform 1 0 4528 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8001
timestamp 1677677812
transform 1 0 4536 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_299
timestamp 1677677812
transform 1 0 4544 0 -1 1570
box -8 -3 46 105
use FILL  FILL_8002
timestamp 1677677812
transform 1 0 4584 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_301
timestamp 1677677812
transform 1 0 4592 0 -1 1570
box -8 -3 46 105
use FILL  FILL_8004
timestamp 1677677812
transform 1 0 4632 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_302
timestamp 1677677812
transform 1 0 4640 0 -1 1570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_431
timestamp 1677677812
transform 1 0 4680 0 -1 1570
box -8 -3 104 105
use INVX2  INVX2_505
timestamp 1677677812
transform -1 0 4792 0 -1 1570
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_65
timestamp 1677677812
transform 1 0 4843 0 1 1470
box -10 -3 10 3
use M3_M2  M3_M2_6110
timestamp 1677677812
transform 1 0 116 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6111
timestamp 1677677812
transform 1 0 148 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6123
timestamp 1677677812
transform 1 0 164 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6144
timestamp 1677677812
transform 1 0 132 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6145
timestamp 1677677812
transform 1 0 172 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6845
timestamp 1677677812
transform 1 0 132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6846
timestamp 1677677812
transform 1 0 164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6847
timestamp 1677677812
transform 1 0 172 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6848
timestamp 1677677812
transform 1 0 180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6849
timestamp 1677677812
transform 1 0 188 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6946
timestamp 1677677812
transform 1 0 84 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6210
timestamp 1677677812
transform 1 0 148 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6211
timestamp 1677677812
transform 1 0 164 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6124
timestamp 1677677812
transform 1 0 204 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6850
timestamp 1677677812
transform 1 0 212 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6947
timestamp 1677677812
transform 1 0 196 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6948
timestamp 1677677812
transform 1 0 204 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6949
timestamp 1677677812
transform 1 0 220 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6950
timestamp 1677677812
transform 1 0 244 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6102
timestamp 1677677812
transform 1 0 316 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6125
timestamp 1677677812
transform 1 0 308 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6851
timestamp 1677677812
transform 1 0 268 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6852
timestamp 1677677812
transform 1 0 284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6853
timestamp 1677677812
transform 1 0 300 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6951
timestamp 1677677812
transform 1 0 276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6952
timestamp 1677677812
transform 1 0 292 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6854
timestamp 1677677812
transform 1 0 372 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6855
timestamp 1677677812
transform 1 0 380 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6953
timestamp 1677677812
transform 1 0 404 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6095
timestamp 1677677812
transform 1 0 420 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6096
timestamp 1677677812
transform 1 0 476 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6097
timestamp 1677677812
transform 1 0 492 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6103
timestamp 1677677812
transform 1 0 428 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6112
timestamp 1677677812
transform 1 0 436 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6146
timestamp 1677677812
transform 1 0 468 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6856
timestamp 1677677812
transform 1 0 468 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6857
timestamp 1677677812
transform 1 0 500 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6858
timestamp 1677677812
transform 1 0 508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6954
timestamp 1677677812
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6230
timestamp 1677677812
transform 1 0 500 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6261
timestamp 1677677812
transform 1 0 444 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6147
timestamp 1677677812
transform 1 0 516 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6859
timestamp 1677677812
transform 1 0 516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6955
timestamp 1677677812
transform 1 0 516 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6148
timestamp 1677677812
transform 1 0 540 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6860
timestamp 1677677812
transform 1 0 532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6956
timestamp 1677677812
transform 1 0 540 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6126
timestamp 1677677812
transform 1 0 556 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6861
timestamp 1677677812
transform 1 0 556 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6176
timestamp 1677677812
transform 1 0 572 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6149
timestamp 1677677812
transform 1 0 596 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6862
timestamp 1677677812
transform 1 0 596 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6177
timestamp 1677677812
transform 1 0 604 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6863
timestamp 1677677812
transform 1 0 612 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6957
timestamp 1677677812
transform 1 0 572 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6958
timestamp 1677677812
transform 1 0 580 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6959
timestamp 1677677812
transform 1 0 612 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6960
timestamp 1677677812
transform 1 0 620 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6231
timestamp 1677677812
transform 1 0 612 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6864
timestamp 1677677812
transform 1 0 636 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6262
timestamp 1677677812
transform 1 0 620 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6178
timestamp 1677677812
transform 1 0 652 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6961
timestamp 1677677812
transform 1 0 644 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6232
timestamp 1677677812
transform 1 0 644 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6263
timestamp 1677677812
transform 1 0 644 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6865
timestamp 1677677812
transform 1 0 676 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6179
timestamp 1677677812
transform 1 0 684 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6866
timestamp 1677677812
transform 1 0 692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6962
timestamp 1677677812
transform 1 0 684 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6212
timestamp 1677677812
transform 1 0 692 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6963
timestamp 1677677812
transform 1 0 700 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6233
timestamp 1677677812
transform 1 0 700 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6867
timestamp 1677677812
transform 1 0 740 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6127
timestamp 1677677812
transform 1 0 772 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6868
timestamp 1677677812
transform 1 0 772 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6150
timestamp 1677677812
transform 1 0 812 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6869
timestamp 1677677812
transform 1 0 812 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6180
timestamp 1677677812
transform 1 0 820 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6113
timestamp 1677677812
transform 1 0 852 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6870
timestamp 1677677812
transform 1 0 828 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6871
timestamp 1677677812
transform 1 0 844 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6964
timestamp 1677677812
transform 1 0 812 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6965
timestamp 1677677812
transform 1 0 820 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6966
timestamp 1677677812
transform 1 0 836 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6234
timestamp 1677677812
transform 1 0 836 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7027
timestamp 1677677812
transform 1 0 852 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6181
timestamp 1677677812
transform 1 0 868 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7028
timestamp 1677677812
transform 1 0 892 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6264
timestamp 1677677812
transform 1 0 892 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6967
timestamp 1677677812
transform 1 0 908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6872
timestamp 1677677812
transform 1 0 932 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6213
timestamp 1677677812
transform 1 0 948 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7029
timestamp 1677677812
transform 1 0 948 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6265
timestamp 1677677812
transform 1 0 948 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6968
timestamp 1677677812
transform 1 0 964 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6266
timestamp 1677677812
transform 1 0 980 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6873
timestamp 1677677812
transform 1 0 996 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6267
timestamp 1677677812
transform 1 0 996 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6969
timestamp 1677677812
transform 1 0 1052 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6128
timestamp 1677677812
transform 1 0 1092 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6874
timestamp 1677677812
transform 1 0 1092 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6214
timestamp 1677677812
transform 1 0 1092 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6151
timestamp 1677677812
transform 1 0 1132 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6875
timestamp 1677677812
transform 1 0 1124 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6876
timestamp 1677677812
transform 1 0 1132 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6152
timestamp 1677677812
transform 1 0 1164 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6970
timestamp 1677677812
transform 1 0 1164 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6235
timestamp 1677677812
transform 1 0 1156 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7030
timestamp 1677677812
transform 1 0 1164 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6114
timestamp 1677677812
transform 1 0 1188 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6182
timestamp 1677677812
transform 1 0 1180 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6877
timestamp 1677677812
transform 1 0 1188 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6183
timestamp 1677677812
transform 1 0 1196 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6878
timestamp 1677677812
transform 1 0 1204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6879
timestamp 1677677812
transform 1 0 1220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6971
timestamp 1677677812
transform 1 0 1212 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6236
timestamp 1677677812
transform 1 0 1196 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6153
timestamp 1677677812
transform 1 0 1244 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6184
timestamp 1677677812
transform 1 0 1244 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6129
timestamp 1677677812
transform 1 0 1260 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6880
timestamp 1677677812
transform 1 0 1276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6881
timestamp 1677677812
transform 1 0 1292 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6185
timestamp 1677677812
transform 1 0 1300 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6882
timestamp 1677677812
transform 1 0 1308 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6215
timestamp 1677677812
transform 1 0 1292 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6972
timestamp 1677677812
transform 1 0 1300 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6154
timestamp 1677677812
transform 1 0 1404 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6883
timestamp 1677677812
transform 1 0 1388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6884
timestamp 1677677812
transform 1 0 1404 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6885
timestamp 1677677812
transform 1 0 1420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6973
timestamp 1677677812
transform 1 0 1396 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6237
timestamp 1677677812
transform 1 0 1396 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6115
timestamp 1677677812
transform 1 0 1436 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6116
timestamp 1677677812
transform 1 0 1452 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6886
timestamp 1677677812
transform 1 0 1444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6974
timestamp 1677677812
transform 1 0 1436 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6268
timestamp 1677677812
transform 1 0 1452 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6155
timestamp 1677677812
transform 1 0 1460 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6975
timestamp 1677677812
transform 1 0 1460 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6156
timestamp 1677677812
transform 1 0 1508 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6157
timestamp 1677677812
transform 1 0 1548 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6887
timestamp 1677677812
transform 1 0 1508 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6888
timestamp 1677677812
transform 1 0 1516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6889
timestamp 1677677812
transform 1 0 1548 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6976
timestamp 1677677812
transform 1 0 1596 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6238
timestamp 1677677812
transform 1 0 1516 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6239
timestamp 1677677812
transform 1 0 1580 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6890
timestamp 1677677812
transform 1 0 1652 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6240
timestamp 1677677812
transform 1 0 1668 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6891
timestamp 1677677812
transform 1 0 1676 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6186
timestamp 1677677812
transform 1 0 1708 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6892
timestamp 1677677812
transform 1 0 1716 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6893
timestamp 1677677812
transform 1 0 1732 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6977
timestamp 1677677812
transform 1 0 1700 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6978
timestamp 1677677812
transform 1 0 1708 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6979
timestamp 1677677812
transform 1 0 1724 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6216
timestamp 1677677812
transform 1 0 1732 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6894
timestamp 1677677812
transform 1 0 1756 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6130
timestamp 1677677812
transform 1 0 1772 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6895
timestamp 1677677812
transform 1 0 1772 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6117
timestamp 1677677812
transform 1 0 1860 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6158
timestamp 1677677812
transform 1 0 1836 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6896
timestamp 1677677812
transform 1 0 1836 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6187
timestamp 1677677812
transform 1 0 1860 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6980
timestamp 1677677812
transform 1 0 1860 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6241
timestamp 1677677812
transform 1 0 1812 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6242
timestamp 1677677812
transform 1 0 1844 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6159
timestamp 1677677812
transform 1 0 1876 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6897
timestamp 1677677812
transform 1 0 1876 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6188
timestamp 1677677812
transform 1 0 1900 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6898
timestamp 1677677812
transform 1 0 1924 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6104
timestamp 1677677812
transform 1 0 1948 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6160
timestamp 1677677812
transform 1 0 1964 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6899
timestamp 1677677812
transform 1 0 1964 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6131
timestamp 1677677812
transform 1 0 1980 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6161
timestamp 1677677812
transform 1 0 1996 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6900
timestamp 1677677812
transform 1 0 1988 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6901
timestamp 1677677812
transform 1 0 2004 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6981
timestamp 1677677812
transform 1 0 1972 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6982
timestamp 1677677812
transform 1 0 1980 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6983
timestamp 1677677812
transform 1 0 1996 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6984
timestamp 1677677812
transform 1 0 2020 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6105
timestamp 1677677812
transform 1 0 2036 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6162
timestamp 1677677812
transform 1 0 2092 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6902
timestamp 1677677812
transform 1 0 2092 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6985
timestamp 1677677812
transform 1 0 2116 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6824
timestamp 1677677812
transform 1 0 2172 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_6826
timestamp 1677677812
transform 1 0 2164 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6189
timestamp 1677677812
transform 1 0 2164 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6986
timestamp 1677677812
transform 1 0 2180 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6132
timestamp 1677677812
transform 1 0 2196 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6827
timestamp 1677677812
transform 1 0 2196 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6217
timestamp 1677677812
transform 1 0 2204 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6133
timestamp 1677677812
transform 1 0 2252 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6903
timestamp 1677677812
transform 1 0 2220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6904
timestamp 1677677812
transform 1 0 2252 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6218
timestamp 1677677812
transform 1 0 2252 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6987
timestamp 1677677812
transform 1 0 2300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6905
timestamp 1677677812
transform 1 0 2388 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6906
timestamp 1677677812
transform 1 0 2420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6988
timestamp 1677677812
transform 1 0 2340 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6243
timestamp 1677677812
transform 1 0 2420 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6190
timestamp 1677677812
transform 1 0 2524 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6907
timestamp 1677677812
transform 1 0 2540 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6989
timestamp 1677677812
transform 1 0 2556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7031
timestamp 1677677812
transform 1 0 2452 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6244
timestamp 1677677812
transform 1 0 2556 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6163
timestamp 1677677812
transform 1 0 2636 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6191
timestamp 1677677812
transform 1 0 2588 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6908
timestamp 1677677812
transform 1 0 2636 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6192
timestamp 1677677812
transform 1 0 2660 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6990
timestamp 1677677812
transform 1 0 2660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6909
timestamp 1677677812
transform 1 0 2676 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6193
timestamp 1677677812
transform 1 0 2684 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6910
timestamp 1677677812
transform 1 0 2740 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6194
timestamp 1677677812
transform 1 0 2764 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6991
timestamp 1677677812
transform 1 0 2764 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6245
timestamp 1677677812
transform 1 0 2740 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6164
timestamp 1677677812
transform 1 0 2788 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6195
timestamp 1677677812
transform 1 0 2780 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6911
timestamp 1677677812
transform 1 0 2788 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6992
timestamp 1677677812
transform 1 0 2788 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6246
timestamp 1677677812
transform 1 0 2788 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6912
timestamp 1677677812
transform 1 0 2812 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7032
timestamp 1677677812
transform 1 0 2900 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6118
timestamp 1677677812
transform 1 0 2916 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6196
timestamp 1677677812
transform 1 0 2932 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7037
timestamp 1677677812
transform 1 0 2940 0 1 1385
box -2 -2 2 2
use M3_M2  M3_M2_6098
timestamp 1677677812
transform 1 0 2964 0 1 1465
box -3 -3 3 3
use M2_M1  M2_M1_7038
timestamp 1677677812
transform 1 0 2972 0 1 1385
box -2 -2 2 2
use M3_M2  M3_M2_6247
timestamp 1677677812
transform 1 0 2996 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6165
timestamp 1677677812
transform 1 0 3012 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6825
timestamp 1677677812
transform 1 0 3052 0 1 1435
box -2 -2 2 2
use M3_M2  M3_M2_6134
timestamp 1677677812
transform 1 0 3060 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6828
timestamp 1677677812
transform 1 0 3044 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6166
timestamp 1677677812
transform 1 0 3052 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6913
timestamp 1677677812
transform 1 0 3060 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6219
timestamp 1677677812
transform 1 0 3044 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6269
timestamp 1677677812
transform 1 0 3068 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6119
timestamp 1677677812
transform 1 0 3084 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6197
timestamp 1677677812
transform 1 0 3084 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6993
timestamp 1677677812
transform 1 0 3084 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6135
timestamp 1677677812
transform 1 0 3092 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6829
timestamp 1677677812
transform 1 0 3092 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6994
timestamp 1677677812
transform 1 0 3116 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6248
timestamp 1677677812
transform 1 0 3116 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6167
timestamp 1677677812
transform 1 0 3132 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6830
timestamp 1677677812
transform 1 0 3140 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6914
timestamp 1677677812
transform 1 0 3132 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6220
timestamp 1677677812
transform 1 0 3132 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6168
timestamp 1677677812
transform 1 0 3164 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6915
timestamp 1677677812
transform 1 0 3164 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6198
timestamp 1677677812
transform 1 0 3172 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6995
timestamp 1677677812
transform 1 0 3172 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6106
timestamp 1677677812
transform 1 0 3220 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6136
timestamp 1677677812
transform 1 0 3220 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6916
timestamp 1677677812
transform 1 0 3204 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6917
timestamp 1677677812
transform 1 0 3220 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6221
timestamp 1677677812
transform 1 0 3212 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6996
timestamp 1677677812
transform 1 0 3228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6997
timestamp 1677677812
transform 1 0 3236 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6270
timestamp 1677677812
transform 1 0 3236 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6107
timestamp 1677677812
transform 1 0 3252 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_6918
timestamp 1677677812
transform 1 0 3276 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6919
timestamp 1677677812
transform 1 0 3284 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6271
timestamp 1677677812
transform 1 0 3276 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6222
timestamp 1677677812
transform 1 0 3300 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6249
timestamp 1677677812
transform 1 0 3292 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7033
timestamp 1677677812
transform 1 0 3324 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_7034
timestamp 1677677812
transform 1 0 3332 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6108
timestamp 1677677812
transform 1 0 3364 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_6920
timestamp 1677677812
transform 1 0 3340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6921
timestamp 1677677812
transform 1 0 3348 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6199
timestamp 1677677812
transform 1 0 3356 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6998
timestamp 1677677812
transform 1 0 3364 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6120
timestamp 1677677812
transform 1 0 3380 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6999
timestamp 1677677812
transform 1 0 3380 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6223
timestamp 1677677812
transform 1 0 3396 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6099
timestamp 1677677812
transform 1 0 3524 0 1 1465
box -3 -3 3 3
use M3_M2  M3_M2_6121
timestamp 1677677812
transform 1 0 3412 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_6137
timestamp 1677677812
transform 1 0 3444 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6138
timestamp 1677677812
transform 1 0 3532 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6922
timestamp 1677677812
transform 1 0 3412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6923
timestamp 1677677812
transform 1 0 3420 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6924
timestamp 1677677812
transform 1 0 3524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7000
timestamp 1677677812
transform 1 0 3404 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6250
timestamp 1677677812
transform 1 0 3388 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6224
timestamp 1677677812
transform 1 0 3412 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6109
timestamp 1677677812
transform 1 0 3572 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_6139
timestamp 1677677812
transform 1 0 3588 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_6140
timestamp 1677677812
transform 1 0 3612 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6925
timestamp 1677677812
transform 1 0 3556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6926
timestamp 1677677812
transform 1 0 3564 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6200
timestamp 1677677812
transform 1 0 3652 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6831
timestamp 1677677812
transform 1 0 3668 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6927
timestamp 1677677812
transform 1 0 3668 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7001
timestamp 1677677812
transform 1 0 3516 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7002
timestamp 1677677812
transform 1 0 3540 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7003
timestamp 1677677812
transform 1 0 3548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7004
timestamp 1677677812
transform 1 0 3660 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7035
timestamp 1677677812
transform 1 0 3508 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6251
timestamp 1677677812
transform 1 0 3516 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6272
timestamp 1677677812
transform 1 0 3508 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6273
timestamp 1677677812
transform 1 0 3532 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6252
timestamp 1677677812
transform 1 0 3564 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_7036
timestamp 1677677812
transform 1 0 3652 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_6253
timestamp 1677677812
transform 1 0 3660 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6274
timestamp 1677677812
transform 1 0 3564 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6141
timestamp 1677677812
transform 1 0 3692 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6832
timestamp 1677677812
transform 1 0 3684 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6254
timestamp 1677677812
transform 1 0 3684 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6833
timestamp 1677677812
transform 1 0 3708 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6201
timestamp 1677677812
transform 1 0 3724 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6202
timestamp 1677677812
transform 1 0 3756 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7005
timestamp 1677677812
transform 1 0 3748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7006
timestamp 1677677812
transform 1 0 3756 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6275
timestamp 1677677812
transform 1 0 3748 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6928
timestamp 1677677812
transform 1 0 3780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6834
timestamp 1677677812
transform 1 0 3820 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6203
timestamp 1677677812
transform 1 0 3820 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6100
timestamp 1677677812
transform 1 0 3844 0 1 1465
box -3 -3 3 3
use M2_M1  M2_M1_6929
timestamp 1677677812
transform 1 0 3836 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6930
timestamp 1677677812
transform 1 0 3844 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6101
timestamp 1677677812
transform 1 0 3876 0 1 1465
box -3 -3 3 3
use M2_M1  M2_M1_7007
timestamp 1677677812
transform 1 0 3868 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7008
timestamp 1677677812
transform 1 0 3892 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7009
timestamp 1677677812
transform 1 0 3908 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6835
timestamp 1677677812
transform 1 0 3956 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6931
timestamp 1677677812
transform 1 0 3940 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6204
timestamp 1677677812
transform 1 0 3956 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6932
timestamp 1677677812
transform 1 0 3972 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7010
timestamp 1677677812
transform 1 0 3964 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6225
timestamp 1677677812
transform 1 0 3972 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7011
timestamp 1677677812
transform 1 0 4004 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6255
timestamp 1677677812
transform 1 0 4004 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6122
timestamp 1677677812
transform 1 0 4020 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_6933
timestamp 1677677812
transform 1 0 4020 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6169
timestamp 1677677812
transform 1 0 4060 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6836
timestamp 1677677812
transform 1 0 4068 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6837
timestamp 1677677812
transform 1 0 4076 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6205
timestamp 1677677812
transform 1 0 4076 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_6170
timestamp 1677677812
transform 1 0 4124 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6206
timestamp 1677677812
transform 1 0 4116 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7012
timestamp 1677677812
transform 1 0 4116 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6226
timestamp 1677677812
transform 1 0 4124 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_6171
timestamp 1677677812
transform 1 0 4140 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6172
timestamp 1677677812
transform 1 0 4236 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6838
timestamp 1677677812
transform 1 0 4252 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6934
timestamp 1677677812
transform 1 0 4164 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6935
timestamp 1677677812
transform 1 0 4220 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6936
timestamp 1677677812
transform 1 0 4228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7013
timestamp 1677677812
transform 1 0 4140 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6227
timestamp 1677677812
transform 1 0 4164 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7014
timestamp 1677677812
transform 1 0 4228 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7015
timestamp 1677677812
transform 1 0 4260 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6937
timestamp 1677677812
transform 1 0 4276 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6228
timestamp 1677677812
transform 1 0 4284 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_6938
timestamp 1677677812
transform 1 0 4356 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6229
timestamp 1677677812
transform 1 0 4356 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_7016
timestamp 1677677812
transform 1 0 4404 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7017
timestamp 1677677812
transform 1 0 4420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6256
timestamp 1677677812
transform 1 0 4420 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6839
timestamp 1677677812
transform 1 0 4444 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_7018
timestamp 1677677812
transform 1 0 4468 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6840
timestamp 1677677812
transform 1 0 4484 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_7019
timestamp 1677677812
transform 1 0 4484 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6173
timestamp 1677677812
transform 1 0 4500 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6257
timestamp 1677677812
transform 1 0 4492 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6276
timestamp 1677677812
transform 1 0 4484 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_6939
timestamp 1677677812
transform 1 0 4516 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6142
timestamp 1677677812
transform 1 0 4524 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6841
timestamp 1677677812
transform 1 0 4524 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6258
timestamp 1677677812
transform 1 0 4524 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_6842
timestamp 1677677812
transform 1 0 4556 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6207
timestamp 1677677812
transform 1 0 4556 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_7020
timestamp 1677677812
transform 1 0 4548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7021
timestamp 1677677812
transform 1 0 4556 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6843
timestamp 1677677812
transform 1 0 4572 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_6143
timestamp 1677677812
transform 1 0 4588 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_6844
timestamp 1677677812
transform 1 0 4588 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_6940
timestamp 1677677812
transform 1 0 4596 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7022
timestamp 1677677812
transform 1 0 4620 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_6941
timestamp 1677677812
transform 1 0 4636 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_6174
timestamp 1677677812
transform 1 0 4668 0 1 1425
box -3 -3 3 3
use M3_M2  M3_M2_6175
timestamp 1677677812
transform 1 0 4692 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_6942
timestamp 1677677812
transform 1 0 4652 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6943
timestamp 1677677812
transform 1 0 4692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_6944
timestamp 1677677812
transform 1 0 4748 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7023
timestamp 1677677812
transform 1 0 4636 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7024
timestamp 1677677812
transform 1 0 4644 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_7025
timestamp 1677677812
transform 1 0 4668 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6259
timestamp 1677677812
transform 1 0 4668 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6260
timestamp 1677677812
transform 1 0 4692 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_6277
timestamp 1677677812
transform 1 0 4652 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6278
timestamp 1677677812
transform 1 0 4684 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_6208
timestamp 1677677812
transform 1 0 4764 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_6945
timestamp 1677677812
transform 1 0 4772 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_7026
timestamp 1677677812
transform 1 0 4764 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_6209
timestamp 1677677812
transform 1 0 4788 0 1 1415
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_66
timestamp 1677677812
transform 1 0 48 0 1 1370
box -10 -3 10 3
use M3_M2  M3_M2_6279
timestamp 1677677812
transform 1 0 92 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6280
timestamp 1677677812
transform 1 0 124 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_432
timestamp 1677677812
transform 1 0 72 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_506
timestamp 1677677812
transform -1 0 184 0 1 1370
box -9 -3 26 105
use FILL  FILL_8010
timestamp 1677677812
transform 1 0 184 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_296
timestamp 1677677812
transform -1 0 232 0 1 1370
box -8 -3 46 105
use FILL  FILL_8011
timestamp 1677677812
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_8021
timestamp 1677677812
transform 1 0 240 0 1 1370
box -8 -3 16 105
use FILL  FILL_8022
timestamp 1677677812
transform 1 0 248 0 1 1370
box -8 -3 16 105
use FILL  FILL_8023
timestamp 1677677812
transform 1 0 256 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_297
timestamp 1677677812
transform 1 0 264 0 1 1370
box -8 -3 46 105
use FILL  FILL_8024
timestamp 1677677812
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_8025
timestamp 1677677812
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8026
timestamp 1677677812
transform 1 0 320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8027
timestamp 1677677812
transform 1 0 328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8028
timestamp 1677677812
transform 1 0 336 0 1 1370
box -8 -3 16 105
use FILL  FILL_8029
timestamp 1677677812
transform 1 0 344 0 1 1370
box -8 -3 16 105
use FILL  FILL_8030
timestamp 1677677812
transform 1 0 352 0 1 1370
box -8 -3 16 105
use FILL  FILL_8031
timestamp 1677677812
transform 1 0 360 0 1 1370
box -8 -3 16 105
use FILL  FILL_8032
timestamp 1677677812
transform 1 0 368 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_507
timestamp 1677677812
transform -1 0 392 0 1 1370
box -9 -3 26 105
use FILL  FILL_8033
timestamp 1677677812
transform 1 0 392 0 1 1370
box -8 -3 16 105
use FILL  FILL_8034
timestamp 1677677812
transform 1 0 400 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_434
timestamp 1677677812
transform 1 0 408 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_508
timestamp 1677677812
transform -1 0 520 0 1 1370
box -9 -3 26 105
use INVX2  INVX2_509
timestamp 1677677812
transform -1 0 536 0 1 1370
box -9 -3 26 105
use FILL  FILL_8035
timestamp 1677677812
transform 1 0 536 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_510
timestamp 1677677812
transform -1 0 560 0 1 1370
box -9 -3 26 105
use FILL  FILL_8036
timestamp 1677677812
transform 1 0 560 0 1 1370
box -8 -3 16 105
use FILL  FILL_8037
timestamp 1677677812
transform 1 0 568 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_298
timestamp 1677677812
transform 1 0 576 0 1 1370
box -8 -3 46 105
use BUFX2  BUFX2_100
timestamp 1677677812
transform -1 0 640 0 1 1370
box -5 -3 28 105
use FILL  FILL_8038
timestamp 1677677812
transform 1 0 640 0 1 1370
box -8 -3 16 105
use FILL  FILL_8039
timestamp 1677677812
transform 1 0 648 0 1 1370
box -8 -3 16 105
use FILL  FILL_8040
timestamp 1677677812
transform 1 0 656 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_303
timestamp 1677677812
transform 1 0 664 0 1 1370
box -8 -3 46 105
use FILL  FILL_8041
timestamp 1677677812
transform 1 0 704 0 1 1370
box -8 -3 16 105
use FILL  FILL_8042
timestamp 1677677812
transform 1 0 712 0 1 1370
box -8 -3 16 105
use FILL  FILL_8043
timestamp 1677677812
transform 1 0 720 0 1 1370
box -8 -3 16 105
use FILL  FILL_8044
timestamp 1677677812
transform 1 0 728 0 1 1370
box -8 -3 16 105
use FILL  FILL_8045
timestamp 1677677812
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_8046
timestamp 1677677812
transform 1 0 744 0 1 1370
box -8 -3 16 105
use FILL  FILL_8047
timestamp 1677677812
transform 1 0 752 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_511
timestamp 1677677812
transform -1 0 776 0 1 1370
box -9 -3 26 105
use FILL  FILL_8048
timestamp 1677677812
transform 1 0 776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8064
timestamp 1677677812
transform 1 0 784 0 1 1370
box -8 -3 16 105
use FILL  FILL_8066
timestamp 1677677812
transform 1 0 792 0 1 1370
box -8 -3 16 105
use FILL  FILL_8068
timestamp 1677677812
transform 1 0 800 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_300
timestamp 1677677812
transform 1 0 808 0 1 1370
box -8 -3 46 105
use FILL  FILL_8070
timestamp 1677677812
transform 1 0 848 0 1 1370
box -8 -3 16 105
use FILL  FILL_8077
timestamp 1677677812
transform 1 0 856 0 1 1370
box -8 -3 16 105
use FILL  FILL_8079
timestamp 1677677812
transform 1 0 864 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_81
timestamp 1677677812
transform 1 0 872 0 1 1370
box -8 -3 32 105
use FILL  FILL_8081
timestamp 1677677812
transform 1 0 896 0 1 1370
box -8 -3 16 105
use FILL  FILL_8086
timestamp 1677677812
transform 1 0 904 0 1 1370
box -8 -3 16 105
use FILL  FILL_8088
timestamp 1677677812
transform 1 0 912 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6281
timestamp 1677677812
transform 1 0 932 0 1 1375
box -3 -3 3 3
use FILL  FILL_8090
timestamp 1677677812
transform 1 0 920 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_82
timestamp 1677677812
transform 1 0 928 0 1 1370
box -8 -3 32 105
use FILL  FILL_8092
timestamp 1677677812
transform 1 0 952 0 1 1370
box -8 -3 16 105
use FILL  FILL_8093
timestamp 1677677812
transform 1 0 960 0 1 1370
box -8 -3 16 105
use FILL  FILL_8094
timestamp 1677677812
transform 1 0 968 0 1 1370
box -8 -3 16 105
use FILL  FILL_8098
timestamp 1677677812
transform 1 0 976 0 1 1370
box -8 -3 16 105
use FILL  FILL_8100
timestamp 1677677812
transform 1 0 984 0 1 1370
box -8 -3 16 105
use FILL  FILL_8102
timestamp 1677677812
transform 1 0 992 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_84
timestamp 1677677812
transform 1 0 1000 0 1 1370
box -8 -3 32 105
use FILL  FILL_8104
timestamp 1677677812
transform 1 0 1024 0 1 1370
box -8 -3 16 105
use FILL  FILL_8105
timestamp 1677677812
transform 1 0 1032 0 1 1370
box -8 -3 16 105
use FILL  FILL_8106
timestamp 1677677812
transform 1 0 1040 0 1 1370
box -8 -3 16 105
use FILL  FILL_8111
timestamp 1677677812
transform 1 0 1048 0 1 1370
box -8 -3 16 105
use FILL  FILL_8113
timestamp 1677677812
transform 1 0 1056 0 1 1370
box -8 -3 16 105
use FILL  FILL_8115
timestamp 1677677812
transform 1 0 1064 0 1 1370
box -8 -3 16 105
use FILL  FILL_8117
timestamp 1677677812
transform 1 0 1072 0 1 1370
box -8 -3 16 105
use FILL  FILL_8119
timestamp 1677677812
transform 1 0 1080 0 1 1370
box -8 -3 16 105
use FILL  FILL_8121
timestamp 1677677812
transform 1 0 1088 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_514
timestamp 1677677812
transform -1 0 1112 0 1 1370
box -9 -3 26 105
use FILL  FILL_8122
timestamp 1677677812
transform 1 0 1112 0 1 1370
box -8 -3 16 105
use FILL  FILL_8127
timestamp 1677677812
transform 1 0 1120 0 1 1370
box -8 -3 16 105
use FILL  FILL_8129
timestamp 1677677812
transform 1 0 1128 0 1 1370
box -8 -3 16 105
use FILL  FILL_8131
timestamp 1677677812
transform 1 0 1136 0 1 1370
box -8 -3 16 105
use FILL  FILL_8133
timestamp 1677677812
transform 1 0 1144 0 1 1370
box -8 -3 16 105
use FILL  FILL_8135
timestamp 1677677812
transform 1 0 1152 0 1 1370
box -8 -3 16 105
use FILL  FILL_8137
timestamp 1677677812
transform 1 0 1160 0 1 1370
box -8 -3 16 105
use FILL  FILL_8139
timestamp 1677677812
transform 1 0 1168 0 1 1370
box -8 -3 16 105
use FILL  FILL_8141
timestamp 1677677812
transform 1 0 1176 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_301
timestamp 1677677812
transform 1 0 1184 0 1 1370
box -8 -3 46 105
use FILL  FILL_8143
timestamp 1677677812
transform 1 0 1224 0 1 1370
box -8 -3 16 105
use FILL  FILL_8147
timestamp 1677677812
transform 1 0 1232 0 1 1370
box -8 -3 16 105
use FILL  FILL_8149
timestamp 1677677812
transform 1 0 1240 0 1 1370
box -8 -3 16 105
use FILL  FILL_8150
timestamp 1677677812
transform 1 0 1248 0 1 1370
box -8 -3 16 105
use FILL  FILL_8151
timestamp 1677677812
transform 1 0 1256 0 1 1370
box -8 -3 16 105
use FILL  FILL_8152
timestamp 1677677812
transform 1 0 1264 0 1 1370
box -8 -3 16 105
use FILL  FILL_8153
timestamp 1677677812
transform 1 0 1272 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_306
timestamp 1677677812
transform -1 0 1320 0 1 1370
box -8 -3 46 105
use FILL  FILL_8154
timestamp 1677677812
transform 1 0 1320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8155
timestamp 1677677812
transform 1 0 1328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8156
timestamp 1677677812
transform 1 0 1336 0 1 1370
box -8 -3 16 105
use FILL  FILL_8157
timestamp 1677677812
transform 1 0 1344 0 1 1370
box -8 -3 16 105
use FILL  FILL_8158
timestamp 1677677812
transform 1 0 1352 0 1 1370
box -8 -3 16 105
use FILL  FILL_8159
timestamp 1677677812
transform 1 0 1360 0 1 1370
box -8 -3 16 105
use FILL  FILL_8160
timestamp 1677677812
transform 1 0 1368 0 1 1370
box -8 -3 16 105
use FILL  FILL_8161
timestamp 1677677812
transform 1 0 1376 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_302
timestamp 1677677812
transform -1 0 1424 0 1 1370
box -8 -3 46 105
use FILL  FILL_8162
timestamp 1677677812
transform 1 0 1424 0 1 1370
box -8 -3 16 105
use FILL  FILL_8163
timestamp 1677677812
transform 1 0 1432 0 1 1370
box -8 -3 16 105
use FILL  FILL_8164
timestamp 1677677812
transform 1 0 1440 0 1 1370
box -8 -3 16 105
use FILL  FILL_8165
timestamp 1677677812
transform 1 0 1448 0 1 1370
box -8 -3 16 105
use FILL  FILL_8166
timestamp 1677677812
transform 1 0 1456 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_515
timestamp 1677677812
transform 1 0 1464 0 1 1370
box -9 -3 26 105
use FILL  FILL_8167
timestamp 1677677812
transform 1 0 1480 0 1 1370
box -8 -3 16 105
use FILL  FILL_8177
timestamp 1677677812
transform 1 0 1488 0 1 1370
box -8 -3 16 105
use FILL  FILL_8178
timestamp 1677677812
transform 1 0 1496 0 1 1370
box -8 -3 16 105
use FILL  FILL_8179
timestamp 1677677812
transform 1 0 1504 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_439
timestamp 1677677812
transform -1 0 1608 0 1 1370
box -8 -3 104 105
use FILL  FILL_8180
timestamp 1677677812
transform 1 0 1608 0 1 1370
box -8 -3 16 105
use FILL  FILL_8181
timestamp 1677677812
transform 1 0 1616 0 1 1370
box -8 -3 16 105
use FILL  FILL_8182
timestamp 1677677812
transform 1 0 1624 0 1 1370
box -8 -3 16 105
use FILL  FILL_8183
timestamp 1677677812
transform 1 0 1632 0 1 1370
box -8 -3 16 105
use FILL  FILL_8188
timestamp 1677677812
transform 1 0 1640 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6282
timestamp 1677677812
transform 1 0 1668 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_516
timestamp 1677677812
transform -1 0 1664 0 1 1370
box -9 -3 26 105
use FILL  FILL_8189
timestamp 1677677812
transform 1 0 1664 0 1 1370
box -8 -3 16 105
use FILL  FILL_8190
timestamp 1677677812
transform 1 0 1672 0 1 1370
box -8 -3 16 105
use FILL  FILL_8191
timestamp 1677677812
transform 1 0 1680 0 1 1370
box -8 -3 16 105
use FILL  FILL_8192
timestamp 1677677812
transform 1 0 1688 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_304
timestamp 1677677812
transform 1 0 1696 0 1 1370
box -8 -3 46 105
use FILL  FILL_8195
timestamp 1677677812
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_8196
timestamp 1677677812
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_8197
timestamp 1677677812
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_8198
timestamp 1677677812
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_8203
timestamp 1677677812
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_441
timestamp 1677677812
transform -1 0 1872 0 1 1370
box -8 -3 104 105
use FILL  FILL_8204
timestamp 1677677812
transform 1 0 1872 0 1 1370
box -8 -3 16 105
use FILL  FILL_8205
timestamp 1677677812
transform 1 0 1880 0 1 1370
box -8 -3 16 105
use FILL  FILL_8209
timestamp 1677677812
transform 1 0 1888 0 1 1370
box -8 -3 16 105
use FILL  FILL_8211
timestamp 1677677812
transform 1 0 1896 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_517
timestamp 1677677812
transform -1 0 1920 0 1 1370
box -9 -3 26 105
use FILL  FILL_8212
timestamp 1677677812
transform 1 0 1920 0 1 1370
box -8 -3 16 105
use FILL  FILL_8217
timestamp 1677677812
transform 1 0 1928 0 1 1370
box -8 -3 16 105
use FILL  FILL_8219
timestamp 1677677812
transform 1 0 1936 0 1 1370
box -8 -3 16 105
use FILL  FILL_8220
timestamp 1677677812
transform 1 0 1944 0 1 1370
box -8 -3 16 105
use FILL  FILL_8221
timestamp 1677677812
transform 1 0 1952 0 1 1370
box -8 -3 16 105
use FILL  FILL_8222
timestamp 1677677812
transform 1 0 1960 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_306
timestamp 1677677812
transform -1 0 2008 0 1 1370
box -8 -3 46 105
use FILL  FILL_8223
timestamp 1677677812
transform 1 0 2008 0 1 1370
box -8 -3 16 105
use FILL  FILL_8224
timestamp 1677677812
transform 1 0 2016 0 1 1370
box -8 -3 16 105
use FILL  FILL_8225
timestamp 1677677812
transform 1 0 2024 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_443
timestamp 1677677812
transform -1 0 2128 0 1 1370
box -8 -3 104 105
use FILL  FILL_8226
timestamp 1677677812
transform 1 0 2128 0 1 1370
box -8 -3 16 105
use FILL  FILL_8227
timestamp 1677677812
transform 1 0 2136 0 1 1370
box -8 -3 16 105
use FILL  FILL_8228
timestamp 1677677812
transform 1 0 2144 0 1 1370
box -8 -3 16 105
use FILL  FILL_8237
timestamp 1677677812
transform 1 0 2152 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_62
timestamp 1677677812
transform -1 0 2192 0 1 1370
box -8 -3 40 105
use FILL  FILL_8239
timestamp 1677677812
transform 1 0 2192 0 1 1370
box -8 -3 16 105
use FILL  FILL_8240
timestamp 1677677812
transform 1 0 2200 0 1 1370
box -8 -3 16 105
use FILL  FILL_8241
timestamp 1677677812
transform 1 0 2208 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_445
timestamp 1677677812
transform -1 0 2312 0 1 1370
box -8 -3 104 105
use FILL  FILL_8242
timestamp 1677677812
transform 1 0 2312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8243
timestamp 1677677812
transform 1 0 2320 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_446
timestamp 1677677812
transform 1 0 2328 0 1 1370
box -8 -3 104 105
use FILL  FILL_8244
timestamp 1677677812
transform 1 0 2424 0 1 1370
box -8 -3 16 105
use FILL  FILL_8245
timestamp 1677677812
transform 1 0 2432 0 1 1370
box -8 -3 16 105
use FAX1  FAX1_4
timestamp 1677677812
transform -1 0 2560 0 1 1370
box -5 -3 126 105
use FILL  FILL_8246
timestamp 1677677812
transform 1 0 2560 0 1 1370
box -8 -3 16 105
use FILL  FILL_8247
timestamp 1677677812
transform 1 0 2568 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6283
timestamp 1677677812
transform 1 0 2652 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6284
timestamp 1677677812
transform 1 0 2676 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_447
timestamp 1677677812
transform -1 0 2672 0 1 1370
box -8 -3 104 105
use FILL  FILL_8248
timestamp 1677677812
transform 1 0 2672 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6285
timestamp 1677677812
transform 1 0 2732 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6286
timestamp 1677677812
transform 1 0 2756 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_448
timestamp 1677677812
transform -1 0 2776 0 1 1370
box -8 -3 104 105
use FILL  FILL_8249
timestamp 1677677812
transform 1 0 2776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8265
timestamp 1677677812
transform 1 0 2784 0 1 1370
box -8 -3 16 105
use FAX1  FAX1_6
timestamp 1677677812
transform 1 0 2792 0 1 1370
box -5 -3 126 105
use FILL  FILL_8266
timestamp 1677677812
transform 1 0 2912 0 1 1370
box -8 -3 16 105
use FILL  FILL_8267
timestamp 1677677812
transform 1 0 2920 0 1 1370
box -8 -3 16 105
use FILL  FILL_8268
timestamp 1677677812
transform 1 0 2928 0 1 1370
box -8 -3 16 105
use FILL  FILL_8270
timestamp 1677677812
transform 1 0 2936 0 1 1370
box -8 -3 16 105
use FILL  FILL_8272
timestamp 1677677812
transform 1 0 2944 0 1 1370
box -8 -3 16 105
use FILL  FILL_8274
timestamp 1677677812
transform 1 0 2952 0 1 1370
box -8 -3 16 105
use FILL  FILL_8276
timestamp 1677677812
transform 1 0 2960 0 1 1370
box -8 -3 16 105
use FILL  FILL_8278
timestamp 1677677812
transform 1 0 2968 0 1 1370
box -8 -3 16 105
use FILL  FILL_8279
timestamp 1677677812
transform 1 0 2976 0 1 1370
box -8 -3 16 105
use FILL  FILL_8280
timestamp 1677677812
transform 1 0 2984 0 1 1370
box -8 -3 16 105
use FILL  FILL_8281
timestamp 1677677812
transform 1 0 2992 0 1 1370
box -8 -3 16 105
use FILL  FILL_8282
timestamp 1677677812
transform 1 0 3000 0 1 1370
box -8 -3 16 105
use FILL  FILL_8284
timestamp 1677677812
transform 1 0 3008 0 1 1370
box -8 -3 16 105
use FILL  FILL_8285
timestamp 1677677812
transform 1 0 3016 0 1 1370
box -8 -3 16 105
use FILL  FILL_8286
timestamp 1677677812
transform 1 0 3024 0 1 1370
box -8 -3 16 105
use FILL  FILL_8287
timestamp 1677677812
transform 1 0 3032 0 1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_64
timestamp 1677677812
transform -1 0 3072 0 1 1370
box -8 -3 40 105
use FILL  FILL_8288
timestamp 1677677812
transform 1 0 3072 0 1 1370
box -8 -3 16 105
use FILL  FILL_8291
timestamp 1677677812
transform 1 0 3080 0 1 1370
box -8 -3 16 105
use FILL  FILL_8293
timestamp 1677677812
transform 1 0 3088 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_520
timestamp 1677677812
transform 1 0 3096 0 1 1370
box -9 -3 26 105
use FILL  FILL_8295
timestamp 1677677812
transform 1 0 3112 0 1 1370
box -8 -3 16 105
use FILL  FILL_8296
timestamp 1677677812
transform 1 0 3120 0 1 1370
box -8 -3 16 105
use FILL  FILL_8299
timestamp 1677677812
transform 1 0 3128 0 1 1370
box -8 -3 16 105
use FILL  FILL_8300
timestamp 1677677812
transform 1 0 3136 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_141
timestamp 1677677812
transform -1 0 3176 0 1 1370
box -8 -3 34 105
use FILL  FILL_8301
timestamp 1677677812
transform 1 0 3176 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6287
timestamp 1677677812
transform 1 0 3196 0 1 1375
box -3 -3 3 3
use FILL  FILL_8302
timestamp 1677677812
transform 1 0 3184 0 1 1370
box -8 -3 16 105
use FILL  FILL_8303
timestamp 1677677812
transform 1 0 3192 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6288
timestamp 1677677812
transform 1 0 3228 0 1 1375
box -3 -3 3 3
use AOI22X1  AOI22X1_309
timestamp 1677677812
transform 1 0 3200 0 1 1370
box -8 -3 46 105
use FILL  FILL_8304
timestamp 1677677812
transform 1 0 3240 0 1 1370
box -8 -3 16 105
use FILL  FILL_8305
timestamp 1677677812
transform 1 0 3248 0 1 1370
box -8 -3 16 105
use FILL  FILL_8306
timestamp 1677677812
transform 1 0 3256 0 1 1370
box -8 -3 16 105
use FILL  FILL_8307
timestamp 1677677812
transform 1 0 3264 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6289
timestamp 1677677812
transform 1 0 3284 0 1 1375
box -3 -3 3 3
use FILL  FILL_8313
timestamp 1677677812
transform 1 0 3272 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_7
timestamp 1677677812
transform 1 0 3280 0 1 1370
box -7 -3 39 105
use FILL  FILL_8315
timestamp 1677677812
transform 1 0 3312 0 1 1370
box -8 -3 16 105
use FILL  FILL_8316
timestamp 1677677812
transform 1 0 3320 0 1 1370
box -8 -3 16 105
use FILL  FILL_8317
timestamp 1677677812
transform 1 0 3328 0 1 1370
box -8 -3 16 105
use FILL  FILL_8321
timestamp 1677677812
transform 1 0 3336 0 1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_8
timestamp 1677677812
transform -1 0 3376 0 1 1370
box -7 -3 39 105
use FILL  FILL_8322
timestamp 1677677812
transform 1 0 3376 0 1 1370
box -8 -3 16 105
use FILL  FILL_8323
timestamp 1677677812
transform 1 0 3384 0 1 1370
box -8 -3 16 105
use FILL  FILL_8324
timestamp 1677677812
transform 1 0 3392 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6290
timestamp 1677677812
transform 1 0 3484 0 1 1375
box -3 -3 3 3
use FAX1  FAX1_8
timestamp 1677677812
transform 1 0 3400 0 1 1370
box -5 -3 126 105
use BUFX2  BUFX2_103
timestamp 1677677812
transform 1 0 3520 0 1 1370
box -5 -3 28 105
use M3_M2  M3_M2_6291
timestamp 1677677812
transform 1 0 3668 0 1 1375
box -3 -3 3 3
use FAX1  FAX1_9
timestamp 1677677812
transform 1 0 3544 0 1 1370
box -5 -3 126 105
use FILL  FILL_8325
timestamp 1677677812
transform 1 0 3664 0 1 1370
box -8 -3 16 105
use FILL  FILL_8339
timestamp 1677677812
transform 1 0 3672 0 1 1370
box -8 -3 16 105
use FILL  FILL_8340
timestamp 1677677812
transform 1 0 3680 0 1 1370
box -8 -3 16 105
use FILL  FILL_8341
timestamp 1677677812
transform 1 0 3688 0 1 1370
box -8 -3 16 105
use FILL  FILL_8342
timestamp 1677677812
transform 1 0 3696 0 1 1370
box -8 -3 16 105
use FILL  FILL_8343
timestamp 1677677812
transform 1 0 3704 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_13
timestamp 1677677812
transform -1 0 3736 0 1 1370
box -8 -3 32 105
use FILL  FILL_8344
timestamp 1677677812
transform 1 0 3736 0 1 1370
box -8 -3 16 105
use FILL  FILL_8349
timestamp 1677677812
transform 1 0 3744 0 1 1370
box -8 -3 16 105
use FILL  FILL_8351
timestamp 1677677812
transform 1 0 3752 0 1 1370
box -8 -3 16 105
use FILL  FILL_8353
timestamp 1677677812
transform 1 0 3760 0 1 1370
box -8 -3 16 105
use FILL  FILL_8354
timestamp 1677677812
transform 1 0 3768 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_143
timestamp 1677677812
transform 1 0 3776 0 1 1370
box -8 -3 34 105
use FILL  FILL_8355
timestamp 1677677812
transform 1 0 3808 0 1 1370
box -8 -3 16 105
use FILL  FILL_8358
timestamp 1677677812
transform 1 0 3816 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_14
timestamp 1677677812
transform -1 0 3848 0 1 1370
box -8 -3 32 105
use FILL  FILL_8359
timestamp 1677677812
transform 1 0 3848 0 1 1370
box -8 -3 16 105
use FILL  FILL_8360
timestamp 1677677812
transform 1 0 3856 0 1 1370
box -8 -3 16 105
use FILL  FILL_8361
timestamp 1677677812
transform 1 0 3864 0 1 1370
box -8 -3 16 105
use BUFX2  BUFX2_104
timestamp 1677677812
transform 1 0 3872 0 1 1370
box -5 -3 28 105
use FILL  FILL_8362
timestamp 1677677812
transform 1 0 3896 0 1 1370
box -8 -3 16 105
use FILL  FILL_8363
timestamp 1677677812
transform 1 0 3904 0 1 1370
box -8 -3 16 105
use FILL  FILL_8364
timestamp 1677677812
transform 1 0 3912 0 1 1370
box -8 -3 16 105
use FILL  FILL_8365
timestamp 1677677812
transform 1 0 3920 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_144
timestamp 1677677812
transform 1 0 3928 0 1 1370
box -8 -3 34 105
use FILL  FILL_8366
timestamp 1677677812
transform 1 0 3960 0 1 1370
box -8 -3 16 105
use FILL  FILL_8367
timestamp 1677677812
transform 1 0 3968 0 1 1370
box -8 -3 16 105
use FILL  FILL_8368
timestamp 1677677812
transform 1 0 3976 0 1 1370
box -8 -3 16 105
use FILL  FILL_8369
timestamp 1677677812
transform 1 0 3984 0 1 1370
box -8 -3 16 105
use FILL  FILL_8370
timestamp 1677677812
transform 1 0 3992 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1677677812
transform 1 0 4000 0 1 1370
box -8 -3 32 105
use FILL  FILL_8371
timestamp 1677677812
transform 1 0 4024 0 1 1370
box -8 -3 16 105
use FILL  FILL_8375
timestamp 1677677812
transform 1 0 4032 0 1 1370
box -8 -3 16 105
use FILL  FILL_8377
timestamp 1677677812
transform 1 0 4040 0 1 1370
box -8 -3 16 105
use FILL  FILL_8378
timestamp 1677677812
transform 1 0 4048 0 1 1370
box -8 -3 16 105
use FILL  FILL_8379
timestamp 1677677812
transform 1 0 4056 0 1 1370
box -8 -3 16 105
use FILL  FILL_8380
timestamp 1677677812
transform 1 0 4064 0 1 1370
box -8 -3 16 105
use FILL  FILL_8381
timestamp 1677677812
transform 1 0 4072 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6292
timestamp 1677677812
transform 1 0 4108 0 1 1375
box -3 -3 3 3
use NAND2X1  NAND2X1_16
timestamp 1677677812
transform -1 0 4104 0 1 1370
box -8 -3 32 105
use FILL  FILL_8382
timestamp 1677677812
transform 1 0 4104 0 1 1370
box -8 -3 16 105
use FILL  FILL_8383
timestamp 1677677812
transform 1 0 4112 0 1 1370
box -8 -3 16 105
use FILL  FILL_8384
timestamp 1677677812
transform 1 0 4120 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6293
timestamp 1677677812
transform 1 0 4140 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_453
timestamp 1677677812
transform 1 0 4128 0 1 1370
box -8 -3 104 105
use OAI21X1  OAI21X1_145
timestamp 1677677812
transform 1 0 4224 0 1 1370
box -8 -3 34 105
use FILL  FILL_8385
timestamp 1677677812
transform 1 0 4256 0 1 1370
box -8 -3 16 105
use FILL  FILL_8401
timestamp 1677677812
transform 1 0 4264 0 1 1370
box -8 -3 16 105
use FILL  FILL_8402
timestamp 1677677812
transform 1 0 4272 0 1 1370
box -8 -3 16 105
use FILL  FILL_8403
timestamp 1677677812
transform 1 0 4280 0 1 1370
box -8 -3 16 105
use FILL  FILL_8404
timestamp 1677677812
transform 1 0 4288 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_527
timestamp 1677677812
transform -1 0 4312 0 1 1370
box -9 -3 26 105
use FILL  FILL_8405
timestamp 1677677812
transform 1 0 4312 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6294
timestamp 1677677812
transform 1 0 4348 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_6295
timestamp 1677677812
transform 1 0 4404 0 1 1375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_454
timestamp 1677677812
transform -1 0 4416 0 1 1370
box -8 -3 104 105
use FILL  FILL_8406
timestamp 1677677812
transform 1 0 4416 0 1 1370
box -8 -3 16 105
use FILL  FILL_8407
timestamp 1677677812
transform 1 0 4424 0 1 1370
box -8 -3 16 105
use FILL  FILL_8408
timestamp 1677677812
transform 1 0 4432 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_147
timestamp 1677677812
transform -1 0 4472 0 1 1370
box -8 -3 34 105
use FILL  FILL_8409
timestamp 1677677812
transform 1 0 4472 0 1 1370
box -8 -3 16 105
use FILL  FILL_8410
timestamp 1677677812
transform 1 0 4480 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6296
timestamp 1677677812
transform 1 0 4500 0 1 1375
box -3 -3 3 3
use FILL  FILL_8418
timestamp 1677677812
transform 1 0 4488 0 1 1370
box -8 -3 16 105
use FILL  FILL_8419
timestamp 1677677812
transform 1 0 4496 0 1 1370
box -8 -3 16 105
use FILL  FILL_8420
timestamp 1677677812
transform 1 0 4504 0 1 1370
box -8 -3 16 105
use FILL  FILL_8421
timestamp 1677677812
transform 1 0 4512 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_149
timestamp 1677677812
transform -1 0 4552 0 1 1370
box -8 -3 34 105
use FILL  FILL_8422
timestamp 1677677812
transform 1 0 4552 0 1 1370
box -8 -3 16 105
use FILL  FILL_8423
timestamp 1677677812
transform 1 0 4560 0 1 1370
box -8 -3 16 105
use FILL  FILL_8424
timestamp 1677677812
transform 1 0 4568 0 1 1370
box -8 -3 16 105
use FILL  FILL_8425
timestamp 1677677812
transform 1 0 4576 0 1 1370
box -8 -3 16 105
use FILL  FILL_8426
timestamp 1677677812
transform 1 0 4584 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_150
timestamp 1677677812
transform -1 0 4624 0 1 1370
box -8 -3 34 105
use FILL  FILL_8427
timestamp 1677677812
transform 1 0 4624 0 1 1370
box -8 -3 16 105
use FILL  FILL_8432
timestamp 1677677812
transform 1 0 4632 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_529
timestamp 1677677812
transform 1 0 4640 0 1 1370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_457
timestamp 1677677812
transform 1 0 4656 0 1 1370
box -8 -3 104 105
use INVX2  INVX2_530
timestamp 1677677812
transform -1 0 4768 0 1 1370
box -9 -3 26 105
use FILL  FILL_8434
timestamp 1677677812
transform 1 0 4768 0 1 1370
box -8 -3 16 105
use FILL  FILL_8435
timestamp 1677677812
transform 1 0 4776 0 1 1370
box -8 -3 16 105
use FILL  FILL_8444
timestamp 1677677812
transform 1 0 4784 0 1 1370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_67
timestamp 1677677812
transform 1 0 4819 0 1 1370
box -10 -3 10 3
use M2_M1  M2_M1_7048
timestamp 1677677812
transform 1 0 92 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6379
timestamp 1677677812
transform 1 0 172 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7138
timestamp 1677677812
transform 1 0 140 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7139
timestamp 1677677812
transform 1 0 172 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7140
timestamp 1677677812
transform 1 0 180 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6411
timestamp 1677677812
transform 1 0 140 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6412
timestamp 1677677812
transform 1 0 180 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6297
timestamp 1677677812
transform 1 0 228 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6298
timestamp 1677677812
transform 1 0 260 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6450
timestamp 1677677812
transform 1 0 268 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7039
timestamp 1677677812
transform 1 0 284 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6380
timestamp 1677677812
transform 1 0 292 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6319
timestamp 1677677812
transform 1 0 324 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7049
timestamp 1677677812
transform 1 0 308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7050
timestamp 1677677812
transform 1 0 324 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6381
timestamp 1677677812
transform 1 0 332 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7051
timestamp 1677677812
transform 1 0 340 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7052
timestamp 1677677812
transform 1 0 356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7141
timestamp 1677677812
transform 1 0 316 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7142
timestamp 1677677812
transform 1 0 340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7143
timestamp 1677677812
transform 1 0 380 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7144
timestamp 1677677812
transform 1 0 436 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6413
timestamp 1677677812
transform 1 0 340 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6414
timestamp 1677677812
transform 1 0 444 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6299
timestamp 1677677812
transform 1 0 516 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7053
timestamp 1677677812
transform 1 0 460 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7145
timestamp 1677677812
transform 1 0 508 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6300
timestamp 1677677812
transform 1 0 572 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6344
timestamp 1677677812
transform 1 0 556 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6345
timestamp 1677677812
transform 1 0 580 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7054
timestamp 1677677812
transform 1 0 556 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7055
timestamp 1677677812
transform 1 0 580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7146
timestamp 1677677812
transform 1 0 548 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7147
timestamp 1677677812
transform 1 0 556 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7148
timestamp 1677677812
transform 1 0 572 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6415
timestamp 1677677812
transform 1 0 548 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6416
timestamp 1677677812
transform 1 0 580 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6451
timestamp 1677677812
transform 1 0 556 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6346
timestamp 1677677812
transform 1 0 604 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7149
timestamp 1677677812
transform 1 0 612 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7150
timestamp 1677677812
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6417
timestamp 1677677812
transform 1 0 612 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7056
timestamp 1677677812
transform 1 0 644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7151
timestamp 1677677812
transform 1 0 652 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6418
timestamp 1677677812
transform 1 0 628 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6419
timestamp 1677677812
transform 1 0 644 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6452
timestamp 1677677812
transform 1 0 636 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6479
timestamp 1677677812
transform 1 0 652 0 1 1285
box -3 -3 3 3
use M2_M1  M2_M1_7057
timestamp 1677677812
transform 1 0 668 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6347
timestamp 1677677812
transform 1 0 676 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6382
timestamp 1677677812
transform 1 0 676 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7152
timestamp 1677677812
transform 1 0 676 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6301
timestamp 1677677812
transform 1 0 756 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6348
timestamp 1677677812
transform 1 0 692 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6349
timestamp 1677677812
transform 1 0 764 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6383
timestamp 1677677812
transform 1 0 700 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7058
timestamp 1677677812
transform 1 0 764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7153
timestamp 1677677812
transform 1 0 740 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6453
timestamp 1677677812
transform 1 0 692 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6480
timestamp 1677677812
transform 1 0 740 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6320
timestamp 1677677812
transform 1 0 780 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7040
timestamp 1677677812
transform 1 0 780 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6474
timestamp 1677677812
transform 1 0 780 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6481
timestamp 1677677812
transform 1 0 780 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6302
timestamp 1677677812
transform 1 0 796 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6350
timestamp 1677677812
transform 1 0 804 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7059
timestamp 1677677812
transform 1 0 884 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7154
timestamp 1677677812
transform 1 0 1020 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7155
timestamp 1677677812
transform 1 0 1028 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6475
timestamp 1677677812
transform 1 0 1020 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7041
timestamp 1677677812
transform 1 0 1052 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6351
timestamp 1677677812
transform 1 0 1164 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7060
timestamp 1677677812
transform 1 0 1180 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6420
timestamp 1677677812
transform 1 0 1188 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6321
timestamp 1677677812
transform 1 0 1204 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6303
timestamp 1677677812
transform 1 0 1220 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6304
timestamp 1677677812
transform 1 0 1268 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6322
timestamp 1677677812
transform 1 0 1244 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6323
timestamp 1677677812
transform 1 0 1268 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6352
timestamp 1677677812
transform 1 0 1236 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7061
timestamp 1677677812
transform 1 0 1228 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7062
timestamp 1677677812
transform 1 0 1236 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6353
timestamp 1677677812
transform 1 0 1260 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6384
timestamp 1677677812
transform 1 0 1284 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6324
timestamp 1677677812
transform 1 0 1308 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6354
timestamp 1677677812
transform 1 0 1300 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7063
timestamp 1677677812
transform 1 0 1292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7156
timestamp 1677677812
transform 1 0 1236 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7157
timestamp 1677677812
transform 1 0 1244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7158
timestamp 1677677812
transform 1 0 1260 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7159
timestamp 1677677812
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6482
timestamp 1677677812
transform 1 0 1244 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6421
timestamp 1677677812
transform 1 0 1276 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6422
timestamp 1677677812
transform 1 0 1292 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6355
timestamp 1677677812
transform 1 0 1316 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7064
timestamp 1677677812
transform 1 0 1316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7160
timestamp 1677677812
transform 1 0 1340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7161
timestamp 1677677812
transform 1 0 1396 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6423
timestamp 1677677812
transform 1 0 1396 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6325
timestamp 1677677812
transform 1 0 1468 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6385
timestamp 1677677812
transform 1 0 1444 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7065
timestamp 1677677812
transform 1 0 1452 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7162
timestamp 1677677812
transform 1 0 1444 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7163
timestamp 1677677812
transform 1 0 1468 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6424
timestamp 1677677812
transform 1 0 1468 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7237
timestamp 1677677812
transform 1 0 1476 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6483
timestamp 1677677812
transform 1 0 1460 0 1 1285
box -3 -3 3 3
use M3_M2  M3_M2_6326
timestamp 1677677812
transform 1 0 1540 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6356
timestamp 1677677812
transform 1 0 1500 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6386
timestamp 1677677812
transform 1 0 1556 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7066
timestamp 1677677812
transform 1 0 1580 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7164
timestamp 1677677812
transform 1 0 1532 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6476
timestamp 1677677812
transform 1 0 1564 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6357
timestamp 1677677812
transform 1 0 1596 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7067
timestamp 1677677812
transform 1 0 1596 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6425
timestamp 1677677812
transform 1 0 1596 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7165
timestamp 1677677812
transform 1 0 1628 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7166
timestamp 1677677812
transform 1 0 1636 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6426
timestamp 1677677812
transform 1 0 1636 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6327
timestamp 1677677812
transform 1 0 1684 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7068
timestamp 1677677812
transform 1 0 1652 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6387
timestamp 1677677812
transform 1 0 1660 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7069
timestamp 1677677812
transform 1 0 1668 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6388
timestamp 1677677812
transform 1 0 1676 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6394
timestamp 1677677812
transform 1 0 1652 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7167
timestamp 1677677812
transform 1 0 1676 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7168
timestamp 1677677812
transform 1 0 1692 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6358
timestamp 1677677812
transform 1 0 1724 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6359
timestamp 1677677812
transform 1 0 1748 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7070
timestamp 1677677812
transform 1 0 1724 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7071
timestamp 1677677812
transform 1 0 1732 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7072
timestamp 1677677812
transform 1 0 1748 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7169
timestamp 1677677812
transform 1 0 1724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7170
timestamp 1677677812
transform 1 0 1740 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7171
timestamp 1677677812
transform 1 0 1756 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6427
timestamp 1677677812
transform 1 0 1740 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6454
timestamp 1677677812
transform 1 0 1724 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6428
timestamp 1677677812
transform 1 0 1764 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6429
timestamp 1677677812
transform 1 0 1780 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6328
timestamp 1677677812
transform 1 0 1868 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7073
timestamp 1677677812
transform 1 0 1868 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7172
timestamp 1677677812
transform 1 0 1820 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6430
timestamp 1677677812
transform 1 0 1820 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6329
timestamp 1677677812
transform 1 0 1892 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6395
timestamp 1677677812
transform 1 0 1884 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7173
timestamp 1677677812
transform 1 0 1940 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7174
timestamp 1677677812
transform 1 0 1964 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7074
timestamp 1677677812
transform 1 0 1996 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7075
timestamp 1677677812
transform 1 0 2004 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7076
timestamp 1677677812
transform 1 0 2020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7175
timestamp 1677677812
transform 1 0 1996 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6396
timestamp 1677677812
transform 1 0 2004 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7176
timestamp 1677677812
transform 1 0 2012 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7177
timestamp 1677677812
transform 1 0 2028 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7178
timestamp 1677677812
transform 1 0 2036 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6455
timestamp 1677677812
transform 1 0 2028 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7077
timestamp 1677677812
transform 1 0 2132 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7179
timestamp 1677677812
transform 1 0 2084 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7238
timestamp 1677677812
transform 1 0 2148 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6360
timestamp 1677677812
transform 1 0 2188 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6389
timestamp 1677677812
transform 1 0 2180 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7078
timestamp 1677677812
transform 1 0 2292 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7079
timestamp 1677677812
transform 1 0 2308 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7180
timestamp 1677677812
transform 1 0 2180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7181
timestamp 1677677812
transform 1 0 2196 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7182
timestamp 1677677812
transform 1 0 2204 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7183
timestamp 1677677812
transform 1 0 2212 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7184
timestamp 1677677812
transform 1 0 2252 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7239
timestamp 1677677812
transform 1 0 2188 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6431
timestamp 1677677812
transform 1 0 2196 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6432
timestamp 1677677812
transform 1 0 2212 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7247
timestamp 1677677812
transform 1 0 2172 0 1 1305
box -2 -2 2 2
use M2_M1  M2_M1_7240
timestamp 1677677812
transform 1 0 2316 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7185
timestamp 1677677812
transform 1 0 2340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7080
timestamp 1677677812
transform 1 0 2356 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7241
timestamp 1677677812
transform 1 0 2348 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6456
timestamp 1677677812
transform 1 0 2356 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6305
timestamp 1677677812
transform 1 0 2380 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7186
timestamp 1677677812
transform 1 0 2372 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6330
timestamp 1677677812
transform 1 0 2396 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6331
timestamp 1677677812
transform 1 0 2420 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6361
timestamp 1677677812
transform 1 0 2404 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7042
timestamp 1677677812
transform 1 0 2412 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7081
timestamp 1677677812
transform 1 0 2396 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7082
timestamp 1677677812
transform 1 0 2404 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6397
timestamp 1677677812
transform 1 0 2468 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7187
timestamp 1677677812
transform 1 0 2500 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6457
timestamp 1677677812
transform 1 0 2436 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6458
timestamp 1677677812
transform 1 0 2460 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6332
timestamp 1677677812
transform 1 0 2532 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6306
timestamp 1677677812
transform 1 0 2548 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6362
timestamp 1677677812
transform 1 0 2540 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7083
timestamp 1677677812
transform 1 0 2532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7188
timestamp 1677677812
transform 1 0 2524 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7084
timestamp 1677677812
transform 1 0 2588 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7189
timestamp 1677677812
transform 1 0 2564 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6477
timestamp 1677677812
transform 1 0 2588 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_7085
timestamp 1677677812
transform 1 0 2604 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6333
timestamp 1677677812
transform 1 0 2620 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6307
timestamp 1677677812
transform 1 0 2676 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6334
timestamp 1677677812
transform 1 0 2660 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7086
timestamp 1677677812
transform 1 0 2644 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7087
timestamp 1677677812
transform 1 0 2660 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6308
timestamp 1677677812
transform 1 0 2716 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7088
timestamp 1677677812
transform 1 0 2692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7190
timestamp 1677677812
transform 1 0 2620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7191
timestamp 1677677812
transform 1 0 2636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7192
timestamp 1677677812
transform 1 0 2652 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7193
timestamp 1677677812
transform 1 0 2668 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7194
timestamp 1677677812
transform 1 0 2684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7195
timestamp 1677677812
transform 1 0 2692 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6433
timestamp 1677677812
transform 1 0 2620 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6434
timestamp 1677677812
transform 1 0 2692 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6478
timestamp 1677677812
transform 1 0 2668 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_6335
timestamp 1677677812
transform 1 0 2748 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7089
timestamp 1677677812
transform 1 0 2740 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7090
timestamp 1677677812
transform 1 0 2748 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6459
timestamp 1677677812
transform 1 0 2700 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6460
timestamp 1677677812
transform 1 0 2756 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6309
timestamp 1677677812
transform 1 0 2812 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6310
timestamp 1677677812
transform 1 0 2908 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6336
timestamp 1677677812
transform 1 0 2892 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7043
timestamp 1677677812
transform 1 0 2892 0 1 1345
box -2 -2 2 2
use M3_M2  M3_M2_6363
timestamp 1677677812
transform 1 0 2900 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7091
timestamp 1677677812
transform 1 0 2900 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7196
timestamp 1677677812
transform 1 0 2796 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7197
timestamp 1677677812
transform 1 0 2804 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7198
timestamp 1677677812
transform 1 0 2908 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6461
timestamp 1677677812
transform 1 0 2796 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6462
timestamp 1677677812
transform 1 0 2844 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6364
timestamp 1677677812
transform 1 0 2932 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7199
timestamp 1677677812
transform 1 0 2932 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7092
timestamp 1677677812
transform 1 0 2964 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6365
timestamp 1677677812
transform 1 0 2980 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6337
timestamp 1677677812
transform 1 0 3004 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7044
timestamp 1677677812
transform 1 0 2996 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7093
timestamp 1677677812
transform 1 0 2980 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6366
timestamp 1677677812
transform 1 0 3020 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7045
timestamp 1677677812
transform 1 0 3044 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7094
timestamp 1677677812
transform 1 0 3012 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7095
timestamp 1677677812
transform 1 0 3020 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7096
timestamp 1677677812
transform 1 0 3036 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7200
timestamp 1677677812
transform 1 0 3004 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6367
timestamp 1677677812
transform 1 0 3052 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7201
timestamp 1677677812
transform 1 0 3052 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7202
timestamp 1677677812
transform 1 0 3060 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7242
timestamp 1677677812
transform 1 0 3068 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7097
timestamp 1677677812
transform 1 0 3100 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6398
timestamp 1677677812
transform 1 0 3100 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6368
timestamp 1677677812
transform 1 0 3124 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7098
timestamp 1677677812
transform 1 0 3124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7203
timestamp 1677677812
transform 1 0 3124 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6435
timestamp 1677677812
transform 1 0 3124 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7243
timestamp 1677677812
transform 1 0 3140 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6338
timestamp 1677677812
transform 1 0 3180 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6339
timestamp 1677677812
transform 1 0 3204 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6369
timestamp 1677677812
transform 1 0 3172 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7099
timestamp 1677677812
transform 1 0 3172 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7100
timestamp 1677677812
transform 1 0 3180 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7101
timestamp 1677677812
transform 1 0 3196 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7102
timestamp 1677677812
transform 1 0 3204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7204
timestamp 1677677812
transform 1 0 3164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7205
timestamp 1677677812
transform 1 0 3172 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7206
timestamp 1677677812
transform 1 0 3188 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6436
timestamp 1677677812
transform 1 0 3164 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6437
timestamp 1677677812
transform 1 0 3180 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6463
timestamp 1677677812
transform 1 0 3172 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6464
timestamp 1677677812
transform 1 0 3212 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6311
timestamp 1677677812
transform 1 0 3228 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7207
timestamp 1677677812
transform 1 0 3228 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7208
timestamp 1677677812
transform 1 0 3244 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6370
timestamp 1677677812
transform 1 0 3268 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7103
timestamp 1677677812
transform 1 0 3260 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6438
timestamp 1677677812
transform 1 0 3244 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6439
timestamp 1677677812
transform 1 0 3260 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7104
timestamp 1677677812
transform 1 0 3300 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7244
timestamp 1677677812
transform 1 0 3308 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7248
timestamp 1677677812
transform 1 0 3324 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_6312
timestamp 1677677812
transform 1 0 3388 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6340
timestamp 1677677812
transform 1 0 3380 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6341
timestamp 1677677812
transform 1 0 3420 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6342
timestamp 1677677812
transform 1 0 3492 0 1 1355
box -3 -3 3 3
use M2_M1  M2_M1_7046
timestamp 1677677812
transform 1 0 3388 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7105
timestamp 1677677812
transform 1 0 3380 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7106
timestamp 1677677812
transform 1 0 3492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7209
timestamp 1677677812
transform 1 0 3476 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7210
timestamp 1677677812
transform 1 0 3484 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6399
timestamp 1677677812
transform 1 0 3492 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6313
timestamp 1677677812
transform 1 0 3548 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6371
timestamp 1677677812
transform 1 0 3524 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6372
timestamp 1677677812
transform 1 0 3540 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7107
timestamp 1677677812
transform 1 0 3524 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7211
timestamp 1677677812
transform 1 0 3572 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6440
timestamp 1677677812
transform 1 0 3572 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7108
timestamp 1677677812
transform 1 0 3652 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6314
timestamp 1677677812
transform 1 0 3692 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7109
timestamp 1677677812
transform 1 0 3692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7110
timestamp 1677677812
transform 1 0 3708 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7212
timestamp 1677677812
transform 1 0 3684 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7213
timestamp 1677677812
transform 1 0 3700 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6441
timestamp 1677677812
transform 1 0 3692 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6465
timestamp 1677677812
transform 1 0 3700 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7111
timestamp 1677677812
transform 1 0 3764 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7112
timestamp 1677677812
transform 1 0 3780 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6390
timestamp 1677677812
transform 1 0 3788 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7214
timestamp 1677677812
transform 1 0 3772 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7215
timestamp 1677677812
transform 1 0 3788 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6466
timestamp 1677677812
transform 1 0 3788 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7113
timestamp 1677677812
transform 1 0 3820 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6315
timestamp 1677677812
transform 1 0 3868 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6343
timestamp 1677677812
transform 1 0 3836 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_6373
timestamp 1677677812
transform 1 0 3876 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6374
timestamp 1677677812
transform 1 0 3908 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_6391
timestamp 1677677812
transform 1 0 3860 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7114
timestamp 1677677812
transform 1 0 3908 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7216
timestamp 1677677812
transform 1 0 3828 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7217
timestamp 1677677812
transform 1 0 3860 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6442
timestamp 1677677812
transform 1 0 3820 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6400
timestamp 1677677812
transform 1 0 3884 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6401
timestamp 1677677812
transform 1 0 3908 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6443
timestamp 1677677812
transform 1 0 3860 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7115
timestamp 1677677812
transform 1 0 3932 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7218
timestamp 1677677812
transform 1 0 3980 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6467
timestamp 1677677812
transform 1 0 3916 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6468
timestamp 1677677812
transform 1 0 3996 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7116
timestamp 1677677812
transform 1 0 4028 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7117
timestamp 1677677812
transform 1 0 4068 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7219
timestamp 1677677812
transform 1 0 4044 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7220
timestamp 1677677812
transform 1 0 4052 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6469
timestamp 1677677812
transform 1 0 4044 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7118
timestamp 1677677812
transform 1 0 4084 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7119
timestamp 1677677812
transform 1 0 4092 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6402
timestamp 1677677812
transform 1 0 4076 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6470
timestamp 1677677812
transform 1 0 4068 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7245
timestamp 1677677812
transform 1 0 4076 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_7120
timestamp 1677677812
transform 1 0 4124 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7121
timestamp 1677677812
transform 1 0 4140 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7221
timestamp 1677677812
transform 1 0 4116 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6403
timestamp 1677677812
transform 1 0 4124 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7222
timestamp 1677677812
transform 1 0 4132 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6444
timestamp 1677677812
transform 1 0 4116 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6471
timestamp 1677677812
transform 1 0 4132 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7223
timestamp 1677677812
transform 1 0 4148 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6445
timestamp 1677677812
transform 1 0 4148 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6404
timestamp 1677677812
transform 1 0 4172 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7224
timestamp 1677677812
transform 1 0 4180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7047
timestamp 1677677812
transform 1 0 4220 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_7122
timestamp 1677677812
transform 1 0 4260 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7123
timestamp 1677677812
transform 1 0 4268 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7124
timestamp 1677677812
transform 1 0 4284 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7225
timestamp 1677677812
transform 1 0 4252 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6405
timestamp 1677677812
transform 1 0 4260 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7226
timestamp 1677677812
transform 1 0 4276 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7227
timestamp 1677677812
transform 1 0 4292 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6446
timestamp 1677677812
transform 1 0 4268 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6447
timestamp 1677677812
transform 1 0 4284 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_6472
timestamp 1677677812
transform 1 0 4268 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_6473
timestamp 1677677812
transform 1 0 4292 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_7125
timestamp 1677677812
transform 1 0 4332 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6375
timestamp 1677677812
transform 1 0 4396 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7126
timestamp 1677677812
transform 1 0 4348 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6316
timestamp 1677677812
transform 1 0 4436 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7127
timestamp 1677677812
transform 1 0 4436 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7228
timestamp 1677677812
transform 1 0 4372 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7229
timestamp 1677677812
transform 1 0 4428 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6406
timestamp 1677677812
transform 1 0 4436 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7246
timestamp 1677677812
transform 1 0 4436 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_6317
timestamp 1677677812
transform 1 0 4460 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_6376
timestamp 1677677812
transform 1 0 4476 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7128
timestamp 1677677812
transform 1 0 4476 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6392
timestamp 1677677812
transform 1 0 4484 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_7230
timestamp 1677677812
transform 1 0 4484 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6318
timestamp 1677677812
transform 1 0 4508 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_7129
timestamp 1677677812
transform 1 0 4500 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6393
timestamp 1677677812
transform 1 0 4564 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_6407
timestamp 1677677812
transform 1 0 4500 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6408
timestamp 1677677812
transform 1 0 4524 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7231
timestamp 1677677812
transform 1 0 4532 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6409
timestamp 1677677812
transform 1 0 4540 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_6410
timestamp 1677677812
transform 1 0 4564 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_7232
timestamp 1677677812
transform 1 0 4620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7130
timestamp 1677677812
transform 1 0 4636 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6377
timestamp 1677677812
transform 1 0 4660 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7131
timestamp 1677677812
transform 1 0 4668 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7132
timestamp 1677677812
transform 1 0 4684 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7133
timestamp 1677677812
transform 1 0 4692 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7233
timestamp 1677677812
transform 1 0 4660 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7234
timestamp 1677677812
transform 1 0 4676 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6448
timestamp 1677677812
transform 1 0 4676 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7134
timestamp 1677677812
transform 1 0 4732 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_6378
timestamp 1677677812
transform 1 0 4772 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_7135
timestamp 1677677812
transform 1 0 4756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7136
timestamp 1677677812
transform 1 0 4772 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_7235
timestamp 1677677812
transform 1 0 4748 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_7236
timestamp 1677677812
transform 1 0 4764 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_6449
timestamp 1677677812
transform 1 0 4740 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_7137
timestamp 1677677812
transform 1 0 4788 0 1 1335
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_68
timestamp 1677677812
transform 1 0 24 0 1 1270
box -10 -3 10 3
use FILL  FILL_8012
timestamp 1677677812
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_433
timestamp 1677677812
transform 1 0 80 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8013
timestamp 1677677812
transform 1 0 176 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8014
timestamp 1677677812
transform 1 0 184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8015
timestamp 1677677812
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8016
timestamp 1677677812
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8017
timestamp 1677677812
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8018
timestamp 1677677812
transform 1 0 216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8019
timestamp 1677677812
transform 1 0 224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8020
timestamp 1677677812
transform 1 0 232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8049
timestamp 1677677812
transform 1 0 240 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_512
timestamp 1677677812
transform -1 0 264 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8050
timestamp 1677677812
transform 1 0 264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8051
timestamp 1677677812
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8052
timestamp 1677677812
transform 1 0 280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8053
timestamp 1677677812
transform 1 0 288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8054
timestamp 1677677812
transform 1 0 296 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_304
timestamp 1677677812
transform -1 0 344 0 -1 1370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_435
timestamp 1677677812
transform 1 0 344 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8055
timestamp 1677677812
transform 1 0 440 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_436
timestamp 1677677812
transform 1 0 448 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8056
timestamp 1677677812
transform 1 0 544 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_299
timestamp 1677677812
transform 1 0 552 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8057
timestamp 1677677812
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8058
timestamp 1677677812
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8059
timestamp 1677677812
transform 1 0 608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8060
timestamp 1677677812
transform 1 0 616 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_305
timestamp 1677677812
transform 1 0 624 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8061
timestamp 1677677812
transform 1 0 664 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8062
timestamp 1677677812
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_437
timestamp 1677677812
transform -1 0 776 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8063
timestamp 1677677812
transform 1 0 776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8065
timestamp 1677677812
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8067
timestamp 1677677812
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8069
timestamp 1677677812
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8071
timestamp 1677677812
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8072
timestamp 1677677812
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8073
timestamp 1677677812
transform 1 0 824 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8074
timestamp 1677677812
transform 1 0 832 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8075
timestamp 1677677812
transform 1 0 840 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8076
timestamp 1677677812
transform 1 0 848 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8078
timestamp 1677677812
transform 1 0 856 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8080
timestamp 1677677812
transform 1 0 864 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8082
timestamp 1677677812
transform 1 0 872 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8083
timestamp 1677677812
transform 1 0 880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8084
timestamp 1677677812
transform 1 0 888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8085
timestamp 1677677812
transform 1 0 896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8087
timestamp 1677677812
transform 1 0 904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8089
timestamp 1677677812
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8091
timestamp 1677677812
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6484
timestamp 1677677812
transform 1 0 940 0 1 1275
box -3 -3 3 3
use FILL  FILL_8095
timestamp 1677677812
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8096
timestamp 1677677812
transform 1 0 936 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6485
timestamp 1677677812
transform 1 0 972 0 1 1275
box -3 -3 3 3
use NOR2X1  NOR2X1_83
timestamp 1677677812
transform 1 0 944 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8097
timestamp 1677677812
transform 1 0 968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8099
timestamp 1677677812
transform 1 0 976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8101
timestamp 1677677812
transform 1 0 984 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8103
timestamp 1677677812
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8107
timestamp 1677677812
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8108
timestamp 1677677812
transform 1 0 1008 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8109
timestamp 1677677812
transform 1 0 1016 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_513
timestamp 1677677812
transform -1 0 1040 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8110
timestamp 1677677812
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8112
timestamp 1677677812
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8114
timestamp 1677677812
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8116
timestamp 1677677812
transform 1 0 1064 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8118
timestamp 1677677812
transform 1 0 1072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8120
timestamp 1677677812
transform 1 0 1080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8123
timestamp 1677677812
transform 1 0 1088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8124
timestamp 1677677812
transform 1 0 1096 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8125
timestamp 1677677812
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8126
timestamp 1677677812
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8128
timestamp 1677677812
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8130
timestamp 1677677812
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8132
timestamp 1677677812
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8134
timestamp 1677677812
transform 1 0 1144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8136
timestamp 1677677812
transform 1 0 1152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8138
timestamp 1677677812
transform 1 0 1160 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8140
timestamp 1677677812
transform 1 0 1168 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8142
timestamp 1677677812
transform 1 0 1176 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_85
timestamp 1677677812
transform 1 0 1184 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8144
timestamp 1677677812
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8145
timestamp 1677677812
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8146
timestamp 1677677812
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8148
timestamp 1677677812
transform 1 0 1232 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_303
timestamp 1677677812
transform 1 0 1240 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8168
timestamp 1677677812
transform 1 0 1280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8169
timestamp 1677677812
transform 1 0 1288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8170
timestamp 1677677812
transform 1 0 1296 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_438
timestamp 1677677812
transform 1 0 1304 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8171
timestamp 1677677812
transform 1 0 1400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8172
timestamp 1677677812
transform 1 0 1408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8173
timestamp 1677677812
transform 1 0 1416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8174
timestamp 1677677812
transform 1 0 1424 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_307
timestamp 1677677812
transform -1 0 1472 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8175
timestamp 1677677812
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8176
timestamp 1677677812
transform 1 0 1480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8184
timestamp 1677677812
transform 1 0 1488 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_440
timestamp 1677677812
transform -1 0 1592 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8185
timestamp 1677677812
transform 1 0 1592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8186
timestamp 1677677812
transform 1 0 1600 0 -1 1370
box -8 -3 16 105
use BUFX2  BUFX2_101
timestamp 1677677812
transform -1 0 1632 0 -1 1370
box -5 -3 28 105
use FILL  FILL_8187
timestamp 1677677812
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8193
timestamp 1677677812
transform 1 0 1640 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_308
timestamp 1677677812
transform 1 0 1648 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8194
timestamp 1677677812
transform 1 0 1688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8199
timestamp 1677677812
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8200
timestamp 1677677812
transform 1 0 1704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8201
timestamp 1677677812
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_305
timestamp 1677677812
transform 1 0 1720 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8202
timestamp 1677677812
transform 1 0 1760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8206
timestamp 1677677812
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8207
timestamp 1677677812
transform 1 0 1776 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_442
timestamp 1677677812
transform -1 0 1880 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8208
timestamp 1677677812
transform 1 0 1880 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8210
timestamp 1677677812
transform 1 0 1888 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8213
timestamp 1677677812
transform 1 0 1896 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8214
timestamp 1677677812
transform 1 0 1904 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8215
timestamp 1677677812
transform 1 0 1912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8216
timestamp 1677677812
transform 1 0 1920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8218
timestamp 1677677812
transform 1 0 1928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8229
timestamp 1677677812
transform 1 0 1936 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_518
timestamp 1677677812
transform -1 0 1960 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8230
timestamp 1677677812
transform 1 0 1960 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8231
timestamp 1677677812
transform 1 0 1968 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8232
timestamp 1677677812
transform 1 0 1976 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8233
timestamp 1677677812
transform 1 0 1984 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_307
timestamp 1677677812
transform -1 0 2032 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8234
timestamp 1677677812
transform 1 0 2032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8235
timestamp 1677677812
transform 1 0 2040 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_444
timestamp 1677677812
transform -1 0 2144 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8236
timestamp 1677677812
transform 1 0 2144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8238
timestamp 1677677812
transform 1 0 2152 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_63
timestamp 1677677812
transform -1 0 2192 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_519
timestamp 1677677812
transform 1 0 2192 0 -1 1370
box -9 -3 26 105
use M3_M2  M3_M2_6486
timestamp 1677677812
transform 1 0 2268 0 1 1275
box -3 -3 3 3
use M3_M2  M3_M2_6487
timestamp 1677677812
transform 1 0 2308 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_449
timestamp 1677677812
transform -1 0 2304 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8250
timestamp 1677677812
transform 1 0 2304 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_140
timestamp 1677677812
transform -1 0 2344 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8251
timestamp 1677677812
transform 1 0 2344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8252
timestamp 1677677812
transform 1 0 2352 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_11
timestamp 1677677812
transform -1 0 2384 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8253
timestamp 1677677812
transform 1 0 2384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8254
timestamp 1677677812
transform 1 0 2392 0 -1 1370
box -8 -3 16 105
use FAX1  FAX1_5
timestamp 1677677812
transform -1 0 2520 0 -1 1370
box -5 -3 126 105
use FILL  FILL_8255
timestamp 1677677812
transform 1 0 2520 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8256
timestamp 1677677812
transform 1 0 2528 0 -1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_0
timestamp 1677677812
transform -1 0 2592 0 -1 1370
box -8 -3 64 105
use FILL  FILL_8257
timestamp 1677677812
transform 1 0 2592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8258
timestamp 1677677812
transform 1 0 2600 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8259
timestamp 1677677812
transform 1 0 2608 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_308
timestamp 1677677812
transform 1 0 2616 0 -1 1370
box -8 -3 46 105
use AND2X2  AND2X2_51
timestamp 1677677812
transform 1 0 2656 0 -1 1370
box -8 -3 40 105
use XOR2X1  XOR2X1_1
timestamp 1677677812
transform -1 0 2744 0 -1 1370
box -8 -3 64 105
use FILL  FILL_8260
timestamp 1677677812
transform 1 0 2744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8261
timestamp 1677677812
transform 1 0 2752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8262
timestamp 1677677812
transform 1 0 2760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8263
timestamp 1677677812
transform 1 0 2768 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8264
timestamp 1677677812
transform 1 0 2776 0 -1 1370
box -8 -3 16 105
use FAX1  FAX1_7
timestamp 1677677812
transform 1 0 2784 0 -1 1370
box -5 -3 126 105
use BUFX2  BUFX2_102
timestamp 1677677812
transform 1 0 2904 0 -1 1370
box -5 -3 28 105
use FILL  FILL_8269
timestamp 1677677812
transform 1 0 2928 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8271
timestamp 1677677812
transform 1 0 2936 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8273
timestamp 1677677812
transform 1 0 2944 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8275
timestamp 1677677812
transform 1 0 2952 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8277
timestamp 1677677812
transform 1 0 2960 0 -1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_5
timestamp 1677677812
transform 1 0 2968 0 -1 1370
box -7 -3 39 105
use FILL  FILL_8283
timestamp 1677677812
transform 1 0 3000 0 -1 1370
box -8 -3 16 105
use AOI21X1  AOI21X1_6
timestamp 1677677812
transform 1 0 3008 0 -1 1370
box -7 -3 39 105
use FILL  FILL_8289
timestamp 1677677812
transform 1 0 3040 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_12
timestamp 1677677812
transform 1 0 3048 0 -1 1370
box -8 -3 32 105
use FILL  FILL_8290
timestamp 1677677812
transform 1 0 3072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8292
timestamp 1677677812
transform 1 0 3080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8294
timestamp 1677677812
transform 1 0 3088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8297
timestamp 1677677812
transform 1 0 3096 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_521
timestamp 1677677812
transform 1 0 3104 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8298
timestamp 1677677812
transform 1 0 3120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8308
timestamp 1677677812
transform 1 0 3128 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_142
timestamp 1677677812
transform -1 0 3168 0 -1 1370
box -8 -3 34 105
use AOI22X1  AOI22X1_310
timestamp 1677677812
transform 1 0 3168 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8309
timestamp 1677677812
transform 1 0 3208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8310
timestamp 1677677812
transform 1 0 3216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8311
timestamp 1677677812
transform 1 0 3224 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_522
timestamp 1677677812
transform 1 0 3232 0 -1 1370
box -9 -3 26 105
use INVX2  INVX2_523
timestamp 1677677812
transform -1 0 3264 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8312
timestamp 1677677812
transform 1 0 3264 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8314
timestamp 1677677812
transform 1 0 3272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8318
timestamp 1677677812
transform 1 0 3280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8319
timestamp 1677677812
transform 1 0 3288 0 -1 1370
box -8 -3 16 105
use AND2X1  AND2X1_0
timestamp 1677677812
transform 1 0 3296 0 -1 1370
box -8 -3 40 105
use FILL  FILL_8320
timestamp 1677677812
transform 1 0 3328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8326
timestamp 1677677812
transform 1 0 3336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8327
timestamp 1677677812
transform 1 0 3344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8328
timestamp 1677677812
transform 1 0 3352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8329
timestamp 1677677812
transform 1 0 3360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8330
timestamp 1677677812
transform 1 0 3368 0 -1 1370
box -8 -3 16 105
use FAX1  FAX1_10
timestamp 1677677812
transform -1 0 3496 0 -1 1370
box -5 -3 126 105
use FILL  FILL_8331
timestamp 1677677812
transform 1 0 3496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8332
timestamp 1677677812
transform 1 0 3504 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_450
timestamp 1677677812
transform 1 0 3512 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8333
timestamp 1677677812
transform 1 0 3608 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8334
timestamp 1677677812
transform 1 0 3616 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8335
timestamp 1677677812
transform 1 0 3624 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_524
timestamp 1677677812
transform 1 0 3632 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8336
timestamp 1677677812
transform 1 0 3648 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8337
timestamp 1677677812
transform 1 0 3656 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8338
timestamp 1677677812
transform 1 0 3664 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_309
timestamp 1677677812
transform 1 0 3672 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8345
timestamp 1677677812
transform 1 0 3712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8346
timestamp 1677677812
transform 1 0 3720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8347
timestamp 1677677812
transform 1 0 3728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8348
timestamp 1677677812
transform 1 0 3736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8350
timestamp 1677677812
transform 1 0 3744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8352
timestamp 1677677812
transform 1 0 3752 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_310
timestamp 1677677812
transform 1 0 3760 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8356
timestamp 1677677812
transform 1 0 3800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8357
timestamp 1677677812
transform 1 0 3808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8372
timestamp 1677677812
transform 1 0 3816 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_451
timestamp 1677677812
transform -1 0 3920 0 -1 1370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_452
timestamp 1677677812
transform 1 0 3920 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8373
timestamp 1677677812
transform 1 0 4016 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8374
timestamp 1677677812
transform 1 0 4024 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8376
timestamp 1677677812
transform 1 0 4032 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_146
timestamp 1677677812
transform 1 0 4040 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8386
timestamp 1677677812
transform 1 0 4072 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8387
timestamp 1677677812
transform 1 0 4080 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8388
timestamp 1677677812
transform 1 0 4088 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8389
timestamp 1677677812
transform 1 0 4096 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_311
timestamp 1677677812
transform 1 0 4104 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8390
timestamp 1677677812
transform 1 0 4144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8391
timestamp 1677677812
transform 1 0 4152 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8392
timestamp 1677677812
transform 1 0 4160 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_525
timestamp 1677677812
transform -1 0 4184 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8393
timestamp 1677677812
transform 1 0 4184 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8394
timestamp 1677677812
transform 1 0 4192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8395
timestamp 1677677812
transform 1 0 4200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8396
timestamp 1677677812
transform 1 0 4208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8397
timestamp 1677677812
transform 1 0 4216 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_526
timestamp 1677677812
transform -1 0 4240 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8398
timestamp 1677677812
transform 1 0 4240 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8399
timestamp 1677677812
transform 1 0 4248 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8400
timestamp 1677677812
transform 1 0 4256 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_312
timestamp 1677677812
transform 1 0 4264 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8411
timestamp 1677677812
transform 1 0 4304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8412
timestamp 1677677812
transform 1 0 4312 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8413
timestamp 1677677812
transform 1 0 4320 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8414
timestamp 1677677812
transform 1 0 4328 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_455
timestamp 1677677812
transform 1 0 4336 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8415
timestamp 1677677812
transform 1 0 4432 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8416
timestamp 1677677812
transform 1 0 4440 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_148
timestamp 1677677812
transform -1 0 4480 0 -1 1370
box -8 -3 34 105
use FILL  FILL_8417
timestamp 1677677812
transform 1 0 4480 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6488
timestamp 1677677812
transform 1 0 4556 0 1 1275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_456
timestamp 1677677812
transform 1 0 4488 0 -1 1370
box -8 -3 104 105
use FILL  FILL_8428
timestamp 1677677812
transform 1 0 4584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8429
timestamp 1677677812
transform 1 0 4592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8430
timestamp 1677677812
transform 1 0 4600 0 -1 1370
box -8 -3 16 105
use M3_M2  M3_M2_6489
timestamp 1677677812
transform 1 0 4636 0 1 1275
box -3 -3 3 3
use INVX2  INVX2_528
timestamp 1677677812
transform 1 0 4608 0 -1 1370
box -9 -3 26 105
use FILL  FILL_8431
timestamp 1677677812
transform 1 0 4624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8433
timestamp 1677677812
transform 1 0 4632 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8436
timestamp 1677677812
transform 1 0 4640 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_313
timestamp 1677677812
transform 1 0 4648 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8437
timestamp 1677677812
transform 1 0 4688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8438
timestamp 1677677812
transform 1 0 4696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8439
timestamp 1677677812
transform 1 0 4704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8440
timestamp 1677677812
transform 1 0 4712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8441
timestamp 1677677812
transform 1 0 4720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8442
timestamp 1677677812
transform 1 0 4728 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_314
timestamp 1677677812
transform -1 0 4776 0 -1 1370
box -8 -3 46 105
use FILL  FILL_8443
timestamp 1677677812
transform 1 0 4776 0 -1 1370
box -8 -3 16 105
use FILL  FILL_8445
timestamp 1677677812
transform 1 0 4784 0 -1 1370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_69
timestamp 1677677812
transform 1 0 4843 0 1 1270
box -10 -3 10 3
use M3_M2  M3_M2_6520
timestamp 1677677812
transform 1 0 188 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6548
timestamp 1677677812
transform 1 0 108 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7255
timestamp 1677677812
transform 1 0 148 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7359
timestamp 1677677812
transform 1 0 108 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7256
timestamp 1677677812
transform 1 0 196 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6619
timestamp 1677677812
transform 1 0 196 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6504
timestamp 1677677812
transform 1 0 268 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7257
timestamp 1677677812
transform 1 0 252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7258
timestamp 1677677812
transform 1 0 268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7360
timestamp 1677677812
transform 1 0 236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7361
timestamp 1677677812
transform 1 0 244 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6589
timestamp 1677677812
transform 1 0 228 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6505
timestamp 1677677812
transform 1 0 300 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7259
timestamp 1677677812
transform 1 0 284 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7260
timestamp 1677677812
transform 1 0 308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7362
timestamp 1677677812
transform 1 0 276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7363
timestamp 1677677812
transform 1 0 300 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7364
timestamp 1677677812
transform 1 0 316 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6620
timestamp 1677677812
transform 1 0 316 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6549
timestamp 1677677812
transform 1 0 356 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6521
timestamp 1677677812
transform 1 0 372 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7261
timestamp 1677677812
transform 1 0 372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7262
timestamp 1677677812
transform 1 0 404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7365
timestamp 1677677812
transform 1 0 396 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7366
timestamp 1677677812
transform 1 0 412 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7367
timestamp 1677677812
transform 1 0 420 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6590
timestamp 1677677812
transform 1 0 412 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7263
timestamp 1677677812
transform 1 0 476 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6522
timestamp 1677677812
transform 1 0 540 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6523
timestamp 1677677812
transform 1 0 580 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7264
timestamp 1677677812
transform 1 0 540 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7265
timestamp 1677677812
transform 1 0 572 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7266
timestamp 1677677812
transform 1 0 580 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7267
timestamp 1677677812
transform 1 0 588 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7368
timestamp 1677677812
transform 1 0 492 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6621
timestamp 1677677812
transform 1 0 572 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6524
timestamp 1677677812
transform 1 0 652 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7268
timestamp 1677677812
transform 1 0 628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7269
timestamp 1677677812
transform 1 0 644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7369
timestamp 1677677812
transform 1 0 612 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7370
timestamp 1677677812
transform 1 0 620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7371
timestamp 1677677812
transform 1 0 636 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6622
timestamp 1677677812
transform 1 0 636 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7372
timestamp 1677677812
transform 1 0 652 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6550
timestamp 1677677812
transform 1 0 668 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6525
timestamp 1677677812
transform 1 0 700 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7270
timestamp 1677677812
transform 1 0 692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7271
timestamp 1677677812
transform 1 0 700 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7373
timestamp 1677677812
transform 1 0 700 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6623
timestamp 1677677812
transform 1 0 700 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6526
timestamp 1677677812
transform 1 0 732 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7272
timestamp 1677677812
transform 1 0 740 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7374
timestamp 1677677812
transform 1 0 732 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6569
timestamp 1677677812
transform 1 0 740 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6527
timestamp 1677677812
transform 1 0 764 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7273
timestamp 1677677812
transform 1 0 780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7375
timestamp 1677677812
transform 1 0 780 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6506
timestamp 1677677812
transform 1 0 820 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7274
timestamp 1677677812
transform 1 0 812 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6551
timestamp 1677677812
transform 1 0 820 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7275
timestamp 1677677812
transform 1 0 836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7376
timestamp 1677677812
transform 1 0 804 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7377
timestamp 1677677812
transform 1 0 820 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7378
timestamp 1677677812
transform 1 0 828 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6591
timestamp 1677677812
transform 1 0 804 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6592
timestamp 1677677812
transform 1 0 860 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6507
timestamp 1677677812
transform 1 0 892 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6528
timestamp 1677677812
transform 1 0 884 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6529
timestamp 1677677812
transform 1 0 932 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7276
timestamp 1677677812
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7277
timestamp 1677677812
transform 1 0 892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7278
timestamp 1677677812
transform 1 0 932 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7379
timestamp 1677677812
transform 1 0 972 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6593
timestamp 1677677812
transform 1 0 972 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7279
timestamp 1677677812
transform 1 0 1028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7380
timestamp 1677677812
transform 1 0 1004 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6570
timestamp 1677677812
transform 1 0 1052 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6594
timestamp 1677677812
transform 1 0 1004 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7446
timestamp 1677677812
transform 1 0 1092 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6530
timestamp 1677677812
transform 1 0 1132 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7280
timestamp 1677677812
transform 1 0 1132 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6571
timestamp 1677677812
transform 1 0 1124 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7381
timestamp 1677677812
transform 1 0 1140 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7382
timestamp 1677677812
transform 1 0 1180 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6531
timestamp 1677677812
transform 1 0 1212 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6532
timestamp 1677677812
transform 1 0 1228 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7281
timestamp 1677677812
transform 1 0 1228 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6624
timestamp 1677677812
transform 1 0 1220 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6496
timestamp 1677677812
transform 1 0 1244 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6595
timestamp 1677677812
transform 1 0 1236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6508
timestamp 1677677812
transform 1 0 1268 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7282
timestamp 1677677812
transform 1 0 1252 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6552
timestamp 1677677812
transform 1 0 1260 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7283
timestamp 1677677812
transform 1 0 1268 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6497
timestamp 1677677812
transform 1 0 1284 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6553
timestamp 1677677812
transform 1 0 1284 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7383
timestamp 1677677812
transform 1 0 1260 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7384
timestamp 1677677812
transform 1 0 1276 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7385
timestamp 1677677812
transform 1 0 1284 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6596
timestamp 1677677812
transform 1 0 1260 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6597
timestamp 1677677812
transform 1 0 1276 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6625
timestamp 1677677812
transform 1 0 1276 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7284
timestamp 1677677812
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7285
timestamp 1677677812
transform 1 0 1348 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7286
timestamp 1677677812
transform 1 0 1364 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7386
timestamp 1677677812
transform 1 0 1332 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6598
timestamp 1677677812
transform 1 0 1332 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6554
timestamp 1677677812
transform 1 0 1372 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6572
timestamp 1677677812
transform 1 0 1348 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7287
timestamp 1677677812
transform 1 0 1396 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7387
timestamp 1677677812
transform 1 0 1372 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7388
timestamp 1677677812
transform 1 0 1380 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6573
timestamp 1677677812
transform 1 0 1388 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6599
timestamp 1677677812
transform 1 0 1388 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6626
timestamp 1677677812
transform 1 0 1396 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7288
timestamp 1677677812
transform 1 0 1420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7289
timestamp 1677677812
transform 1 0 1444 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7290
timestamp 1677677812
transform 1 0 1452 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7291
timestamp 1677677812
transform 1 0 1468 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6574
timestamp 1677677812
transform 1 0 1436 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7292
timestamp 1677677812
transform 1 0 1492 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7389
timestamp 1677677812
transform 1 0 1460 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7390
timestamp 1677677812
transform 1 0 1476 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7391
timestamp 1677677812
transform 1 0 1484 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6600
timestamp 1677677812
transform 1 0 1460 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6627
timestamp 1677677812
transform 1 0 1452 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6575
timestamp 1677677812
transform 1 0 1492 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7293
timestamp 1677677812
transform 1 0 1532 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6498
timestamp 1677677812
transform 1 0 1556 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7294
timestamp 1677677812
transform 1 0 1556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7392
timestamp 1677677812
transform 1 0 1548 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7393
timestamp 1677677812
transform 1 0 1564 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6509
timestamp 1677677812
transform 1 0 1604 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7295
timestamp 1677677812
transform 1 0 1596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7296
timestamp 1677677812
transform 1 0 1604 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6499
timestamp 1677677812
transform 1 0 1636 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6533
timestamp 1677677812
transform 1 0 1628 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7297
timestamp 1677677812
transform 1 0 1636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7394
timestamp 1677677812
transform 1 0 1604 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7395
timestamp 1677677812
transform 1 0 1612 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6601
timestamp 1677677812
transform 1 0 1596 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6576
timestamp 1677677812
transform 1 0 1620 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7396
timestamp 1677677812
transform 1 0 1628 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6510
timestamp 1677677812
transform 1 0 1652 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6534
timestamp 1677677812
transform 1 0 1660 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7397
timestamp 1677677812
transform 1 0 1660 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6535
timestamp 1677677812
transform 1 0 1756 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7298
timestamp 1677677812
transform 1 0 1700 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6555
timestamp 1677677812
transform 1 0 1716 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7299
timestamp 1677677812
transform 1 0 1756 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7398
timestamp 1677677812
transform 1 0 1676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7399
timestamp 1677677812
transform 1 0 1764 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7300
timestamp 1677677812
transform 1 0 1780 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7301
timestamp 1677677812
transform 1 0 1788 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7302
timestamp 1677677812
transform 1 0 1836 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7303
timestamp 1677677812
transform 1 0 1884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7304
timestamp 1677677812
transform 1 0 1940 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6577
timestamp 1677677812
transform 1 0 1788 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6578
timestamp 1677677812
transform 1 0 1804 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7400
timestamp 1677677812
transform 1 0 1868 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6602
timestamp 1677677812
transform 1 0 1868 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7401
timestamp 1677677812
transform 1 0 1964 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6603
timestamp 1677677812
transform 1 0 1900 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6604
timestamp 1677677812
transform 1 0 1964 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7305
timestamp 1677677812
transform 1 0 2028 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7306
timestamp 1677677812
transform 1 0 2108 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7402
timestamp 1677677812
transform 1 0 2132 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6628
timestamp 1677677812
transform 1 0 2196 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6490
timestamp 1677677812
transform 1 0 2308 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6556
timestamp 1677677812
transform 1 0 2220 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6557
timestamp 1677677812
transform 1 0 2244 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6500
timestamp 1677677812
transform 1 0 2324 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7250
timestamp 1677677812
transform 1 0 2324 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7307
timestamp 1677677812
transform 1 0 2268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7308
timestamp 1677677812
transform 1 0 2308 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7309
timestamp 1677677812
transform 1 0 2316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7403
timestamp 1677677812
transform 1 0 2220 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6605
timestamp 1677677812
transform 1 0 2220 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6606
timestamp 1677677812
transform 1 0 2300 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6629
timestamp 1677677812
transform 1 0 2212 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6501
timestamp 1677677812
transform 1 0 2348 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7310
timestamp 1677677812
transform 1 0 2340 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6607
timestamp 1677677812
transform 1 0 2332 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7251
timestamp 1677677812
transform 1 0 2372 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7404
timestamp 1677677812
transform 1 0 2348 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6579
timestamp 1677677812
transform 1 0 2356 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7405
timestamp 1677677812
transform 1 0 2388 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7311
timestamp 1677677812
transform 1 0 2404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7312
timestamp 1677677812
transform 1 0 2436 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7406
timestamp 1677677812
transform 1 0 2420 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7407
timestamp 1677677812
transform 1 0 2436 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6536
timestamp 1677677812
transform 1 0 2452 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7313
timestamp 1677677812
transform 1 0 2460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7447
timestamp 1677677812
transform 1 0 2452 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6537
timestamp 1677677812
transform 1 0 2492 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7314
timestamp 1677677812
transform 1 0 2484 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7315
timestamp 1677677812
transform 1 0 2492 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6580
timestamp 1677677812
transform 1 0 2484 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6581
timestamp 1677677812
transform 1 0 2500 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7448
timestamp 1677677812
transform 1 0 2500 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6491
timestamp 1677677812
transform 1 0 2532 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6538
timestamp 1677677812
transform 1 0 2516 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7316
timestamp 1677677812
transform 1 0 2524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7408
timestamp 1677677812
transform 1 0 2516 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6582
timestamp 1677677812
transform 1 0 2524 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6511
timestamp 1677677812
transform 1 0 2548 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7409
timestamp 1677677812
transform 1 0 2548 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6558
timestamp 1677677812
transform 1 0 2556 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_6539
timestamp 1677677812
transform 1 0 2580 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7317
timestamp 1677677812
transform 1 0 2564 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7318
timestamp 1677677812
transform 1 0 2580 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6559
timestamp 1677677812
transform 1 0 2588 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7410
timestamp 1677677812
transform 1 0 2572 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6502
timestamp 1677677812
transform 1 0 2620 0 1 1245
box -3 -3 3 3
use M2_M1  M2_M1_7411
timestamp 1677677812
transform 1 0 2620 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6503
timestamp 1677677812
transform 1 0 2644 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_6512
timestamp 1677677812
transform 1 0 2636 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6540
timestamp 1677677812
transform 1 0 2636 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7319
timestamp 1677677812
transform 1 0 2636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7320
timestamp 1677677812
transform 1 0 2644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7321
timestamp 1677677812
transform 1 0 2700 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6560
timestamp 1677677812
transform 1 0 2724 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7412
timestamp 1677677812
transform 1 0 2724 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6541
timestamp 1677677812
transform 1 0 2740 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7322
timestamp 1677677812
transform 1 0 2740 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6542
timestamp 1677677812
transform 1 0 2804 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_6561
timestamp 1677677812
transform 1 0 2764 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7323
timestamp 1677677812
transform 1 0 2804 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6562
timestamp 1677677812
transform 1 0 2828 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7413
timestamp 1677677812
transform 1 0 2828 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6608
timestamp 1677677812
transform 1 0 2804 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6543
timestamp 1677677812
transform 1 0 2852 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7324
timestamp 1677677812
transform 1 0 2844 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7414
timestamp 1677677812
transform 1 0 2844 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6609
timestamp 1677677812
transform 1 0 2844 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6513
timestamp 1677677812
transform 1 0 2868 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6514
timestamp 1677677812
transform 1 0 2908 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7325
timestamp 1677677812
transform 1 0 2876 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6583
timestamp 1677677812
transform 1 0 2876 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7415
timestamp 1677677812
transform 1 0 2972 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7416
timestamp 1677677812
transform 1 0 2980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7449
timestamp 1677677812
transform 1 0 2964 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_6584
timestamp 1677677812
transform 1 0 2996 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6515
timestamp 1677677812
transform 1 0 3012 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7252
timestamp 1677677812
transform 1 0 3012 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7253
timestamp 1677677812
transform 1 0 3028 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7326
timestamp 1677677812
transform 1 0 3036 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7249
timestamp 1677677812
transform 1 0 3052 0 1 1235
box -2 -2 2 2
use M3_M2  M3_M2_6516
timestamp 1677677812
transform 1 0 3068 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7327
timestamp 1677677812
transform 1 0 3060 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6610
timestamp 1677677812
transform 1 0 3100 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7328
timestamp 1677677812
transform 1 0 3124 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7329
timestamp 1677677812
transform 1 0 3172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7254
timestamp 1677677812
transform 1 0 3188 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_7330
timestamp 1677677812
transform 1 0 3268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7450
timestamp 1677677812
transform 1 0 3324 0 1 1195
box -2 -2 2 2
use M2_M1  M2_M1_7417
timestamp 1677677812
transform 1 0 3356 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7331
timestamp 1677677812
transform 1 0 3484 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6544
timestamp 1677677812
transform 1 0 3556 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7332
timestamp 1677677812
transform 1 0 3556 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7418
timestamp 1677677812
transform 1 0 3508 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6630
timestamp 1677677812
transform 1 0 3524 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7333
timestamp 1677677812
transform 1 0 3596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7419
timestamp 1677677812
transform 1 0 3604 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6631
timestamp 1677677812
transform 1 0 3604 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6545
timestamp 1677677812
transform 1 0 3628 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7334
timestamp 1677677812
transform 1 0 3620 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7335
timestamp 1677677812
transform 1 0 3636 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7420
timestamp 1677677812
transform 1 0 3628 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6585
timestamp 1677677812
transform 1 0 3636 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7336
timestamp 1677677812
transform 1 0 3660 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6632
timestamp 1677677812
transform 1 0 3652 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6563
timestamp 1677677812
transform 1 0 3676 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7421
timestamp 1677677812
transform 1 0 3676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7422
timestamp 1677677812
transform 1 0 3684 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6564
timestamp 1677677812
transform 1 0 3708 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7337
timestamp 1677677812
transform 1 0 3716 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7423
timestamp 1677677812
transform 1 0 3708 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7338
timestamp 1677677812
transform 1 0 3772 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6492
timestamp 1677677812
transform 1 0 3788 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7339
timestamp 1677677812
transform 1 0 3812 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7424
timestamp 1677677812
transform 1 0 3844 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6586
timestamp 1677677812
transform 1 0 3852 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6517
timestamp 1677677812
transform 1 0 3988 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7340
timestamp 1677677812
transform 1 0 3940 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7341
timestamp 1677677812
transform 1 0 3972 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6565
timestamp 1677677812
transform 1 0 3980 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7342
timestamp 1677677812
transform 1 0 3988 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7425
timestamp 1677677812
transform 1 0 3892 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7426
timestamp 1677677812
transform 1 0 3980 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7427
timestamp 1677677812
transform 1 0 3996 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7428
timestamp 1677677812
transform 1 0 4012 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6611
timestamp 1677677812
transform 1 0 3892 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6633
timestamp 1677677812
transform 1 0 4012 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7343
timestamp 1677677812
transform 1 0 4044 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7429
timestamp 1677677812
transform 1 0 4068 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6634
timestamp 1677677812
transform 1 0 4084 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_6566
timestamp 1677677812
transform 1 0 4140 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7344
timestamp 1677677812
transform 1 0 4164 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7345
timestamp 1677677812
transform 1 0 4220 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7346
timestamp 1677677812
transform 1 0 4260 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7347
timestamp 1677677812
transform 1 0 4316 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7430
timestamp 1677677812
transform 1 0 4140 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6612
timestamp 1677677812
transform 1 0 4140 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7431
timestamp 1677677812
transform 1 0 4236 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6613
timestamp 1677677812
transform 1 0 4236 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6546
timestamp 1677677812
transform 1 0 4332 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7432
timestamp 1677677812
transform 1 0 4332 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6518
timestamp 1677677812
transform 1 0 4356 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_7348
timestamp 1677677812
transform 1 0 4356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7433
timestamp 1677677812
transform 1 0 4364 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7434
timestamp 1677677812
transform 1 0 4380 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7349
timestamp 1677677812
transform 1 0 4404 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7435
timestamp 1677677812
transform 1 0 4428 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6614
timestamp 1677677812
transform 1 0 4420 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6615
timestamp 1677677812
transform 1 0 4444 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7350
timestamp 1677677812
transform 1 0 4460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7351
timestamp 1677677812
transform 1 0 4468 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6587
timestamp 1677677812
transform 1 0 4476 0 1 1205
box -3 -3 3 3
use M3_M2  M3_M2_6616
timestamp 1677677812
transform 1 0 4468 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6567
timestamp 1677677812
transform 1 0 4484 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7436
timestamp 1677677812
transform 1 0 4500 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6493
timestamp 1677677812
transform 1 0 4524 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6547
timestamp 1677677812
transform 1 0 4516 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_7352
timestamp 1677677812
transform 1 0 4508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7353
timestamp 1677677812
transform 1 0 4524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7354
timestamp 1677677812
transform 1 0 4540 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_6568
timestamp 1677677812
transform 1 0 4548 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_7437
timestamp 1677677812
transform 1 0 4516 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6588
timestamp 1677677812
transform 1 0 4524 0 1 1205
box -3 -3 3 3
use M2_M1  M2_M1_7438
timestamp 1677677812
transform 1 0 4532 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7439
timestamp 1677677812
transform 1 0 4548 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6617
timestamp 1677677812
transform 1 0 4540 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_6635
timestamp 1677677812
transform 1 0 4548 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_7440
timestamp 1677677812
transform 1 0 4564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7441
timestamp 1677677812
transform 1 0 4588 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6618
timestamp 1677677812
transform 1 0 4588 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_7355
timestamp 1677677812
transform 1 0 4596 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7356
timestamp 1677677812
transform 1 0 4628 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7357
timestamp 1677677812
transform 1 0 4644 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7442
timestamp 1677677812
transform 1 0 4620 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7443
timestamp 1677677812
transform 1 0 4636 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_7444
timestamp 1677677812
transform 1 0 4652 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_6519
timestamp 1677677812
transform 1 0 4684 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_6494
timestamp 1677677812
transform 1 0 4732 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_6495
timestamp 1677677812
transform 1 0 4748 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_7358
timestamp 1677677812
transform 1 0 4764 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_7445
timestamp 1677677812
transform 1 0 4788 0 1 1205
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_70
timestamp 1677677812
transform 1 0 48 0 1 1170
box -10 -3 10 3
use FILL  FILL_8446
timestamp 1677677812
transform 1 0 72 0 1 1170
box -8 -3 16 105
use FILL  FILL_8448
timestamp 1677677812
transform 1 0 80 0 1 1170
box -8 -3 16 105
use FILL  FILL_8450
timestamp 1677677812
transform 1 0 88 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_458
timestamp 1677677812
transform 1 0 96 0 1 1170
box -8 -3 104 105
use FILL  FILL_8452
timestamp 1677677812
transform 1 0 192 0 1 1170
box -8 -3 16 105
use FILL  FILL_8453
timestamp 1677677812
transform 1 0 200 0 1 1170
box -8 -3 16 105
use FILL  FILL_8454
timestamp 1677677812
transform 1 0 208 0 1 1170
box -8 -3 16 105
use FILL  FILL_8455
timestamp 1677677812
transform 1 0 216 0 1 1170
box -8 -3 16 105
use FILL  FILL_8456
timestamp 1677677812
transform 1 0 224 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_311
timestamp 1677677812
transform 1 0 232 0 1 1170
box -8 -3 46 105
use FILL  FILL_8457
timestamp 1677677812
transform 1 0 272 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6636
timestamp 1677677812
transform 1 0 300 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_315
timestamp 1677677812
transform 1 0 280 0 1 1170
box -8 -3 46 105
use FILL  FILL_8458
timestamp 1677677812
transform 1 0 320 0 1 1170
box -8 -3 16 105
use FILL  FILL_8459
timestamp 1677677812
transform 1 0 328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8460
timestamp 1677677812
transform 1 0 336 0 1 1170
box -8 -3 16 105
use FILL  FILL_8461
timestamp 1677677812
transform 1 0 344 0 1 1170
box -8 -3 16 105
use FILL  FILL_8462
timestamp 1677677812
transform 1 0 352 0 1 1170
box -8 -3 16 105
use FILL  FILL_8463
timestamp 1677677812
transform 1 0 360 0 1 1170
box -8 -3 16 105
use FILL  FILL_8464
timestamp 1677677812
transform 1 0 368 0 1 1170
box -8 -3 16 105
use FILL  FILL_8477
timestamp 1677677812
transform 1 0 376 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_313
timestamp 1677677812
transform -1 0 424 0 1 1170
box -8 -3 46 105
use FILL  FILL_8478
timestamp 1677677812
transform 1 0 424 0 1 1170
box -8 -3 16 105
use FILL  FILL_8486
timestamp 1677677812
transform 1 0 432 0 1 1170
box -8 -3 16 105
use FILL  FILL_8487
timestamp 1677677812
transform 1 0 440 0 1 1170
box -8 -3 16 105
use FILL  FILL_8488
timestamp 1677677812
transform 1 0 448 0 1 1170
box -8 -3 16 105
use FILL  FILL_8489
timestamp 1677677812
transform 1 0 456 0 1 1170
box -8 -3 16 105
use FILL  FILL_8490
timestamp 1677677812
transform 1 0 464 0 1 1170
box -8 -3 16 105
use FILL  FILL_8491
timestamp 1677677812
transform 1 0 472 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_460
timestamp 1677677812
transform 1 0 480 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_534
timestamp 1677677812
transform -1 0 592 0 1 1170
box -9 -3 26 105
use FILL  FILL_8492
timestamp 1677677812
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8507
timestamp 1677677812
transform 1 0 600 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_314
timestamp 1677677812
transform 1 0 608 0 1 1170
box -8 -3 46 105
use FILL  FILL_8509
timestamp 1677677812
transform 1 0 648 0 1 1170
box -8 -3 16 105
use FILL  FILL_8516
timestamp 1677677812
transform 1 0 656 0 1 1170
box -8 -3 16 105
use FILL  FILL_8518
timestamp 1677677812
transform 1 0 664 0 1 1170
box -8 -3 16 105
use BUFX2  BUFX2_105
timestamp 1677677812
transform -1 0 696 0 1 1170
box -5 -3 28 105
use FILL  FILL_8519
timestamp 1677677812
transform 1 0 696 0 1 1170
box -8 -3 16 105
use FILL  FILL_8520
timestamp 1677677812
transform 1 0 704 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_317
timestamp 1677677812
transform 1 0 712 0 1 1170
box -8 -3 46 105
use FILL  FILL_8521
timestamp 1677677812
transform 1 0 752 0 1 1170
box -8 -3 16 105
use FILL  FILL_8522
timestamp 1677677812
transform 1 0 760 0 1 1170
box -8 -3 16 105
use FILL  FILL_8523
timestamp 1677677812
transform 1 0 768 0 1 1170
box -8 -3 16 105
use FILL  FILL_8524
timestamp 1677677812
transform 1 0 776 0 1 1170
box -8 -3 16 105
use FILL  FILL_8525
timestamp 1677677812
transform 1 0 784 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_315
timestamp 1677677812
transform 1 0 792 0 1 1170
box -8 -3 46 105
use FILL  FILL_8530
timestamp 1677677812
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_8531
timestamp 1677677812
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_8532
timestamp 1677677812
transform 1 0 848 0 1 1170
box -8 -3 16 105
use FILL  FILL_8533
timestamp 1677677812
transform 1 0 856 0 1 1170
box -8 -3 16 105
use FILL  FILL_8534
timestamp 1677677812
transform 1 0 864 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_536
timestamp 1677677812
transform 1 0 872 0 1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_462
timestamp 1677677812
transform -1 0 984 0 1 1170
box -8 -3 104 105
use FILL  FILL_8535
timestamp 1677677812
transform 1 0 984 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6637
timestamp 1677677812
transform 1 0 1092 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_463
timestamp 1677677812
transform 1 0 992 0 1 1170
box -8 -3 104 105
use FILL  FILL_8536
timestamp 1677677812
transform 1 0 1088 0 1 1170
box -8 -3 16 105
use FILL  FILL_8537
timestamp 1677677812
transform 1 0 1096 0 1 1170
box -8 -3 16 105
use FILL  FILL_8538
timestamp 1677677812
transform 1 0 1104 0 1 1170
box -8 -3 16 105
use FILL  FILL_8539
timestamp 1677677812
transform 1 0 1112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8552
timestamp 1677677812
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_88
timestamp 1677677812
transform 1 0 1128 0 1 1170
box -8 -3 32 105
use FILL  FILL_8554
timestamp 1677677812
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_8555
timestamp 1677677812
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use FILL  FILL_8556
timestamp 1677677812
transform 1 0 1168 0 1 1170
box -8 -3 16 105
use FILL  FILL_8557
timestamp 1677677812
transform 1 0 1176 0 1 1170
box -8 -3 16 105
use FILL  FILL_8558
timestamp 1677677812
transform 1 0 1184 0 1 1170
box -8 -3 16 105
use FILL  FILL_8559
timestamp 1677677812
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_8564
timestamp 1677677812
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use FILL  FILL_8566
timestamp 1677677812
transform 1 0 1208 0 1 1170
box -8 -3 16 105
use FILL  FILL_8568
timestamp 1677677812
transform 1 0 1216 0 1 1170
box -8 -3 16 105
use FILL  FILL_8570
timestamp 1677677812
transform 1 0 1224 0 1 1170
box -8 -3 16 105
use FILL  FILL_8572
timestamp 1677677812
transform 1 0 1232 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6638
timestamp 1677677812
transform 1 0 1252 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_318
timestamp 1677677812
transform -1 0 1280 0 1 1170
box -8 -3 46 105
use FILL  FILL_8573
timestamp 1677677812
transform 1 0 1280 0 1 1170
box -8 -3 16 105
use FILL  FILL_8581
timestamp 1677677812
transform 1 0 1288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8583
timestamp 1677677812
transform 1 0 1296 0 1 1170
box -8 -3 16 105
use FILL  FILL_8585
timestamp 1677677812
transform 1 0 1304 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_540
timestamp 1677677812
transform 1 0 1312 0 1 1170
box -9 -3 26 105
use FILL  FILL_8586
timestamp 1677677812
transform 1 0 1328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8587
timestamp 1677677812
transform 1 0 1336 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6639
timestamp 1677677812
transform 1 0 1356 0 1 1175
box -3 -3 3 3
use AOI22X1  AOI22X1_318
timestamp 1677677812
transform -1 0 1384 0 1 1170
box -8 -3 46 105
use FILL  FILL_8588
timestamp 1677677812
transform 1 0 1384 0 1 1170
box -8 -3 16 105
use FILL  FILL_8589
timestamp 1677677812
transform 1 0 1392 0 1 1170
box -8 -3 16 105
use FILL  FILL_8590
timestamp 1677677812
transform 1 0 1400 0 1 1170
box -8 -3 16 105
use FILL  FILL_8591
timestamp 1677677812
transform 1 0 1408 0 1 1170
box -8 -3 16 105
use FILL  FILL_8592
timestamp 1677677812
transform 1 0 1416 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_541
timestamp 1677677812
transform 1 0 1424 0 1 1170
box -9 -3 26 105
use FILL  FILL_8593
timestamp 1677677812
transform 1 0 1440 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_319
timestamp 1677677812
transform 1 0 1448 0 1 1170
box -8 -3 46 105
use FILL  FILL_8594
timestamp 1677677812
transform 1 0 1488 0 1 1170
box -8 -3 16 105
use FILL  FILL_8600
timestamp 1677677812
transform 1 0 1496 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_543
timestamp 1677677812
transform 1 0 1504 0 1 1170
box -9 -3 26 105
use FILL  FILL_8601
timestamp 1677677812
transform 1 0 1520 0 1 1170
box -8 -3 16 105
use FILL  FILL_8602
timestamp 1677677812
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_8603
timestamp 1677677812
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_319
timestamp 1677677812
transform -1 0 1584 0 1 1170
box -8 -3 46 105
use FILL  FILL_8604
timestamp 1677677812
transform 1 0 1584 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6640
timestamp 1677677812
transform 1 0 1604 0 1 1175
box -3 -3 3 3
use FILL  FILL_8605
timestamp 1677677812
transform 1 0 1592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8607
timestamp 1677677812
transform 1 0 1600 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_320
timestamp 1677677812
transform 1 0 1608 0 1 1170
box -8 -3 46 105
use FILL  FILL_8609
timestamp 1677677812
transform 1 0 1648 0 1 1170
box -8 -3 16 105
use FILL  FILL_8610
timestamp 1677677812
transform 1 0 1656 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_467
timestamp 1677677812
transform 1 0 1664 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_544
timestamp 1677677812
transform 1 0 1760 0 1 1170
box -9 -3 26 105
use FILL  FILL_8613
timestamp 1677677812
transform 1 0 1776 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_468
timestamp 1677677812
transform -1 0 1880 0 1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_469
timestamp 1677677812
transform -1 0 1976 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_6641
timestamp 1677677812
transform 1 0 1988 0 1 1175
box -3 -3 3 3
use FILL  FILL_8614
timestamp 1677677812
transform 1 0 1976 0 1 1170
box -8 -3 16 105
use FILL  FILL_8615
timestamp 1677677812
transform 1 0 1984 0 1 1170
box -8 -3 16 105
use FILL  FILL_8616
timestamp 1677677812
transform 1 0 1992 0 1 1170
box -8 -3 16 105
use FILL  FILL_8617
timestamp 1677677812
transform 1 0 2000 0 1 1170
box -8 -3 16 105
use FILL  FILL_8638
timestamp 1677677812
transform 1 0 2008 0 1 1170
box -8 -3 16 105
use FILL  FILL_8640
timestamp 1677677812
transform 1 0 2016 0 1 1170
box -8 -3 16 105
use FILL  FILL_8642
timestamp 1677677812
transform 1 0 2024 0 1 1170
box -8 -3 16 105
use FILL  FILL_8643
timestamp 1677677812
transform 1 0 2032 0 1 1170
box -8 -3 16 105
use FILL  FILL_8644
timestamp 1677677812
transform 1 0 2040 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6642
timestamp 1677677812
transform 1 0 2068 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_470
timestamp 1677677812
transform -1 0 2144 0 1 1170
box -8 -3 104 105
use FILL  FILL_8645
timestamp 1677677812
transform 1 0 2144 0 1 1170
box -8 -3 16 105
use FILL  FILL_8646
timestamp 1677677812
transform 1 0 2152 0 1 1170
box -8 -3 16 105
use FILL  FILL_8647
timestamp 1677677812
transform 1 0 2160 0 1 1170
box -8 -3 16 105
use FILL  FILL_8648
timestamp 1677677812
transform 1 0 2168 0 1 1170
box -8 -3 16 105
use FILL  FILL_8649
timestamp 1677677812
transform 1 0 2176 0 1 1170
box -8 -3 16 105
use FILL  FILL_8650
timestamp 1677677812
transform 1 0 2184 0 1 1170
box -8 -3 16 105
use FILL  FILL_8651
timestamp 1677677812
transform 1 0 2192 0 1 1170
box -8 -3 16 105
use FILL  FILL_8654
timestamp 1677677812
transform 1 0 2200 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_472
timestamp 1677677812
transform 1 0 2208 0 1 1170
box -8 -3 104 105
use NAND2X1  NAND2X1_17
timestamp 1677677812
transform 1 0 2304 0 1 1170
box -8 -3 32 105
use FILL  FILL_8656
timestamp 1677677812
transform 1 0 2328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8669
timestamp 1677677812
transform 1 0 2336 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_151
timestamp 1677677812
transform 1 0 2344 0 1 1170
box -8 -3 34 105
use FILL  FILL_8670
timestamp 1677677812
transform 1 0 2376 0 1 1170
box -8 -3 16 105
use FILL  FILL_8674
timestamp 1677677812
transform 1 0 2384 0 1 1170
box -8 -3 16 105
use FILL  FILL_8675
timestamp 1677677812
transform 1 0 2392 0 1 1170
box -8 -3 16 105
use FILL  FILL_8676
timestamp 1677677812
transform 1 0 2400 0 1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_9
timestamp 1677677812
transform 1 0 2408 0 1 1170
box -7 -3 39 105
use FILL  FILL_8677
timestamp 1677677812
transform 1 0 2440 0 1 1170
box -8 -3 16 105
use FILL  FILL_8678
timestamp 1677677812
transform 1 0 2448 0 1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_10
timestamp 1677677812
transform 1 0 2456 0 1 1170
box -7 -3 39 105
use FILL  FILL_8679
timestamp 1677677812
transform 1 0 2488 0 1 1170
box -8 -3 16 105
use FILL  FILL_8680
timestamp 1677677812
transform 1 0 2496 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_551
timestamp 1677677812
transform -1 0 2520 0 1 1170
box -9 -3 26 105
use FILL  FILL_8681
timestamp 1677677812
transform 1 0 2520 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_552
timestamp 1677677812
transform -1 0 2544 0 1 1170
box -9 -3 26 105
use FILL  FILL_8682
timestamp 1677677812
transform 1 0 2544 0 1 1170
box -8 -3 16 105
use FILL  FILL_8683
timestamp 1677677812
transform 1 0 2552 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_325
timestamp 1677677812
transform 1 0 2560 0 1 1170
box -8 -3 46 105
use M3_M2  M3_M2_6643
timestamp 1677677812
transform 1 0 2612 0 1 1175
box -3 -3 3 3
use FILL  FILL_8684
timestamp 1677677812
transform 1 0 2600 0 1 1170
box -8 -3 16 105
use FILL  FILL_8685
timestamp 1677677812
transform 1 0 2608 0 1 1170
box -8 -3 16 105
use FILL  FILL_8686
timestamp 1677677812
transform 1 0 2616 0 1 1170
box -8 -3 16 105
use FILL  FILL_8687
timestamp 1677677812
transform 1 0 2624 0 1 1170
box -8 -3 16 105
use FILL  FILL_8688
timestamp 1677677812
transform 1 0 2632 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6644
timestamp 1677677812
transform 1 0 2668 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_473
timestamp 1677677812
transform -1 0 2736 0 1 1170
box -8 -3 104 105
use FILL  FILL_8689
timestamp 1677677812
transform 1 0 2736 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_474
timestamp 1677677812
transform -1 0 2840 0 1 1170
box -8 -3 104 105
use FILL  FILL_8690
timestamp 1677677812
transform 1 0 2840 0 1 1170
box -8 -3 16 105
use FILL  FILL_8691
timestamp 1677677812
transform 1 0 2848 0 1 1170
box -8 -3 16 105
use FAX1  FAX1_11
timestamp 1677677812
transform 1 0 2856 0 1 1170
box -5 -3 126 105
use NAND2X1  NAND2X1_19
timestamp 1677677812
transform 1 0 2976 0 1 1170
box -8 -3 32 105
use FILL  FILL_8692
timestamp 1677677812
transform 1 0 3000 0 1 1170
box -8 -3 16 105
use FILL  FILL_8693
timestamp 1677677812
transform 1 0 3008 0 1 1170
box -8 -3 16 105
use FILL  FILL_8694
timestamp 1677677812
transform 1 0 3016 0 1 1170
box -8 -3 16 105
use FILL  FILL_8695
timestamp 1677677812
transform 1 0 3024 0 1 1170
box -8 -3 16 105
use FILL  FILL_8696
timestamp 1677677812
transform 1 0 3032 0 1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_67
timestamp 1677677812
transform -1 0 3072 0 1 1170
box -8 -3 40 105
use FILL  FILL_8697
timestamp 1677677812
transform 1 0 3072 0 1 1170
box -8 -3 16 105
use FILL  FILL_8698
timestamp 1677677812
transform 1 0 3080 0 1 1170
box -8 -3 16 105
use FILL  FILL_8699
timestamp 1677677812
transform 1 0 3088 0 1 1170
box -8 -3 16 105
use FILL  FILL_8700
timestamp 1677677812
transform 1 0 3096 0 1 1170
box -8 -3 16 105
use FILL  FILL_8701
timestamp 1677677812
transform 1 0 3104 0 1 1170
box -8 -3 16 105
use FILL  FILL_8702
timestamp 1677677812
transform 1 0 3112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8729
timestamp 1677677812
transform 1 0 3120 0 1 1170
box -8 -3 16 105
use FILL  FILL_8730
timestamp 1677677812
transform 1 0 3128 0 1 1170
box -8 -3 16 105
use FILL  FILL_8731
timestamp 1677677812
transform 1 0 3136 0 1 1170
box -8 -3 16 105
use FILL  FILL_8732
timestamp 1677677812
transform 1 0 3144 0 1 1170
box -8 -3 16 105
use FILL  FILL_8733
timestamp 1677677812
transform 1 0 3152 0 1 1170
box -8 -3 16 105
use FILL  FILL_8735
timestamp 1677677812
transform 1 0 3160 0 1 1170
box -8 -3 16 105
use FILL  FILL_8737
timestamp 1677677812
transform 1 0 3168 0 1 1170
box -8 -3 16 105
use FILL  FILL_8739
timestamp 1677677812
transform 1 0 3176 0 1 1170
box -8 -3 16 105
use FILL  FILL_8740
timestamp 1677677812
transform 1 0 3184 0 1 1170
box -8 -3 16 105
use FILL  FILL_8741
timestamp 1677677812
transform 1 0 3192 0 1 1170
box -8 -3 16 105
use FILL  FILL_8742
timestamp 1677677812
transform 1 0 3200 0 1 1170
box -8 -3 16 105
use FILL  FILL_8743
timestamp 1677677812
transform 1 0 3208 0 1 1170
box -8 -3 16 105
use FILL  FILL_8744
timestamp 1677677812
transform 1 0 3216 0 1 1170
box -8 -3 16 105
use FILL  FILL_8747
timestamp 1677677812
transform 1 0 3224 0 1 1170
box -8 -3 16 105
use FILL  FILL_8749
timestamp 1677677812
transform 1 0 3232 0 1 1170
box -8 -3 16 105
use FILL  FILL_8750
timestamp 1677677812
transform 1 0 3240 0 1 1170
box -8 -3 16 105
use FILL  FILL_8751
timestamp 1677677812
transform 1 0 3248 0 1 1170
box -8 -3 16 105
use FILL  FILL_8753
timestamp 1677677812
transform 1 0 3256 0 1 1170
box -8 -3 16 105
use FILL  FILL_8754
timestamp 1677677812
transform 1 0 3264 0 1 1170
box -8 -3 16 105
use FILL  FILL_8755
timestamp 1677677812
transform 1 0 3272 0 1 1170
box -8 -3 16 105
use FILL  FILL_8756
timestamp 1677677812
transform 1 0 3280 0 1 1170
box -8 -3 16 105
use FILL  FILL_8757
timestamp 1677677812
transform 1 0 3288 0 1 1170
box -8 -3 16 105
use FILL  FILL_8758
timestamp 1677677812
transform 1 0 3296 0 1 1170
box -8 -3 16 105
use FILL  FILL_8760
timestamp 1677677812
transform 1 0 3304 0 1 1170
box -8 -3 16 105
use FILL  FILL_8762
timestamp 1677677812
transform 1 0 3312 0 1 1170
box -8 -3 16 105
use FILL  FILL_8764
timestamp 1677677812
transform 1 0 3320 0 1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_12
timestamp 1677677812
transform -1 0 3360 0 1 1170
box -7 -3 39 105
use FILL  FILL_8765
timestamp 1677677812
transform 1 0 3360 0 1 1170
box -8 -3 16 105
use FILL  FILL_8766
timestamp 1677677812
transform 1 0 3368 0 1 1170
box -8 -3 16 105
use FILL  FILL_8767
timestamp 1677677812
transform 1 0 3376 0 1 1170
box -8 -3 16 105
use FILL  FILL_8768
timestamp 1677677812
transform 1 0 3384 0 1 1170
box -8 -3 16 105
use FILL  FILL_8769
timestamp 1677677812
transform 1 0 3392 0 1 1170
box -8 -3 16 105
use FILL  FILL_8770
timestamp 1677677812
transform 1 0 3400 0 1 1170
box -8 -3 16 105
use FILL  FILL_8771
timestamp 1677677812
transform 1 0 3408 0 1 1170
box -8 -3 16 105
use FILL  FILL_8772
timestamp 1677677812
transform 1 0 3416 0 1 1170
box -8 -3 16 105
use FILL  FILL_8773
timestamp 1677677812
transform 1 0 3424 0 1 1170
box -8 -3 16 105
use FILL  FILL_8774
timestamp 1677677812
transform 1 0 3432 0 1 1170
box -8 -3 16 105
use FILL  FILL_8775
timestamp 1677677812
transform 1 0 3440 0 1 1170
box -8 -3 16 105
use FILL  FILL_8776
timestamp 1677677812
transform 1 0 3448 0 1 1170
box -8 -3 16 105
use FILL  FILL_8777
timestamp 1677677812
transform 1 0 3456 0 1 1170
box -8 -3 16 105
use FILL  FILL_8778
timestamp 1677677812
transform 1 0 3464 0 1 1170
box -8 -3 16 105
use FILL  FILL_8779
timestamp 1677677812
transform 1 0 3472 0 1 1170
box -8 -3 16 105
use FILL  FILL_8780
timestamp 1677677812
transform 1 0 3480 0 1 1170
box -8 -3 16 105
use FILL  FILL_8781
timestamp 1677677812
transform 1 0 3488 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_475
timestamp 1677677812
transform 1 0 3496 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_6645
timestamp 1677677812
transform 1 0 3604 0 1 1175
box -3 -3 3 3
use FILL  FILL_8782
timestamp 1677677812
transform 1 0 3592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8791
timestamp 1677677812
transform 1 0 3600 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_321
timestamp 1677677812
transform 1 0 3608 0 1 1170
box -8 -3 46 105
use FILL  FILL_8792
timestamp 1677677812
transform 1 0 3648 0 1 1170
box -8 -3 16 105
use FILL  FILL_8798
timestamp 1677677812
transform 1 0 3656 0 1 1170
box -8 -3 16 105
use FILL  FILL_8800
timestamp 1677677812
transform 1 0 3664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8802
timestamp 1677677812
transform 1 0 3672 0 1 1170
box -8 -3 16 105
use FILL  FILL_8804
timestamp 1677677812
transform 1 0 3680 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6646
timestamp 1677677812
transform 1 0 3708 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_322
timestamp 1677677812
transform 1 0 3688 0 1 1170
box -8 -3 46 105
use FILL  FILL_8806
timestamp 1677677812
transform 1 0 3728 0 1 1170
box -8 -3 16 105
use FILL  FILL_8813
timestamp 1677677812
transform 1 0 3736 0 1 1170
box -8 -3 16 105
use FILL  FILL_8815
timestamp 1677677812
transform 1 0 3744 0 1 1170
box -8 -3 16 105
use FILL  FILL_8817
timestamp 1677677812
transform 1 0 3752 0 1 1170
box -8 -3 16 105
use FILL  FILL_8819
timestamp 1677677812
transform 1 0 3760 0 1 1170
box -8 -3 16 105
use FILL  FILL_8821
timestamp 1677677812
transform 1 0 3768 0 1 1170
box -8 -3 16 105
use FILL  FILL_8822
timestamp 1677677812
transform 1 0 3776 0 1 1170
box -8 -3 16 105
use FILL  FILL_8823
timestamp 1677677812
transform 1 0 3784 0 1 1170
box -8 -3 16 105
use FILL  FILL_8824
timestamp 1677677812
transform 1 0 3792 0 1 1170
box -8 -3 16 105
use FILL  FILL_8825
timestamp 1677677812
transform 1 0 3800 0 1 1170
box -8 -3 16 105
use FILL  FILL_8826
timestamp 1677677812
transform 1 0 3808 0 1 1170
box -8 -3 16 105
use FILL  FILL_8828
timestamp 1677677812
transform 1 0 3816 0 1 1170
box -8 -3 16 105
use FILL  FILL_8830
timestamp 1677677812
transform 1 0 3824 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_556
timestamp 1677677812
transform -1 0 3848 0 1 1170
box -9 -3 26 105
use FILL  FILL_8831
timestamp 1677677812
transform 1 0 3848 0 1 1170
box -8 -3 16 105
use FILL  FILL_8832
timestamp 1677677812
transform 1 0 3856 0 1 1170
box -8 -3 16 105
use FILL  FILL_8833
timestamp 1677677812
transform 1 0 3864 0 1 1170
box -8 -3 16 105
use FILL  FILL_8835
timestamp 1677677812
transform 1 0 3872 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_476
timestamp 1677677812
transform 1 0 3880 0 1 1170
box -8 -3 104 105
use OAI22X1  OAI22X1_325
timestamp 1677677812
transform -1 0 4016 0 1 1170
box -8 -3 46 105
use FILL  FILL_8837
timestamp 1677677812
transform 1 0 4016 0 1 1170
box -8 -3 16 105
use FILL  FILL_8838
timestamp 1677677812
transform 1 0 4024 0 1 1170
box -8 -3 16 105
use FILL  FILL_8849
timestamp 1677677812
transform 1 0 4032 0 1 1170
box -8 -3 16 105
use FILL  FILL_8851
timestamp 1677677812
transform 1 0 4040 0 1 1170
box -8 -3 16 105
use FILL  FILL_8853
timestamp 1677677812
transform 1 0 4048 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6647
timestamp 1677677812
transform 1 0 4068 0 1 1175
box -3 -3 3 3
use INVX2  INVX2_559
timestamp 1677677812
transform -1 0 4072 0 1 1170
box -9 -3 26 105
use FILL  FILL_8854
timestamp 1677677812
transform 1 0 4072 0 1 1170
box -8 -3 16 105
use FILL  FILL_8855
timestamp 1677677812
transform 1 0 4080 0 1 1170
box -8 -3 16 105
use FILL  FILL_8856
timestamp 1677677812
transform 1 0 4088 0 1 1170
box -8 -3 16 105
use FILL  FILL_8857
timestamp 1677677812
transform 1 0 4096 0 1 1170
box -8 -3 16 105
use FILL  FILL_8858
timestamp 1677677812
transform 1 0 4104 0 1 1170
box -8 -3 16 105
use FILL  FILL_8862
timestamp 1677677812
transform 1 0 4112 0 1 1170
box -8 -3 16 105
use FILL  FILL_8864
timestamp 1677677812
transform 1 0 4120 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_477
timestamp 1677677812
transform 1 0 4128 0 1 1170
box -8 -3 104 105
use M3_M2  M3_M2_6648
timestamp 1677677812
transform 1 0 4284 0 1 1175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_478
timestamp 1677677812
transform 1 0 4224 0 1 1170
box -8 -3 104 105
use FILL  FILL_8866
timestamp 1677677812
transform 1 0 4320 0 1 1170
box -8 -3 16 105
use FILL  FILL_8883
timestamp 1677677812
transform 1 0 4328 0 1 1170
box -8 -3 16 105
use FILL  FILL_8885
timestamp 1677677812
transform 1 0 4336 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6649
timestamp 1677677812
transform 1 0 4380 0 1 1175
box -3 -3 3 3
use OAI22X1  OAI22X1_329
timestamp 1677677812
transform -1 0 4384 0 1 1170
box -8 -3 46 105
use FILL  FILL_8887
timestamp 1677677812
transform 1 0 4384 0 1 1170
box -8 -3 16 105
use FILL  FILL_8889
timestamp 1677677812
transform 1 0 4392 0 1 1170
box -8 -3 16 105
use FILL  FILL_8891
timestamp 1677677812
transform 1 0 4400 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6650
timestamp 1677677812
transform 1 0 4420 0 1 1175
box -3 -3 3 3
use FILL  FILL_8893
timestamp 1677677812
transform 1 0 4408 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_562
timestamp 1677677812
transform -1 0 4432 0 1 1170
box -9 -3 26 105
use FILL  FILL_8894
timestamp 1677677812
transform 1 0 4432 0 1 1170
box -8 -3 16 105
use FILL  FILL_8895
timestamp 1677677812
transform 1 0 4440 0 1 1170
box -8 -3 16 105
use FILL  FILL_8896
timestamp 1677677812
transform 1 0 4448 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_563
timestamp 1677677812
transform -1 0 4472 0 1 1170
box -9 -3 26 105
use FILL  FILL_8897
timestamp 1677677812
transform 1 0 4472 0 1 1170
box -8 -3 16 105
use FILL  FILL_8898
timestamp 1677677812
transform 1 0 4480 0 1 1170
box -8 -3 16 105
use FILL  FILL_8899
timestamp 1677677812
transform 1 0 4488 0 1 1170
box -8 -3 16 105
use FILL  FILL_8900
timestamp 1677677812
transform 1 0 4496 0 1 1170
box -8 -3 16 105
use FILL  FILL_8901
timestamp 1677677812
transform 1 0 4504 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_331
timestamp 1677677812
transform -1 0 4552 0 1 1170
box -8 -3 46 105
use FILL  FILL_8902
timestamp 1677677812
transform 1 0 4552 0 1 1170
box -8 -3 16 105
use FILL  FILL_8903
timestamp 1677677812
transform 1 0 4560 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_564
timestamp 1677677812
transform 1 0 4568 0 1 1170
box -9 -3 26 105
use FILL  FILL_8904
timestamp 1677677812
transform 1 0 4584 0 1 1170
box -8 -3 16 105
use FILL  FILL_8905
timestamp 1677677812
transform 1 0 4592 0 1 1170
box -8 -3 16 105
use FILL  FILL_8906
timestamp 1677677812
transform 1 0 4600 0 1 1170
box -8 -3 16 105
use FILL  FILL_8907
timestamp 1677677812
transform 1 0 4608 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_332
timestamp 1677677812
transform -1 0 4656 0 1 1170
box -8 -3 46 105
use FILL  FILL_8908
timestamp 1677677812
transform 1 0 4656 0 1 1170
box -8 -3 16 105
use FILL  FILL_8920
timestamp 1677677812
transform 1 0 4664 0 1 1170
box -8 -3 16 105
use FILL  FILL_8922
timestamp 1677677812
transform 1 0 4672 0 1 1170
box -8 -3 16 105
use FILL  FILL_8924
timestamp 1677677812
transform 1 0 4680 0 1 1170
box -8 -3 16 105
use FILL  FILL_8926
timestamp 1677677812
transform 1 0 4688 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6651
timestamp 1677677812
transform 1 0 4708 0 1 1175
box -3 -3 3 3
use FILL  FILL_8928
timestamp 1677677812
transform 1 0 4696 0 1 1170
box -8 -3 16 105
use FILL  FILL_8929
timestamp 1677677812
transform 1 0 4704 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_565
timestamp 1677677812
transform -1 0 4728 0 1 1170
box -9 -3 26 105
use FILL  FILL_8930
timestamp 1677677812
transform 1 0 4728 0 1 1170
box -8 -3 16 105
use FILL  FILL_8931
timestamp 1677677812
transform 1 0 4736 0 1 1170
box -8 -3 16 105
use FILL  FILL_8932
timestamp 1677677812
transform 1 0 4744 0 1 1170
box -8 -3 16 105
use FILL  FILL_8933
timestamp 1677677812
transform 1 0 4752 0 1 1170
box -8 -3 16 105
use FILL  FILL_8934
timestamp 1677677812
transform 1 0 4760 0 1 1170
box -8 -3 16 105
use FILL  FILL_8935
timestamp 1677677812
transform 1 0 4768 0 1 1170
box -8 -3 16 105
use FILL  FILL_8936
timestamp 1677677812
transform 1 0 4776 0 1 1170
box -8 -3 16 105
use FILL  FILL_8937
timestamp 1677677812
transform 1 0 4784 0 1 1170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_71
timestamp 1677677812
transform 1 0 4819 0 1 1170
box -10 -3 10 3
use M2_M1  M2_M1_7459
timestamp 1677677812
transform 1 0 100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7558
timestamp 1677677812
transform 1 0 108 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6760
timestamp 1677677812
transform 1 0 100 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7559
timestamp 1677677812
transform 1 0 148 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6652
timestamp 1677677812
transform 1 0 236 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7460
timestamp 1677677812
transform 1 0 204 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7461
timestamp 1677677812
transform 1 0 212 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7462
timestamp 1677677812
transform 1 0 228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7463
timestamp 1677677812
transform 1 0 236 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7560
timestamp 1677677812
transform 1 0 188 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6790
timestamp 1677677812
transform 1 0 180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6730
timestamp 1677677812
transform 1 0 196 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6731
timestamp 1677677812
transform 1 0 212 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7561
timestamp 1677677812
transform 1 0 220 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6761
timestamp 1677677812
transform 1 0 212 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6791
timestamp 1677677812
transform 1 0 228 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6686
timestamp 1677677812
transform 1 0 260 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7464
timestamp 1677677812
transform 1 0 252 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6687
timestamp 1677677812
transform 1 0 356 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7465
timestamp 1677677812
transform 1 0 356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7562
timestamp 1677677812
transform 1 0 268 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7563
timestamp 1677677812
transform 1 0 276 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7564
timestamp 1677677812
transform 1 0 308 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6762
timestamp 1677677812
transform 1 0 268 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6763
timestamp 1677677812
transform 1 0 308 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6792
timestamp 1677677812
transform 1 0 284 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7466
timestamp 1677677812
transform 1 0 396 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7467
timestamp 1677677812
transform 1 0 436 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6688
timestamp 1677677812
transform 1 0 460 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7468
timestamp 1677677812
transform 1 0 460 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7469
timestamp 1677677812
transform 1 0 476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7565
timestamp 1677677812
transform 1 0 452 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7566
timestamp 1677677812
transform 1 0 468 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6793
timestamp 1677677812
transform 1 0 468 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7567
timestamp 1677677812
transform 1 0 516 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6653
timestamp 1677677812
transform 1 0 588 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7568
timestamp 1677677812
transform 1 0 620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6794
timestamp 1677677812
transform 1 0 652 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6709
timestamp 1677677812
transform 1 0 676 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6838
timestamp 1677677812
transform 1 0 684 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6654
timestamp 1677677812
transform 1 0 700 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6655
timestamp 1677677812
transform 1 0 756 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7470
timestamp 1677677812
transform 1 0 700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7569
timestamp 1677677812
transform 1 0 748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7570
timestamp 1677677812
transform 1 0 780 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7571
timestamp 1677677812
transform 1 0 788 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6795
timestamp 1677677812
transform 1 0 748 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6732
timestamp 1677677812
transform 1 0 796 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6796
timestamp 1677677812
transform 1 0 788 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6826
timestamp 1677677812
transform 1 0 780 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6839
timestamp 1677677812
transform 1 0 708 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6668
timestamp 1677677812
transform 1 0 868 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7471
timestamp 1677677812
transform 1 0 836 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7472
timestamp 1677677812
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7473
timestamp 1677677812
transform 1 0 860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7572
timestamp 1677677812
transform 1 0 828 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6733
timestamp 1677677812
transform 1 0 836 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7451
timestamp 1677677812
transform 1 0 876 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6710
timestamp 1677677812
transform 1 0 876 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7573
timestamp 1677677812
transform 1 0 852 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7574
timestamp 1677677812
transform 1 0 868 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6797
timestamp 1677677812
transform 1 0 828 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6764
timestamp 1677677812
transform 1 0 868 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6798
timestamp 1677677812
transform 1 0 852 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6827
timestamp 1677677812
transform 1 0 844 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6734
timestamp 1677677812
transform 1 0 900 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6689
timestamp 1677677812
transform 1 0 916 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7452
timestamp 1677677812
transform 1 0 924 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7575
timestamp 1677677812
transform 1 0 908 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7474
timestamp 1677677812
transform 1 0 932 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7475
timestamp 1677677812
transform 1 0 948 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7576
timestamp 1677677812
transform 1 0 940 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6735
timestamp 1677677812
transform 1 0 948 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6690
timestamp 1677677812
transform 1 0 1052 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7476
timestamp 1677677812
transform 1 0 972 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6711
timestamp 1677677812
transform 1 0 1004 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6712
timestamp 1677677812
transform 1 0 1068 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7577
timestamp 1677677812
transform 1 0 956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7578
timestamp 1677677812
transform 1 0 1020 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7579
timestamp 1677677812
transform 1 0 1052 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7580
timestamp 1677677812
transform 1 0 1060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7581
timestamp 1677677812
transform 1 0 1068 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6799
timestamp 1677677812
transform 1 0 1020 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6800
timestamp 1677677812
transform 1 0 1068 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6828
timestamp 1677677812
transform 1 0 1052 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6840
timestamp 1677677812
transform 1 0 996 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6841
timestamp 1677677812
transform 1 0 1028 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7477
timestamp 1677677812
transform 1 0 1092 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6801
timestamp 1677677812
transform 1 0 1084 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6736
timestamp 1677677812
transform 1 0 1100 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6829
timestamp 1677677812
transform 1 0 1116 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7582
timestamp 1677677812
transform 1 0 1124 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6765
timestamp 1677677812
transform 1 0 1124 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6691
timestamp 1677677812
transform 1 0 1180 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7478
timestamp 1677677812
transform 1 0 1148 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6713
timestamp 1677677812
transform 1 0 1156 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7479
timestamp 1677677812
transform 1 0 1164 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6714
timestamp 1677677812
transform 1 0 1172 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7480
timestamp 1677677812
transform 1 0 1180 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6737
timestamp 1677677812
transform 1 0 1148 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6738
timestamp 1677677812
transform 1 0 1164 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7583
timestamp 1677677812
transform 1 0 1172 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7584
timestamp 1677677812
transform 1 0 1188 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6766
timestamp 1677677812
transform 1 0 1156 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6802
timestamp 1677677812
transform 1 0 1180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6692
timestamp 1677677812
transform 1 0 1308 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7481
timestamp 1677677812
transform 1 0 1308 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7585
timestamp 1677677812
transform 1 0 1324 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6693
timestamp 1677677812
transform 1 0 1356 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7482
timestamp 1677677812
transform 1 0 1348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7483
timestamp 1677677812
transform 1 0 1364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7586
timestamp 1677677812
transform 1 0 1340 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7587
timestamp 1677677812
transform 1 0 1356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7588
timestamp 1677677812
transform 1 0 1380 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7589
timestamp 1677677812
transform 1 0 1388 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6669
timestamp 1677677812
transform 1 0 1476 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7484
timestamp 1677677812
transform 1 0 1476 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7590
timestamp 1677677812
transform 1 0 1444 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6670
timestamp 1677677812
transform 1 0 1500 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7485
timestamp 1677677812
transform 1 0 1508 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6715
timestamp 1677677812
transform 1 0 1548 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6716
timestamp 1677677812
transform 1 0 1588 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7591
timestamp 1677677812
transform 1 0 1556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7592
timestamp 1677677812
transform 1 0 1588 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7593
timestamp 1677677812
transform 1 0 1596 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6803
timestamp 1677677812
transform 1 0 1540 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6804
timestamp 1677677812
transform 1 0 1596 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6671
timestamp 1677677812
transform 1 0 1628 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7486
timestamp 1677677812
transform 1 0 1628 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6717
timestamp 1677677812
transform 1 0 1636 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7487
timestamp 1677677812
transform 1 0 1644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7594
timestamp 1677677812
transform 1 0 1612 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6739
timestamp 1677677812
transform 1 0 1620 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7595
timestamp 1677677812
transform 1 0 1636 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6740
timestamp 1677677812
transform 1 0 1644 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6767
timestamp 1677677812
transform 1 0 1612 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6718
timestamp 1677677812
transform 1 0 1668 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7596
timestamp 1677677812
transform 1 0 1668 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6694
timestamp 1677677812
transform 1 0 1692 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7488
timestamp 1677677812
transform 1 0 1692 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6672
timestamp 1677677812
transform 1 0 1708 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7489
timestamp 1677677812
transform 1 0 1708 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7597
timestamp 1677677812
transform 1 0 1700 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6805
timestamp 1677677812
transform 1 0 1700 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6673
timestamp 1677677812
transform 1 0 1724 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6695
timestamp 1677677812
transform 1 0 1732 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_6719
timestamp 1677677812
transform 1 0 1748 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7490
timestamp 1677677812
transform 1 0 1756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7598
timestamp 1677677812
transform 1 0 1716 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7599
timestamp 1677677812
transform 1 0 1732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7600
timestamp 1677677812
transform 1 0 1748 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7601
timestamp 1677677812
transform 1 0 1756 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6830
timestamp 1677677812
transform 1 0 1716 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6806
timestamp 1677677812
transform 1 0 1756 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6674
timestamp 1677677812
transform 1 0 1772 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6741
timestamp 1677677812
transform 1 0 1804 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7491
timestamp 1677677812
transform 1 0 1828 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7602
timestamp 1677677812
transform 1 0 1836 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6696
timestamp 1677677812
transform 1 0 1980 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7492
timestamp 1677677812
transform 1 0 1908 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7493
timestamp 1677677812
transform 1 0 1916 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7494
timestamp 1677677812
transform 1 0 1940 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7495
timestamp 1677677812
transform 1 0 1956 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7496
timestamp 1677677812
transform 1 0 1964 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7497
timestamp 1677677812
transform 1 0 1972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7498
timestamp 1677677812
transform 1 0 1988 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7603
timestamp 1677677812
transform 1 0 1908 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6742
timestamp 1677677812
transform 1 0 1916 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7604
timestamp 1677677812
transform 1 0 1924 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7605
timestamp 1677677812
transform 1 0 1940 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7606
timestamp 1677677812
transform 1 0 1948 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6743
timestamp 1677677812
transform 1 0 1956 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7607
timestamp 1677677812
transform 1 0 1964 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7608
timestamp 1677677812
transform 1 0 1980 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7609
timestamp 1677677812
transform 1 0 1996 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6768
timestamp 1677677812
transform 1 0 1932 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6769
timestamp 1677677812
transform 1 0 1964 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6807
timestamp 1677677812
transform 1 0 1908 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6831
timestamp 1677677812
transform 1 0 1940 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6744
timestamp 1677677812
transform 1 0 2004 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6808
timestamp 1677677812
transform 1 0 1996 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6832
timestamp 1677677812
transform 1 0 1972 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6833
timestamp 1677677812
transform 1 0 2012 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_7610
timestamp 1677677812
transform 1 0 2028 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6842
timestamp 1677677812
transform 1 0 2036 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6697
timestamp 1677677812
transform 1 0 2052 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7499
timestamp 1677677812
transform 1 0 2044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7500
timestamp 1677677812
transform 1 0 2052 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6656
timestamp 1677677812
transform 1 0 2092 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6720
timestamp 1677677812
transform 1 0 2100 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7501
timestamp 1677677812
transform 1 0 2148 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7611
timestamp 1677677812
transform 1 0 2060 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7612
timestamp 1677677812
transform 1 0 2068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7613
timestamp 1677677812
transform 1 0 2100 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6770
timestamp 1677677812
transform 1 0 2060 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6771
timestamp 1677677812
transform 1 0 2100 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7614
timestamp 1677677812
transform 1 0 2180 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7667
timestamp 1677677812
transform 1 0 2164 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7680
timestamp 1677677812
transform 1 0 2172 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_6809
timestamp 1677677812
transform 1 0 2180 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6721
timestamp 1677677812
transform 1 0 2204 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6745
timestamp 1677677812
transform 1 0 2196 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7668
timestamp 1677677812
transform 1 0 2196 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7681
timestamp 1677677812
transform 1 0 2188 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_7682
timestamp 1677677812
transform 1 0 2196 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_6834
timestamp 1677677812
transform 1 0 2188 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6843
timestamp 1677677812
transform 1 0 2172 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6657
timestamp 1677677812
transform 1 0 2228 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7669
timestamp 1677677812
transform 1 0 2220 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6810
timestamp 1677677812
transform 1 0 2220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6835
timestamp 1677677812
transform 1 0 2220 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6844
timestamp 1677677812
transform 1 0 2212 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6746
timestamp 1677677812
transform 1 0 2252 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7683
timestamp 1677677812
transform 1 0 2252 0 1 1105
box -2 -2 2 2
use M2_M1  M2_M1_7670
timestamp 1677677812
transform 1 0 2284 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7615
timestamp 1677677812
transform 1 0 2332 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7671
timestamp 1677677812
transform 1 0 2324 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7502
timestamp 1677677812
transform 1 0 2372 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6836
timestamp 1677677812
transform 1 0 2372 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6658
timestamp 1677677812
transform 1 0 2396 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7453
timestamp 1677677812
transform 1 0 2492 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7616
timestamp 1677677812
transform 1 0 2396 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7617
timestamp 1677677812
transform 1 0 2404 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6747
timestamp 1677677812
transform 1 0 2436 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7503
timestamp 1677677812
transform 1 0 2508 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6811
timestamp 1677677812
transform 1 0 2452 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6812
timestamp 1677677812
transform 1 0 2476 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6813
timestamp 1677677812
transform 1 0 2500 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6698
timestamp 1677677812
transform 1 0 2516 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7504
timestamp 1677677812
transform 1 0 2516 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6837
timestamp 1677677812
transform 1 0 2508 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_6845
timestamp 1677677812
transform 1 0 2500 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7505
timestamp 1677677812
transform 1 0 2572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7618
timestamp 1677677812
transform 1 0 2540 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7619
timestamp 1677677812
transform 1 0 2556 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7620
timestamp 1677677812
transform 1 0 2564 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6772
timestamp 1677677812
transform 1 0 2532 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6773
timestamp 1677677812
transform 1 0 2564 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7506
timestamp 1677677812
transform 1 0 2604 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7507
timestamp 1677677812
transform 1 0 2620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7508
timestamp 1677677812
transform 1 0 2636 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7621
timestamp 1677677812
transform 1 0 2612 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7622
timestamp 1677677812
transform 1 0 2628 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6846
timestamp 1677677812
transform 1 0 2612 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6659
timestamp 1677677812
transform 1 0 2644 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7623
timestamp 1677677812
transform 1 0 2700 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6699
timestamp 1677677812
transform 1 0 2740 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7509
timestamp 1677677812
transform 1 0 2740 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6660
timestamp 1677677812
transform 1 0 2852 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7454
timestamp 1677677812
transform 1 0 2852 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6700
timestamp 1677677812
transform 1 0 2868 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7510
timestamp 1677677812
transform 1 0 2860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7511
timestamp 1677677812
transform 1 0 2868 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7624
timestamp 1677677812
transform 1 0 2756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7625
timestamp 1677677812
transform 1 0 2764 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6774
timestamp 1677677812
transform 1 0 2756 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6661
timestamp 1677677812
transform 1 0 3004 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6675
timestamp 1677677812
transform 1 0 2988 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7455
timestamp 1677677812
transform 1 0 2988 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6722
timestamp 1677677812
transform 1 0 2884 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7512
timestamp 1677677812
transform 1 0 2996 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7513
timestamp 1677677812
transform 1 0 3004 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7626
timestamp 1677677812
transform 1 0 2884 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7627
timestamp 1677677812
transform 1 0 2900 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6775
timestamp 1677677812
transform 1 0 2884 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6676
timestamp 1677677812
transform 1 0 3020 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7514
timestamp 1677677812
transform 1 0 3020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7628
timestamp 1677677812
transform 1 0 3028 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7672
timestamp 1677677812
transform 1 0 3020 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6814
timestamp 1677677812
transform 1 0 3028 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6701
timestamp 1677677812
transform 1 0 3044 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7515
timestamp 1677677812
transform 1 0 3044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7673
timestamp 1677677812
transform 1 0 3044 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7629
timestamp 1677677812
transform 1 0 3068 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7674
timestamp 1677677812
transform 1 0 3060 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6776
timestamp 1677677812
transform 1 0 3068 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6677
timestamp 1677677812
transform 1 0 3084 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7516
timestamp 1677677812
transform 1 0 3084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7517
timestamp 1677677812
transform 1 0 3108 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7630
timestamp 1677677812
transform 1 0 3084 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7631
timestamp 1677677812
transform 1 0 3100 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7675
timestamp 1677677812
transform 1 0 3084 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6815
timestamp 1677677812
transform 1 0 3084 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6748
timestamp 1677677812
transform 1 0 3108 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7632
timestamp 1677677812
transform 1 0 3124 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6678
timestamp 1677677812
transform 1 0 3148 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7456
timestamp 1677677812
transform 1 0 3148 0 1 1145
box -2 -2 2 2
use M2_M1  M2_M1_7676
timestamp 1677677812
transform 1 0 3164 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7633
timestamp 1677677812
transform 1 0 3180 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6679
timestamp 1677677812
transform 1 0 3220 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6723
timestamp 1677677812
transform 1 0 3212 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7518
timestamp 1677677812
transform 1 0 3220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7634
timestamp 1677677812
transform 1 0 3204 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6777
timestamp 1677677812
transform 1 0 3204 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7684
timestamp 1677677812
transform 1 0 3196 0 1 1105
box -2 -2 2 2
use M3_M2  M3_M2_6778
timestamp 1677677812
transform 1 0 3220 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7677
timestamp 1677677812
transform 1 0 3228 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6816
timestamp 1677677812
transform 1 0 3228 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7519
timestamp 1677677812
transform 1 0 3284 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7635
timestamp 1677677812
transform 1 0 3260 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7636
timestamp 1677677812
transform 1 0 3276 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6817
timestamp 1677677812
transform 1 0 3276 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7520
timestamp 1677677812
transform 1 0 3300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7521
timestamp 1677677812
transform 1 0 3308 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6779
timestamp 1677677812
transform 1 0 3308 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6680
timestamp 1677677812
transform 1 0 3332 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6724
timestamp 1677677812
transform 1 0 3324 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7522
timestamp 1677677812
transform 1 0 3356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7637
timestamp 1677677812
transform 1 0 3324 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7638
timestamp 1677677812
transform 1 0 3332 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6749
timestamp 1677677812
transform 1 0 3340 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7639
timestamp 1677677812
transform 1 0 3348 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6681
timestamp 1677677812
transform 1 0 3492 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6702
timestamp 1677677812
transform 1 0 3380 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7457
timestamp 1677677812
transform 1 0 3388 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6703
timestamp 1677677812
transform 1 0 3476 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7523
timestamp 1677677812
transform 1 0 3380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7640
timestamp 1677677812
transform 1 0 3372 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6780
timestamp 1677677812
transform 1 0 3372 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6725
timestamp 1677677812
transform 1 0 3388 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7524
timestamp 1677677812
transform 1 0 3492 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7525
timestamp 1677677812
transform 1 0 3500 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7641
timestamp 1677677812
transform 1 0 3476 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7642
timestamp 1677677812
transform 1 0 3484 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6781
timestamp 1677677812
transform 1 0 3484 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6726
timestamp 1677677812
transform 1 0 3508 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_6750
timestamp 1677677812
transform 1 0 3508 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6751
timestamp 1677677812
transform 1 0 3548 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7678
timestamp 1677677812
transform 1 0 3564 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_6818
timestamp 1677677812
transform 1 0 3564 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7526
timestamp 1677677812
transform 1 0 3588 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7527
timestamp 1677677812
transform 1 0 3596 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7643
timestamp 1677677812
transform 1 0 3604 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7644
timestamp 1677677812
transform 1 0 3620 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6819
timestamp 1677677812
transform 1 0 3628 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6847
timestamp 1677677812
transform 1 0 3636 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6820
timestamp 1677677812
transform 1 0 3668 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7528
timestamp 1677677812
transform 1 0 3684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7645
timestamp 1677677812
transform 1 0 3748 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6848
timestamp 1677677812
transform 1 0 3764 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7529
timestamp 1677677812
transform 1 0 3788 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7646
timestamp 1677677812
transform 1 0 3796 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7530
timestamp 1677677812
transform 1 0 3812 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6752
timestamp 1677677812
transform 1 0 3812 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6704
timestamp 1677677812
transform 1 0 3860 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7531
timestamp 1677677812
transform 1 0 3828 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7532
timestamp 1677677812
transform 1 0 3844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7533
timestamp 1677677812
transform 1 0 3860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7647
timestamp 1677677812
transform 1 0 3820 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6782
timestamp 1677677812
transform 1 0 3820 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7648
timestamp 1677677812
transform 1 0 3852 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6849
timestamp 1677677812
transform 1 0 3828 0 1 1085
box -3 -3 3 3
use M2_M1  M2_M1_7649
timestamp 1677677812
transform 1 0 3868 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6783
timestamp 1677677812
transform 1 0 3868 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6662
timestamp 1677677812
transform 1 0 3908 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6705
timestamp 1677677812
transform 1 0 3908 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7534
timestamp 1677677812
transform 1 0 3900 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7535
timestamp 1677677812
transform 1 0 3908 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6753
timestamp 1677677812
transform 1 0 3900 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6706
timestamp 1677677812
transform 1 0 3972 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7536
timestamp 1677677812
transform 1 0 3956 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7537
timestamp 1677677812
transform 1 0 3972 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7650
timestamp 1677677812
transform 1 0 3948 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6754
timestamp 1677677812
transform 1 0 3972 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6784
timestamp 1677677812
transform 1 0 3948 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6850
timestamp 1677677812
transform 1 0 3972 0 1 1085
box -3 -3 3 3
use M3_M2  M3_M2_6785
timestamp 1677677812
transform 1 0 3988 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6707
timestamp 1677677812
transform 1 0 4020 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7538
timestamp 1677677812
transform 1 0 4020 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7651
timestamp 1677677812
transform 1 0 4012 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6663
timestamp 1677677812
transform 1 0 4036 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7539
timestamp 1677677812
transform 1 0 4036 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6664
timestamp 1677677812
transform 1 0 4084 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7540
timestamp 1677677812
transform 1 0 4084 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7541
timestamp 1677677812
transform 1 0 4100 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7652
timestamp 1677677812
transform 1 0 4076 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7653
timestamp 1677677812
transform 1 0 4092 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6755
timestamp 1677677812
transform 1 0 4100 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6821
timestamp 1677677812
transform 1 0 4076 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_6665
timestamp 1677677812
transform 1 0 4164 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7654
timestamp 1677677812
transform 1 0 4164 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7458
timestamp 1677677812
transform 1 0 4220 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_6727
timestamp 1677677812
transform 1 0 4220 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7542
timestamp 1677677812
transform 1 0 4228 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7655
timestamp 1677677812
transform 1 0 4228 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6786
timestamp 1677677812
transform 1 0 4228 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_7543
timestamp 1677677812
transform 1 0 4260 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7656
timestamp 1677677812
transform 1 0 4268 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6822
timestamp 1677677812
transform 1 0 4268 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7657
timestamp 1677677812
transform 1 0 4284 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6787
timestamp 1677677812
transform 1 0 4284 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6682
timestamp 1677677812
transform 1 0 4300 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7544
timestamp 1677677812
transform 1 0 4300 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6823
timestamp 1677677812
transform 1 0 4300 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7545
timestamp 1677677812
transform 1 0 4316 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6756
timestamp 1677677812
transform 1 0 4324 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6683
timestamp 1677677812
transform 1 0 4332 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7546
timestamp 1677677812
transform 1 0 4332 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7547
timestamp 1677677812
transform 1 0 4348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7548
timestamp 1677677812
transform 1 0 4364 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7658
timestamp 1677677812
transform 1 0 4332 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6757
timestamp 1677677812
transform 1 0 4340 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6728
timestamp 1677677812
transform 1 0 4372 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7549
timestamp 1677677812
transform 1 0 4380 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7659
timestamp 1677677812
transform 1 0 4356 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7660
timestamp 1677677812
transform 1 0 4372 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6788
timestamp 1677677812
transform 1 0 4364 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6824
timestamp 1677677812
transform 1 0 4348 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7550
timestamp 1677677812
transform 1 0 4420 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7661
timestamp 1677677812
transform 1 0 4444 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7662
timestamp 1677677812
transform 1 0 4500 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6789
timestamp 1677677812
transform 1 0 4444 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_6666
timestamp 1677677812
transform 1 0 4540 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_7551
timestamp 1677677812
transform 1 0 4532 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7552
timestamp 1677677812
transform 1 0 4548 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7663
timestamp 1677677812
transform 1 0 4540 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6667
timestamp 1677677812
transform 1 0 4580 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_6684
timestamp 1677677812
transform 1 0 4580 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_7553
timestamp 1677677812
transform 1 0 4580 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7664
timestamp 1677677812
transform 1 0 4580 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_6708
timestamp 1677677812
transform 1 0 4588 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_7554
timestamp 1677677812
transform 1 0 4588 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6758
timestamp 1677677812
transform 1 0 4588 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_6759
timestamp 1677677812
transform 1 0 4604 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_7679
timestamp 1677677812
transform 1 0 4588 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_7555
timestamp 1677677812
transform 1 0 4620 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_7556
timestamp 1677677812
transform 1 0 4636 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6685
timestamp 1677677812
transform 1 0 4652 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_6825
timestamp 1677677812
transform 1 0 4692 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_7557
timestamp 1677677812
transform 1 0 4708 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_6729
timestamp 1677677812
transform 1 0 4772 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_7665
timestamp 1677677812
transform 1 0 4756 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_7666
timestamp 1677677812
transform 1 0 4788 0 1 1125
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_72
timestamp 1677677812
transform 1 0 24 0 1 1070
box -10 -3 10 3
use FILL  FILL_8447
timestamp 1677677812
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8449
timestamp 1677677812
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8451
timestamp 1677677812
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_531
timestamp 1677677812
transform 1 0 96 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8465
timestamp 1677677812
transform 1 0 112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8466
timestamp 1677677812
transform 1 0 120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8467
timestamp 1677677812
transform 1 0 128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8468
timestamp 1677677812
transform 1 0 136 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_532
timestamp 1677677812
transform -1 0 160 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8469
timestamp 1677677812
transform 1 0 160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8470
timestamp 1677677812
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8471
timestamp 1677677812
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8472
timestamp 1677677812
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8473
timestamp 1677677812
transform 1 0 192 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_312
timestamp 1677677812
transform -1 0 240 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8474
timestamp 1677677812
transform 1 0 240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8475
timestamp 1677677812
transform 1 0 248 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_533
timestamp 1677677812
transform 1 0 256 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_459
timestamp 1677677812
transform -1 0 368 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8476
timestamp 1677677812
transform 1 0 368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8479
timestamp 1677677812
transform 1 0 376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8480
timestamp 1677677812
transform 1 0 384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8481
timestamp 1677677812
transform 1 0 392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8482
timestamp 1677677812
transform 1 0 400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8483
timestamp 1677677812
transform 1 0 408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8484
timestamp 1677677812
transform 1 0 416 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8485
timestamp 1677677812
transform 1 0 424 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8493
timestamp 1677677812
transform 1 0 432 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_316
timestamp 1677677812
transform -1 0 480 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8494
timestamp 1677677812
transform 1 0 480 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8495
timestamp 1677677812
transform 1 0 488 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8496
timestamp 1677677812
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8497
timestamp 1677677812
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8498
timestamp 1677677812
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8499
timestamp 1677677812
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8500
timestamp 1677677812
transform 1 0 528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8501
timestamp 1677677812
transform 1 0 536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8502
timestamp 1677677812
transform 1 0 544 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_535
timestamp 1677677812
transform -1 0 568 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8503
timestamp 1677677812
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8504
timestamp 1677677812
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8505
timestamp 1677677812
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8506
timestamp 1677677812
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8508
timestamp 1677677812
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8510
timestamp 1677677812
transform 1 0 608 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8511
timestamp 1677677812
transform 1 0 616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8512
timestamp 1677677812
transform 1 0 624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8513
timestamp 1677677812
transform 1 0 632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8514
timestamp 1677677812
transform 1 0 640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8515
timestamp 1677677812
transform 1 0 648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8517
timestamp 1677677812
transform 1 0 656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8526
timestamp 1677677812
transform 1 0 664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8527
timestamp 1677677812
transform 1 0 672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8528
timestamp 1677677812
transform 1 0 680 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_461
timestamp 1677677812
transform 1 0 688 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8529
timestamp 1677677812
transform 1 0 784 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8540
timestamp 1677677812
transform 1 0 792 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_537
timestamp 1677677812
transform -1 0 816 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8541
timestamp 1677677812
transform 1 0 816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8542
timestamp 1677677812
transform 1 0 824 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_316
timestamp 1677677812
transform -1 0 872 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8543
timestamp 1677677812
transform 1 0 872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8544
timestamp 1677677812
transform 1 0 880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8545
timestamp 1677677812
transform 1 0 888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8546
timestamp 1677677812
transform 1 0 896 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_86
timestamp 1677677812
transform 1 0 904 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8547
timestamp 1677677812
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6851
timestamp 1677677812
transform 1 0 956 0 1 1075
box -3 -3 3 3
use NOR2X1  NOR2X1_87
timestamp 1677677812
transform 1 0 936 0 -1 1170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_464
timestamp 1677677812
transform 1 0 960 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_538
timestamp 1677677812
transform -1 0 1072 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8548
timestamp 1677677812
transform 1 0 1072 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8549
timestamp 1677677812
transform 1 0 1080 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8550
timestamp 1677677812
transform 1 0 1088 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_539
timestamp 1677677812
transform -1 0 1112 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8551
timestamp 1677677812
transform 1 0 1112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8553
timestamp 1677677812
transform 1 0 1120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8560
timestamp 1677677812
transform 1 0 1128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8561
timestamp 1677677812
transform 1 0 1136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8562
timestamp 1677677812
transform 1 0 1144 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_317
timestamp 1677677812
transform 1 0 1152 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8563
timestamp 1677677812
transform 1 0 1192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8565
timestamp 1677677812
transform 1 0 1200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8567
timestamp 1677677812
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8569
timestamp 1677677812
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8571
timestamp 1677677812
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8574
timestamp 1677677812
transform 1 0 1232 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8575
timestamp 1677677812
transform 1 0 1240 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8576
timestamp 1677677812
transform 1 0 1248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8577
timestamp 1677677812
transform 1 0 1256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8578
timestamp 1677677812
transform 1 0 1264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8579
timestamp 1677677812
transform 1 0 1272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8580
timestamp 1677677812
transform 1 0 1280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8582
timestamp 1677677812
transform 1 0 1288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8584
timestamp 1677677812
transform 1 0 1296 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_542
timestamp 1677677812
transform 1 0 1304 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8595
timestamp 1677677812
transform 1 0 1320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8596
timestamp 1677677812
transform 1 0 1328 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_320
timestamp 1677677812
transform -1 0 1376 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8597
timestamp 1677677812
transform 1 0 1376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8598
timestamp 1677677812
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_465
timestamp 1677677812
transform -1 0 1488 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8599
timestamp 1677677812
transform 1 0 1488 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_466
timestamp 1677677812
transform 1 0 1496 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8606
timestamp 1677677812
transform 1 0 1592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8608
timestamp 1677677812
transform 1 0 1600 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8611
timestamp 1677677812
transform 1 0 1608 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_321
timestamp 1677677812
transform 1 0 1616 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8612
timestamp 1677677812
transform 1 0 1656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8618
timestamp 1677677812
transform 1 0 1664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8619
timestamp 1677677812
transform 1 0 1672 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_6852
timestamp 1677677812
transform 1 0 1692 0 1 1075
box -3 -3 3 3
use FILL  FILL_8620
timestamp 1677677812
transform 1 0 1680 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_545
timestamp 1677677812
transform 1 0 1688 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8621
timestamp 1677677812
transform 1 0 1704 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_322
timestamp 1677677812
transform 1 0 1712 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8622
timestamp 1677677812
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8623
timestamp 1677677812
transform 1 0 1760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8624
timestamp 1677677812
transform 1 0 1768 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_546
timestamp 1677677812
transform -1 0 1792 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8625
timestamp 1677677812
transform 1 0 1792 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8626
timestamp 1677677812
transform 1 0 1800 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8627
timestamp 1677677812
transform 1 0 1808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8628
timestamp 1677677812
transform 1 0 1816 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8629
timestamp 1677677812
transform 1 0 1824 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_547
timestamp 1677677812
transform -1 0 1848 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8630
timestamp 1677677812
transform 1 0 1848 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8631
timestamp 1677677812
transform 1 0 1856 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8632
timestamp 1677677812
transform 1 0 1864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8633
timestamp 1677677812
transform 1 0 1872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8634
timestamp 1677677812
transform 1 0 1880 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8635
timestamp 1677677812
transform 1 0 1888 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8636
timestamp 1677677812
transform 1 0 1896 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_323
timestamp 1677677812
transform -1 0 1944 0 -1 1170
box -8 -3 46 105
use INVX2  INVX2_548
timestamp 1677677812
transform -1 0 1960 0 -1 1170
box -9 -3 26 105
use AOI22X1  AOI22X1_324
timestamp 1677677812
transform 1 0 1960 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8637
timestamp 1677677812
transform 1 0 2000 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8639
timestamp 1677677812
transform 1 0 2008 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8641
timestamp 1677677812
transform 1 0 2016 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8652
timestamp 1677677812
transform 1 0 2024 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_549
timestamp 1677677812
transform -1 0 2048 0 -1 1170
box -9 -3 26 105
use INVX2  INVX2_550
timestamp 1677677812
transform 1 0 2048 0 -1 1170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_471
timestamp 1677677812
transform -1 0 2160 0 -1 1170
box -8 -3 104 105
use NAND3X1  NAND3X1_65
timestamp 1677677812
transform -1 0 2192 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8653
timestamp 1677677812
transform 1 0 2192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8655
timestamp 1677677812
transform 1 0 2200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8657
timestamp 1677677812
transform 1 0 2208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8658
timestamp 1677677812
transform 1 0 2216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8659
timestamp 1677677812
transform 1 0 2224 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_66
timestamp 1677677812
transform 1 0 2232 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8660
timestamp 1677677812
transform 1 0 2264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8661
timestamp 1677677812
transform 1 0 2272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8662
timestamp 1677677812
transform 1 0 2280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8663
timestamp 1677677812
transform 1 0 2288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8664
timestamp 1677677812
transform 1 0 2296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8665
timestamp 1677677812
transform 1 0 2304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8666
timestamp 1677677812
transform 1 0 2312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8667
timestamp 1677677812
transform 1 0 2320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8668
timestamp 1677677812
transform 1 0 2328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8671
timestamp 1677677812
transform 1 0 2336 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_18
timestamp 1677677812
transform -1 0 2368 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8672
timestamp 1677677812
transform 1 0 2368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8673
timestamp 1677677812
transform 1 0 2376 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_12
timestamp 1677677812
transform 1 0 2384 0 -1 1170
box -5 -3 126 105
use FILL  FILL_8703
timestamp 1677677812
transform 1 0 2504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8704
timestamp 1677677812
transform 1 0 2512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8705
timestamp 1677677812
transform 1 0 2520 0 -1 1170
box -8 -3 16 105
use AND2X2  AND2X2_52
timestamp 1677677812
transform 1 0 2528 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8706
timestamp 1677677812
transform 1 0 2560 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8707
timestamp 1677677812
transform 1 0 2568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8708
timestamp 1677677812
transform 1 0 2576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8709
timestamp 1677677812
transform 1 0 2584 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_326
timestamp 1677677812
transform 1 0 2592 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8710
timestamp 1677677812
transform 1 0 2632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8711
timestamp 1677677812
transform 1 0 2640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8712
timestamp 1677677812
transform 1 0 2648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8713
timestamp 1677677812
transform 1 0 2656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8714
timestamp 1677677812
transform 1 0 2664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8715
timestamp 1677677812
transform 1 0 2672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8716
timestamp 1677677812
transform 1 0 2680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8717
timestamp 1677677812
transform 1 0 2688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8718
timestamp 1677677812
transform 1 0 2696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8719
timestamp 1677677812
transform 1 0 2704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8720
timestamp 1677677812
transform 1 0 2712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8721
timestamp 1677677812
transform 1 0 2720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8722
timestamp 1677677812
transform 1 0 2728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8723
timestamp 1677677812
transform 1 0 2736 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_13
timestamp 1677677812
transform 1 0 2744 0 -1 1170
box -5 -3 126 105
use FILL  FILL_8724
timestamp 1677677812
transform 1 0 2864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8725
timestamp 1677677812
transform 1 0 2872 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_14
timestamp 1677677812
transform 1 0 2880 0 -1 1170
box -5 -3 126 105
use NAND2X1  NAND2X1_20
timestamp 1677677812
transform 1 0 3000 0 -1 1170
box -8 -3 32 105
use NAND2X1  NAND2X1_21
timestamp 1677677812
transform 1 0 3024 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8726
timestamp 1677677812
transform 1 0 3048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8727
timestamp 1677677812
transform 1 0 3056 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_553
timestamp 1677677812
transform 1 0 3064 0 -1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_152
timestamp 1677677812
transform -1 0 3112 0 -1 1170
box -8 -3 34 105
use FILL  FILL_8728
timestamp 1677677812
transform 1 0 3112 0 -1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_11
timestamp 1677677812
transform 1 0 3120 0 -1 1170
box -7 -3 39 105
use FILL  FILL_8734
timestamp 1677677812
transform 1 0 3152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8736
timestamp 1677677812
transform 1 0 3160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8738
timestamp 1677677812
transform 1 0 3168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8745
timestamp 1677677812
transform 1 0 3176 0 -1 1170
box -8 -3 16 105
use NAND3X1  NAND3X1_68
timestamp 1677677812
transform -1 0 3216 0 -1 1170
box -8 -3 40 105
use FILL  FILL_8746
timestamp 1677677812
transform 1 0 3216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8748
timestamp 1677677812
transform 1 0 3224 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_554
timestamp 1677677812
transform 1 0 3232 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8752
timestamp 1677677812
transform 1 0 3248 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_327
timestamp 1677677812
transform 1 0 3256 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8759
timestamp 1677677812
transform 1 0 3296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8761
timestamp 1677677812
transform 1 0 3304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8763
timestamp 1677677812
transform 1 0 3312 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8783
timestamp 1677677812
transform 1 0 3320 0 -1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_328
timestamp 1677677812
transform -1 0 3368 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8784
timestamp 1677677812
transform 1 0 3368 0 -1 1170
box -8 -3 16 105
use FAX1  FAX1_15
timestamp 1677677812
transform -1 0 3496 0 -1 1170
box -5 -3 126 105
use NAND2X1  NAND2X1_22
timestamp 1677677812
transform 1 0 3496 0 -1 1170
box -8 -3 32 105
use FILL  FILL_8785
timestamp 1677677812
transform 1 0 3520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8786
timestamp 1677677812
transform 1 0 3528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8787
timestamp 1677677812
transform 1 0 3536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8788
timestamp 1677677812
transform 1 0 3544 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8789
timestamp 1677677812
transform 1 0 3552 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_153
timestamp 1677677812
transform -1 0 3592 0 -1 1170
box -8 -3 34 105
use FILL  FILL_8790
timestamp 1677677812
transform 1 0 3592 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_555
timestamp 1677677812
transform 1 0 3600 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8793
timestamp 1677677812
transform 1 0 3616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8794
timestamp 1677677812
transform 1 0 3624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8795
timestamp 1677677812
transform 1 0 3632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8796
timestamp 1677677812
transform 1 0 3640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8797
timestamp 1677677812
transform 1 0 3648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8799
timestamp 1677677812
transform 1 0 3656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8801
timestamp 1677677812
transform 1 0 3664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8803
timestamp 1677677812
transform 1 0 3672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8805
timestamp 1677677812
transform 1 0 3680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8807
timestamp 1677677812
transform 1 0 3688 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8808
timestamp 1677677812
transform 1 0 3696 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8809
timestamp 1677677812
transform 1 0 3704 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8810
timestamp 1677677812
transform 1 0 3712 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8811
timestamp 1677677812
transform 1 0 3720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8812
timestamp 1677677812
transform 1 0 3728 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8814
timestamp 1677677812
transform 1 0 3736 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8816
timestamp 1677677812
transform 1 0 3744 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8818
timestamp 1677677812
transform 1 0 3752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8820
timestamp 1677677812
transform 1 0 3760 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_323
timestamp 1677677812
transform 1 0 3768 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8827
timestamp 1677677812
transform 1 0 3808 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8829
timestamp 1677677812
transform 1 0 3816 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_324
timestamp 1677677812
transform 1 0 3824 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8834
timestamp 1677677812
transform 1 0 3864 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8836
timestamp 1677677812
transform 1 0 3872 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8839
timestamp 1677677812
transform 1 0 3880 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_557
timestamp 1677677812
transform -1 0 3904 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8840
timestamp 1677677812
transform 1 0 3904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8841
timestamp 1677677812
transform 1 0 3912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8842
timestamp 1677677812
transform 1 0 3920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8843
timestamp 1677677812
transform 1 0 3928 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_326
timestamp 1677677812
transform -1 0 3976 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8844
timestamp 1677677812
transform 1 0 3976 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8845
timestamp 1677677812
transform 1 0 3984 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8846
timestamp 1677677812
transform 1 0 3992 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8847
timestamp 1677677812
transform 1 0 4000 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_558
timestamp 1677677812
transform -1 0 4024 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8848
timestamp 1677677812
transform 1 0 4024 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8850
timestamp 1677677812
transform 1 0 4032 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8852
timestamp 1677677812
transform 1 0 4040 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8859
timestamp 1677677812
transform 1 0 4048 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8860
timestamp 1677677812
transform 1 0 4056 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_327
timestamp 1677677812
transform -1 0 4104 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8861
timestamp 1677677812
transform 1 0 4104 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8863
timestamp 1677677812
transform 1 0 4112 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8865
timestamp 1677677812
transform 1 0 4120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8867
timestamp 1677677812
transform 1 0 4128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8868
timestamp 1677677812
transform 1 0 4136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8869
timestamp 1677677812
transform 1 0 4144 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8870
timestamp 1677677812
transform 1 0 4152 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_560
timestamp 1677677812
transform -1 0 4176 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8871
timestamp 1677677812
transform 1 0 4176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8872
timestamp 1677677812
transform 1 0 4184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8873
timestamp 1677677812
transform 1 0 4192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8874
timestamp 1677677812
transform 1 0 4200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8875
timestamp 1677677812
transform 1 0 4208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8876
timestamp 1677677812
transform 1 0 4216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8877
timestamp 1677677812
transform 1 0 4224 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8878
timestamp 1677677812
transform 1 0 4232 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_328
timestamp 1677677812
transform 1 0 4240 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8879
timestamp 1677677812
transform 1 0 4280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8880
timestamp 1677677812
transform 1 0 4288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8881
timestamp 1677677812
transform 1 0 4296 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_561
timestamp 1677677812
transform -1 0 4320 0 -1 1170
box -9 -3 26 105
use FILL  FILL_8882
timestamp 1677677812
transform 1 0 4320 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8884
timestamp 1677677812
transform 1 0 4328 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8886
timestamp 1677677812
transform 1 0 4336 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_330
timestamp 1677677812
transform -1 0 4384 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8888
timestamp 1677677812
transform 1 0 4384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8890
timestamp 1677677812
transform 1 0 4392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8892
timestamp 1677677812
transform 1 0 4400 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_479
timestamp 1677677812
transform 1 0 4408 0 -1 1170
box -8 -3 104 105
use FILL  FILL_8909
timestamp 1677677812
transform 1 0 4504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8910
timestamp 1677677812
transform 1 0 4512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8911
timestamp 1677677812
transform 1 0 4520 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_333
timestamp 1677677812
transform -1 0 4568 0 -1 1170
box -8 -3 46 105
use FILL  FILL_8912
timestamp 1677677812
transform 1 0 4568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8913
timestamp 1677677812
transform 1 0 4576 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_154
timestamp 1677677812
transform -1 0 4616 0 -1 1170
box -8 -3 34 105
use FILL  FILL_8914
timestamp 1677677812
transform 1 0 4616 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8915
timestamp 1677677812
transform 1 0 4624 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8916
timestamp 1677677812
transform 1 0 4632 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8917
timestamp 1677677812
transform 1 0 4640 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8918
timestamp 1677677812
transform 1 0 4648 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8919
timestamp 1677677812
transform 1 0 4656 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8921
timestamp 1677677812
transform 1 0 4664 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8923
timestamp 1677677812
transform 1 0 4672 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8925
timestamp 1677677812
transform 1 0 4680 0 -1 1170
box -8 -3 16 105
use FILL  FILL_8927
timestamp 1677677812
transform 1 0 4688 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_480
timestamp 1677677812
transform 1 0 4696 0 -1 1170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_73
timestamp 1677677812
transform 1 0 4843 0 1 1070
box -10 -3 10 3
use M2_M1  M2_M1_7694
timestamp 1677677812
transform 1 0 108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7823
timestamp 1677677812
transform 1 0 84 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6920
timestamp 1677677812
transform 1 0 172 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6921
timestamp 1677677812
transform 1 0 228 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7695
timestamp 1677677812
transform 1 0 196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7696
timestamp 1677677812
transform 1 0 212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7697
timestamp 1677677812
transform 1 0 228 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6984
timestamp 1677677812
transform 1 0 196 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7824
timestamp 1677677812
transform 1 0 204 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7825
timestamp 1677677812
transform 1 0 220 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7826
timestamp 1677677812
transform 1 0 228 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7009
timestamp 1677677812
transform 1 0 204 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6895
timestamp 1677677812
transform 1 0 252 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6922
timestamp 1677677812
transform 1 0 244 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6923
timestamp 1677677812
transform 1 0 260 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7698
timestamp 1677677812
transform 1 0 252 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6985
timestamp 1677677812
transform 1 0 244 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7699
timestamp 1677677812
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7827
timestamp 1677677812
transform 1 0 260 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7828
timestamp 1677677812
transform 1 0 276 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7050
timestamp 1677677812
transform 1 0 220 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7051
timestamp 1677677812
transform 1 0 236 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7010
timestamp 1677677812
transform 1 0 276 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7052
timestamp 1677677812
transform 1 0 252 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6858
timestamp 1677677812
transform 1 0 300 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6859
timestamp 1677677812
transform 1 0 356 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6924
timestamp 1677677812
transform 1 0 388 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7700
timestamp 1677677812
transform 1 0 348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7701
timestamp 1677677812
transform 1 0 380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7702
timestamp 1677677812
transform 1 0 388 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7829
timestamp 1677677812
transform 1 0 300 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6986
timestamp 1677677812
transform 1 0 348 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6964
timestamp 1677677812
transform 1 0 396 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6925
timestamp 1677677812
transform 1 0 428 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7703
timestamp 1677677812
transform 1 0 404 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7704
timestamp 1677677812
transform 1 0 420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7830
timestamp 1677677812
transform 1 0 396 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7831
timestamp 1677677812
transform 1 0 412 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6987
timestamp 1677677812
transform 1 0 420 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7053
timestamp 1677677812
transform 1 0 412 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6896
timestamp 1677677812
transform 1 0 452 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7705
timestamp 1677677812
transform 1 0 460 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6965
timestamp 1677677812
transform 1 0 476 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7706
timestamp 1677677812
transform 1 0 516 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7832
timestamp 1677677812
transform 1 0 452 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7833
timestamp 1677677812
transform 1 0 476 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7011
timestamp 1677677812
transform 1 0 476 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7012
timestamp 1677677812
transform 1 0 500 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7054
timestamp 1677677812
transform 1 0 452 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6926
timestamp 1677677812
transform 1 0 612 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7707
timestamp 1677677812
transform 1 0 596 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7708
timestamp 1677677812
transform 1 0 604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7834
timestamp 1677677812
transform 1 0 580 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7835
timestamp 1677677812
transform 1 0 588 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7013
timestamp 1677677812
transform 1 0 596 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7055
timestamp 1677677812
transform 1 0 588 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6966
timestamp 1677677812
transform 1 0 612 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7709
timestamp 1677677812
transform 1 0 620 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7710
timestamp 1677677812
transform 1 0 636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7836
timestamp 1677677812
transform 1 0 628 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7014
timestamp 1677677812
transform 1 0 628 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7711
timestamp 1677677812
transform 1 0 652 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6897
timestamp 1677677812
transform 1 0 668 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6898
timestamp 1677677812
transform 1 0 684 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7712
timestamp 1677677812
transform 1 0 684 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6988
timestamp 1677677812
transform 1 0 660 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7837
timestamp 1677677812
transform 1 0 676 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6989
timestamp 1677677812
transform 1 0 684 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6853
timestamp 1677677812
transform 1 0 708 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_7056
timestamp 1677677812
transform 1 0 700 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6927
timestamp 1677677812
transform 1 0 788 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7713
timestamp 1677677812
transform 1 0 732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7714
timestamp 1677677812
transform 1 0 788 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6990
timestamp 1677677812
transform 1 0 772 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7838
timestamp 1677677812
transform 1 0 812 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7015
timestamp 1677677812
transform 1 0 732 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7057
timestamp 1677677812
transform 1 0 732 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7058
timestamp 1677677812
transform 1 0 812 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6928
timestamp 1677677812
transform 1 0 828 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7715
timestamp 1677677812
transform 1 0 828 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7059
timestamp 1677677812
transform 1 0 836 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7716
timestamp 1677677812
transform 1 0 852 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7717
timestamp 1677677812
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6967
timestamp 1677677812
transform 1 0 876 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6875
timestamp 1677677812
transform 1 0 916 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6929
timestamp 1677677812
transform 1 0 916 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6968
timestamp 1677677812
transform 1 0 892 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7718
timestamp 1677677812
transform 1 0 900 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7719
timestamp 1677677812
transform 1 0 916 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7839
timestamp 1677677812
transform 1 0 876 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7840
timestamp 1677677812
transform 1 0 884 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6991
timestamp 1677677812
transform 1 0 892 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7841
timestamp 1677677812
transform 1 0 908 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7016
timestamp 1677677812
transform 1 0 884 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7060
timestamp 1677677812
transform 1 0 900 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6969
timestamp 1677677812
transform 1 0 940 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7842
timestamp 1677677812
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6930
timestamp 1677677812
transform 1 0 1012 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7720
timestamp 1677677812
transform 1 0 1012 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7843
timestamp 1677677812
transform 1 0 964 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7017
timestamp 1677677812
transform 1 0 964 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7018
timestamp 1677677812
transform 1 0 996 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6931
timestamp 1677677812
transform 1 0 1060 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6876
timestamp 1677677812
transform 1 0 1092 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7721
timestamp 1677677812
transform 1 0 1084 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7722
timestamp 1677677812
transform 1 0 1092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7723
timestamp 1677677812
transform 1 0 1108 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7019
timestamp 1677677812
transform 1 0 1084 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7844
timestamp 1677677812
transform 1 0 1100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7845
timestamp 1677677812
transform 1 0 1124 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7020
timestamp 1677677812
transform 1 0 1124 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7931
timestamp 1677677812
transform 1 0 1132 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_7061
timestamp 1677677812
transform 1 0 1116 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6932
timestamp 1677677812
transform 1 0 1148 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7724
timestamp 1677677812
transform 1 0 1148 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7846
timestamp 1677677812
transform 1 0 1140 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6933
timestamp 1677677812
transform 1 0 1188 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7847
timestamp 1677677812
transform 1 0 1188 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7021
timestamp 1677677812
transform 1 0 1188 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7725
timestamp 1677677812
transform 1 0 1220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7726
timestamp 1677677812
transform 1 0 1236 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6970
timestamp 1677677812
transform 1 0 1244 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7727
timestamp 1677677812
transform 1 0 1260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7848
timestamp 1677677812
transform 1 0 1244 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7849
timestamp 1677677812
transform 1 0 1348 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6877
timestamp 1677677812
transform 1 0 1364 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7728
timestamp 1677677812
transform 1 0 1380 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7850
timestamp 1677677812
transform 1 0 1380 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7851
timestamp 1677677812
transform 1 0 1388 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7062
timestamp 1677677812
transform 1 0 1388 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7729
timestamp 1677677812
transform 1 0 1420 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7730
timestamp 1677677812
transform 1 0 1436 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7731
timestamp 1677677812
transform 1 0 1444 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7852
timestamp 1677677812
transform 1 0 1436 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6860
timestamp 1677677812
transform 1 0 1556 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7732
timestamp 1677677812
transform 1 0 1524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7853
timestamp 1677677812
transform 1 0 1556 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6861
timestamp 1677677812
transform 1 0 1580 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7733
timestamp 1677677812
transform 1 0 1572 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6899
timestamp 1677677812
transform 1 0 1644 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7734
timestamp 1677677812
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7735
timestamp 1677677812
transform 1 0 1644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7854
timestamp 1677677812
transform 1 0 1660 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6934
timestamp 1677677812
transform 1 0 1676 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7736
timestamp 1677677812
transform 1 0 1700 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7855
timestamp 1677677812
transform 1 0 1676 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7856
timestamp 1677677812
transform 1 0 1692 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7063
timestamp 1677677812
transform 1 0 1676 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6971
timestamp 1677677812
transform 1 0 1716 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6862
timestamp 1677677812
transform 1 0 1780 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7737
timestamp 1677677812
transform 1 0 1748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7738
timestamp 1677677812
transform 1 0 1764 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6972
timestamp 1677677812
transform 1 0 1772 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7739
timestamp 1677677812
transform 1 0 1780 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7857
timestamp 1677677812
transform 1 0 1748 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7858
timestamp 1677677812
transform 1 0 1772 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7859
timestamp 1677677812
transform 1 0 1780 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6935
timestamp 1677677812
transform 1 0 1836 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6936
timestamp 1677677812
transform 1 0 1892 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7740
timestamp 1677677812
transform 1 0 1828 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7741
timestamp 1677677812
transform 1 0 1836 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7742
timestamp 1677677812
transform 1 0 1892 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7860
timestamp 1677677812
transform 1 0 1916 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7022
timestamp 1677677812
transform 1 0 1916 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6973
timestamp 1677677812
transform 1 0 1932 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7861
timestamp 1677677812
transform 1 0 1932 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6937
timestamp 1677677812
transform 1 0 1948 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7743
timestamp 1677677812
transform 1 0 1972 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6863
timestamp 1677677812
transform 1 0 2020 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6878
timestamp 1677677812
transform 1 0 2028 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7744
timestamp 1677677812
transform 1 0 1988 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7745
timestamp 1677677812
transform 1 0 2004 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7746
timestamp 1677677812
transform 1 0 2020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7862
timestamp 1677677812
transform 1 0 2012 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7023
timestamp 1677677812
transform 1 0 1996 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7747
timestamp 1677677812
transform 1 0 2036 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6864
timestamp 1677677812
transform 1 0 2060 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6879
timestamp 1677677812
transform 1 0 2108 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7748
timestamp 1677677812
transform 1 0 2100 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7863
timestamp 1677677812
transform 1 0 2124 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6865
timestamp 1677677812
transform 1 0 2148 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6880
timestamp 1677677812
transform 1 0 2148 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6900
timestamp 1677677812
transform 1 0 2140 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7686
timestamp 1677677812
transform 1 0 2140 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6854
timestamp 1677677812
transform 1 0 2164 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6881
timestamp 1677677812
transform 1 0 2164 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7685
timestamp 1677677812
transform 1 0 2172 0 1 1035
box -2 -2 2 2
use M3_M2  M3_M2_6901
timestamp 1677677812
transform 1 0 2180 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7687
timestamp 1677677812
transform 1 0 2180 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7749
timestamp 1677677812
transform 1 0 2180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7750
timestamp 1677677812
transform 1 0 2196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7864
timestamp 1677677812
transform 1 0 2196 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7024
timestamp 1677677812
transform 1 0 2196 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7064
timestamp 1677677812
transform 1 0 2196 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6866
timestamp 1677677812
transform 1 0 2212 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6902
timestamp 1677677812
transform 1 0 2268 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6938
timestamp 1677677812
transform 1 0 2276 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7751
timestamp 1677677812
transform 1 0 2220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7752
timestamp 1677677812
transform 1 0 2276 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7865
timestamp 1677677812
transform 1 0 2300 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7025
timestamp 1677677812
transform 1 0 2220 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7065
timestamp 1677677812
transform 1 0 2252 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6939
timestamp 1677677812
transform 1 0 2316 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7866
timestamp 1677677812
transform 1 0 2316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7688
timestamp 1677677812
transform 1 0 2332 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6882
timestamp 1677677812
transform 1 0 2356 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6867
timestamp 1677677812
transform 1 0 2380 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7753
timestamp 1677677812
transform 1 0 2348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7754
timestamp 1677677812
transform 1 0 2356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7755
timestamp 1677677812
transform 1 0 2372 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7867
timestamp 1677677812
transform 1 0 2356 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6992
timestamp 1677677812
transform 1 0 2364 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7026
timestamp 1677677812
transform 1 0 2356 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7027
timestamp 1677677812
transform 1 0 2404 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7756
timestamp 1677677812
transform 1 0 2436 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6993
timestamp 1677677812
transform 1 0 2436 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6994
timestamp 1677677812
transform 1 0 2452 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7757
timestamp 1677677812
transform 1 0 2476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7758
timestamp 1677677812
transform 1 0 2484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7868
timestamp 1677677812
transform 1 0 2468 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7869
timestamp 1677677812
transform 1 0 2476 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7932
timestamp 1677677812
transform 1 0 2452 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_6995
timestamp 1677677812
transform 1 0 2484 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6940
timestamp 1677677812
transform 1 0 2564 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7759
timestamp 1677677812
transform 1 0 2532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7760
timestamp 1677677812
transform 1 0 2556 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7870
timestamp 1677677812
transform 1 0 2500 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7871
timestamp 1677677812
transform 1 0 2508 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7872
timestamp 1677677812
transform 1 0 2556 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7066
timestamp 1677677812
transform 1 0 2524 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6883
timestamp 1677677812
transform 1 0 2604 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6941
timestamp 1677677812
transform 1 0 2604 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6884
timestamp 1677677812
transform 1 0 2644 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6885
timestamp 1677677812
transform 1 0 2684 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7761
timestamp 1677677812
transform 1 0 2604 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7762
timestamp 1677677812
transform 1 0 2628 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7763
timestamp 1677677812
transform 1 0 2684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7873
timestamp 1677677812
transform 1 0 2572 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7028
timestamp 1677677812
transform 1 0 2572 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7874
timestamp 1677677812
transform 1 0 2620 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6996
timestamp 1677677812
transform 1 0 2628 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7875
timestamp 1677677812
transform 1 0 2708 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7067
timestamp 1677677812
transform 1 0 2692 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7764
timestamp 1677677812
transform 1 0 2732 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7876
timestamp 1677677812
transform 1 0 2724 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7029
timestamp 1677677812
transform 1 0 2724 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7068
timestamp 1677677812
transform 1 0 2732 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6868
timestamp 1677677812
transform 1 0 2860 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6869
timestamp 1677677812
transform 1 0 2876 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6903
timestamp 1677677812
transform 1 0 2764 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6904
timestamp 1677677812
transform 1 0 2852 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6942
timestamp 1677677812
transform 1 0 2748 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7765
timestamp 1677677812
transform 1 0 2748 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7766
timestamp 1677677812
transform 1 0 2756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7877
timestamp 1677677812
transform 1 0 2852 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7933
timestamp 1677677812
transform 1 0 2844 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_6886
timestamp 1677677812
transform 1 0 2868 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6905
timestamp 1677677812
transform 1 0 2868 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6906
timestamp 1677677812
transform 1 0 2900 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6943
timestamp 1677677812
transform 1 0 2972 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7767
timestamp 1677677812
transform 1 0 2964 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7768
timestamp 1677677812
transform 1 0 2972 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7878
timestamp 1677677812
transform 1 0 2868 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7879
timestamp 1677677812
transform 1 0 2980 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7880
timestamp 1677677812
transform 1 0 2988 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7934
timestamp 1677677812
transform 1 0 2876 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_7069
timestamp 1677677812
transform 1 0 2876 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6907
timestamp 1677677812
transform 1 0 3028 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7689
timestamp 1677677812
transform 1 0 3020 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7769
timestamp 1677677812
transform 1 0 3028 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7881
timestamp 1677677812
transform 1 0 3020 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7070
timestamp 1677677812
transform 1 0 3020 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6908
timestamp 1677677812
transform 1 0 3052 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7690
timestamp 1677677812
transform 1 0 3044 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7691
timestamp 1677677812
transform 1 0 3052 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7770
timestamp 1677677812
transform 1 0 3060 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7882
timestamp 1677677812
transform 1 0 3068 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7030
timestamp 1677677812
transform 1 0 3060 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7071
timestamp 1677677812
transform 1 0 3068 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6944
timestamp 1677677812
transform 1 0 3092 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6945
timestamp 1677677812
transform 1 0 3116 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7771
timestamp 1677677812
transform 1 0 3092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7772
timestamp 1677677812
transform 1 0 3100 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6974
timestamp 1677677812
transform 1 0 3108 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7773
timestamp 1677677812
transform 1 0 3124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7883
timestamp 1677677812
transform 1 0 3100 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6997
timestamp 1677677812
transform 1 0 3108 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7884
timestamp 1677677812
transform 1 0 3116 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7935
timestamp 1677677812
transform 1 0 3100 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_7072
timestamp 1677677812
transform 1 0 3100 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6909
timestamp 1677677812
transform 1 0 3180 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6975
timestamp 1677677812
transform 1 0 3172 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7774
timestamp 1677677812
transform 1 0 3180 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7885
timestamp 1677677812
transform 1 0 3188 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7031
timestamp 1677677812
transform 1 0 3180 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7775
timestamp 1677677812
transform 1 0 3212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7776
timestamp 1677677812
transform 1 0 3228 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7886
timestamp 1677677812
transform 1 0 3220 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6998
timestamp 1677677812
transform 1 0 3228 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7887
timestamp 1677677812
transform 1 0 3244 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7032
timestamp 1677677812
transform 1 0 3212 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6910
timestamp 1677677812
transform 1 0 3260 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7777
timestamp 1677677812
transform 1 0 3260 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7778
timestamp 1677677812
transform 1 0 3276 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6946
timestamp 1677677812
transform 1 0 3300 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7779
timestamp 1677677812
transform 1 0 3308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7888
timestamp 1677677812
transform 1 0 3300 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7889
timestamp 1677677812
transform 1 0 3316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7890
timestamp 1677677812
transform 1 0 3324 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6911
timestamp 1677677812
transform 1 0 3356 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7780
timestamp 1677677812
transform 1 0 3348 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7781
timestamp 1677677812
transform 1 0 3356 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7782
timestamp 1677677812
transform 1 0 3372 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6999
timestamp 1677677812
transform 1 0 3348 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7000
timestamp 1677677812
transform 1 0 3460 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7936
timestamp 1677677812
transform 1 0 3460 0 1 995
box -2 -2 2 2
use M2_M1  M2_M1_7783
timestamp 1677677812
transform 1 0 3476 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6887
timestamp 1677677812
transform 1 0 3492 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6947
timestamp 1677677812
transform 1 0 3484 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7784
timestamp 1677677812
transform 1 0 3484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7891
timestamp 1677677812
transform 1 0 3484 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7033
timestamp 1677677812
transform 1 0 3484 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7892
timestamp 1677677812
transform 1 0 3508 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6948
timestamp 1677677812
transform 1 0 3540 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7785
timestamp 1677677812
transform 1 0 3532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7786
timestamp 1677677812
transform 1 0 3548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7893
timestamp 1677677812
transform 1 0 3548 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7034
timestamp 1677677812
transform 1 0 3548 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7787
timestamp 1677677812
transform 1 0 3564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7788
timestamp 1677677812
transform 1 0 3580 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7035
timestamp 1677677812
transform 1 0 3572 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7789
timestamp 1677677812
transform 1 0 3620 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7073
timestamp 1677677812
transform 1 0 3612 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6912
timestamp 1677677812
transform 1 0 3644 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6870
timestamp 1677677812
transform 1 0 3684 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6913
timestamp 1677677812
transform 1 0 3668 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6949
timestamp 1677677812
transform 1 0 3660 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7790
timestamp 1677677812
transform 1 0 3660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7791
timestamp 1677677812
transform 1 0 3668 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7792
timestamp 1677677812
transform 1 0 3684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7894
timestamp 1677677812
transform 1 0 3676 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7074
timestamp 1677677812
transform 1 0 3676 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6871
timestamp 1677677812
transform 1 0 3716 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6855
timestamp 1677677812
transform 1 0 3748 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6950
timestamp 1677677812
transform 1 0 3740 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6951
timestamp 1677677812
transform 1 0 3764 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6976
timestamp 1677677812
transform 1 0 3732 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7793
timestamp 1677677812
transform 1 0 3748 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6977
timestamp 1677677812
transform 1 0 3756 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7794
timestamp 1677677812
transform 1 0 3764 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7895
timestamp 1677677812
transform 1 0 3732 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7896
timestamp 1677677812
transform 1 0 3740 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7001
timestamp 1677677812
transform 1 0 3748 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6888
timestamp 1677677812
transform 1 0 3780 0 1 1045
box -3 -3 3 3
use M2_M1  M2_M1_7897
timestamp 1677677812
transform 1 0 3756 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7898
timestamp 1677677812
transform 1 0 3772 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7036
timestamp 1677677812
transform 1 0 3740 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7075
timestamp 1677677812
transform 1 0 3732 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7076
timestamp 1677677812
transform 1 0 3772 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6889
timestamp 1677677812
transform 1 0 3796 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6952
timestamp 1677677812
transform 1 0 3796 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7002
timestamp 1677677812
transform 1 0 3796 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7037
timestamp 1677677812
transform 1 0 3788 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7795
timestamp 1677677812
transform 1 0 3812 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6978
timestamp 1677677812
transform 1 0 3828 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7796
timestamp 1677677812
transform 1 0 3844 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7003
timestamp 1677677812
transform 1 0 3852 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7899
timestamp 1677677812
transform 1 0 3892 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7077
timestamp 1677677812
transform 1 0 3820 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6914
timestamp 1677677812
transform 1 0 3908 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7797
timestamp 1677677812
transform 1 0 3908 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6872
timestamp 1677677812
transform 1 0 3956 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6953
timestamp 1677677812
transform 1 0 3964 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7798
timestamp 1677677812
transform 1 0 3956 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7900
timestamp 1677677812
transform 1 0 3932 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7901
timestamp 1677677812
transform 1 0 3948 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7038
timestamp 1677677812
transform 1 0 3932 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6856
timestamp 1677677812
transform 1 0 4036 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6890
timestamp 1677677812
transform 1 0 4020 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6954
timestamp 1677677812
transform 1 0 4028 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7799
timestamp 1677677812
transform 1 0 4020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7800
timestamp 1677677812
transform 1 0 4036 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7902
timestamp 1677677812
transform 1 0 4012 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7903
timestamp 1677677812
transform 1 0 4028 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7904
timestamp 1677677812
transform 1 0 4044 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7039
timestamp 1677677812
transform 1 0 4044 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7004
timestamp 1677677812
transform 1 0 4060 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6873
timestamp 1677677812
transform 1 0 4092 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_6915
timestamp 1677677812
transform 1 0 4108 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7801
timestamp 1677677812
transform 1 0 4092 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7802
timestamp 1677677812
transform 1 0 4108 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7803
timestamp 1677677812
transform 1 0 4116 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7905
timestamp 1677677812
transform 1 0 4084 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7906
timestamp 1677677812
transform 1 0 4100 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7005
timestamp 1677677812
transform 1 0 4108 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7907
timestamp 1677677812
transform 1 0 4148 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7040
timestamp 1677677812
transform 1 0 4148 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6857
timestamp 1677677812
transform 1 0 4188 0 1 1065
box -3 -3 3 3
use M3_M2  M3_M2_6891
timestamp 1677677812
transform 1 0 4172 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6916
timestamp 1677677812
transform 1 0 4196 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6955
timestamp 1677677812
transform 1 0 4188 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7804
timestamp 1677677812
transform 1 0 4172 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7805
timestamp 1677677812
transform 1 0 4188 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7806
timestamp 1677677812
transform 1 0 4196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7908
timestamp 1677677812
transform 1 0 4164 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7909
timestamp 1677677812
transform 1 0 4180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7910
timestamp 1677677812
transform 1 0 4196 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7041
timestamp 1677677812
transform 1 0 4196 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_6874
timestamp 1677677812
transform 1 0 4252 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_7807
timestamp 1677677812
transform 1 0 4252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7911
timestamp 1677677812
transform 1 0 4228 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7912
timestamp 1677677812
transform 1 0 4244 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7042
timestamp 1677677812
transform 1 0 4252 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7913
timestamp 1677677812
transform 1 0 4292 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6892
timestamp 1677677812
transform 1 0 4308 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6956
timestamp 1677677812
transform 1 0 4324 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7808
timestamp 1677677812
transform 1 0 4308 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7809
timestamp 1677677812
transform 1 0 4324 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7914
timestamp 1677677812
transform 1 0 4316 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7915
timestamp 1677677812
transform 1 0 4332 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7078
timestamp 1677677812
transform 1 0 4308 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6917
timestamp 1677677812
transform 1 0 4348 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_7810
timestamp 1677677812
transform 1 0 4348 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6918
timestamp 1677677812
transform 1 0 4396 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6957
timestamp 1677677812
transform 1 0 4372 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6979
timestamp 1677677812
transform 1 0 4388 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7811
timestamp 1677677812
transform 1 0 4396 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7916
timestamp 1677677812
transform 1 0 4372 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7006
timestamp 1677677812
transform 1 0 4380 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_6919
timestamp 1677677812
transform 1 0 4420 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_6958
timestamp 1677677812
transform 1 0 4412 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7812
timestamp 1677677812
transform 1 0 4412 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7917
timestamp 1677677812
transform 1 0 4388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7918
timestamp 1677677812
transform 1 0 4404 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7043
timestamp 1677677812
transform 1 0 4396 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7919
timestamp 1677677812
transform 1 0 4436 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6959
timestamp 1677677812
transform 1 0 4444 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_7044
timestamp 1677677812
transform 1 0 4452 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7079
timestamp 1677677812
transform 1 0 4444 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7692
timestamp 1677677812
transform 1 0 4468 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_7813
timestamp 1677677812
transform 1 0 4468 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7080
timestamp 1677677812
transform 1 0 4460 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_7814
timestamp 1677677812
transform 1 0 4484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7920
timestamp 1677677812
transform 1 0 4492 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7693
timestamp 1677677812
transform 1 0 4500 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_6980
timestamp 1677677812
transform 1 0 4500 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_6981
timestamp 1677677812
transform 1 0 4516 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_7007
timestamp 1677677812
transform 1 0 4508 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_7045
timestamp 1677677812
transform 1 0 4500 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7081
timestamp 1677677812
transform 1 0 4508 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6960
timestamp 1677677812
transform 1 0 4540 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7921
timestamp 1677677812
transform 1 0 4532 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_6961
timestamp 1677677812
transform 1 0 4564 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_7815
timestamp 1677677812
transform 1 0 4548 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_6982
timestamp 1677677812
transform 1 0 4556 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7816
timestamp 1677677812
transform 1 0 4564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7817
timestamp 1677677812
transform 1 0 4580 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7922
timestamp 1677677812
transform 1 0 4556 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7008
timestamp 1677677812
transform 1 0 4564 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_7923
timestamp 1677677812
transform 1 0 4572 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7818
timestamp 1677677812
transform 1 0 4596 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_7082
timestamp 1677677812
transform 1 0 4612 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_6962
timestamp 1677677812
transform 1 0 4628 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6893
timestamp 1677677812
transform 1 0 4644 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6894
timestamp 1677677812
transform 1 0 4676 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_6963
timestamp 1677677812
transform 1 0 4660 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_6983
timestamp 1677677812
transform 1 0 4652 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_7819
timestamp 1677677812
transform 1 0 4660 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7820
timestamp 1677677812
transform 1 0 4676 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7924
timestamp 1677677812
transform 1 0 4644 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7925
timestamp 1677677812
transform 1 0 4652 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7926
timestamp 1677677812
transform 1 0 4668 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7927
timestamp 1677677812
transform 1 0 4684 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_7928
timestamp 1677677812
transform 1 0 4692 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7046
timestamp 1677677812
transform 1 0 4644 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_7083
timestamp 1677677812
transform 1 0 4644 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_7047
timestamp 1677677812
transform 1 0 4684 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7821
timestamp 1677677812
transform 1 0 4740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7822
timestamp 1677677812
transform 1 0 4756 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_7929
timestamp 1677677812
transform 1 0 4748 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7048
timestamp 1677677812
transform 1 0 4756 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_7930
timestamp 1677677812
transform 1 0 4772 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_7049
timestamp 1677677812
transform 1 0 4796 0 1 995
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_74
timestamp 1677677812
transform 1 0 48 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_7084
timestamp 1677677812
transform 1 0 68 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7085
timestamp 1677677812
transform 1 0 92 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_481
timestamp 1677677812
transform 1 0 72 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_7086
timestamp 1677677812
transform 1 0 180 0 1 975
box -3 -3 3 3
use FILL  FILL_8938
timestamp 1677677812
transform 1 0 168 0 1 970
box -8 -3 16 105
use FILL  FILL_8939
timestamp 1677677812
transform 1 0 176 0 1 970
box -8 -3 16 105
use FILL  FILL_8940
timestamp 1677677812
transform 1 0 184 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7087
timestamp 1677677812
transform 1 0 212 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_329
timestamp 1677677812
transform -1 0 232 0 1 970
box -8 -3 46 105
use FILL  FILL_8941
timestamp 1677677812
transform 1 0 232 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7088
timestamp 1677677812
transform 1 0 260 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_334
timestamp 1677677812
transform -1 0 280 0 1 970
box -8 -3 46 105
use FILL  FILL_8942
timestamp 1677677812
transform 1 0 280 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_482
timestamp 1677677812
transform 1 0 288 0 1 970
box -8 -3 104 105
use AOI22X1  AOI22X1_330
timestamp 1677677812
transform -1 0 424 0 1 970
box -8 -3 46 105
use FILL  FILL_8943
timestamp 1677677812
transform 1 0 424 0 1 970
box -8 -3 16 105
use FILL  FILL_8952
timestamp 1677677812
transform 1 0 432 0 1 970
box -8 -3 16 105
use FILL  FILL_8953
timestamp 1677677812
transform 1 0 440 0 1 970
box -8 -3 16 105
use INVX2  INVX2_570
timestamp 1677677812
transform 1 0 448 0 1 970
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_485
timestamp 1677677812
transform 1 0 464 0 1 970
box -8 -3 104 105
use FILL  FILL_8954
timestamp 1677677812
transform 1 0 560 0 1 970
box -8 -3 16 105
use FILL  FILL_8960
timestamp 1677677812
transform 1 0 568 0 1 970
box -8 -3 16 105
use FILL  FILL_8961
timestamp 1677677812
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_8962
timestamp 1677677812
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_8963
timestamp 1677677812
transform 1 0 592 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_332
timestamp 1677677812
transform 1 0 600 0 1 970
box -8 -3 46 105
use FILL  FILL_8964
timestamp 1677677812
transform 1 0 640 0 1 970
box -8 -3 16 105
use FILL  FILL_8965
timestamp 1677677812
transform 1 0 648 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_335
timestamp 1677677812
transform 1 0 656 0 1 970
box -8 -3 46 105
use FILL  FILL_8966
timestamp 1677677812
transform 1 0 696 0 1 970
box -8 -3 16 105
use FILL  FILL_8974
timestamp 1677677812
transform 1 0 704 0 1 970
box -8 -3 16 105
use FILL  FILL_8976
timestamp 1677677812
transform 1 0 712 0 1 970
box -8 -3 16 105
use FILL  FILL_8978
timestamp 1677677812
transform 1 0 720 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_487
timestamp 1677677812
transform -1 0 824 0 1 970
box -8 -3 104 105
use FILL  FILL_8979
timestamp 1677677812
transform 1 0 824 0 1 970
box -8 -3 16 105
use FILL  FILL_8982
timestamp 1677677812
transform 1 0 832 0 1 970
box -8 -3 16 105
use INVX2  INVX2_571
timestamp 1677677812
transform -1 0 856 0 1 970
box -9 -3 26 105
use FILL  FILL_8984
timestamp 1677677812
transform 1 0 856 0 1 970
box -8 -3 16 105
use FILL  FILL_8986
timestamp 1677677812
transform 1 0 864 0 1 970
box -8 -3 16 105
use FILL  FILL_8988
timestamp 1677677812
transform 1 0 872 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_334
timestamp 1677677812
transform -1 0 920 0 1 970
box -8 -3 46 105
use FILL  FILL_8989
timestamp 1677677812
transform 1 0 920 0 1 970
box -8 -3 16 105
use FILL  FILL_8990
timestamp 1677677812
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_8991
timestamp 1677677812
transform 1 0 936 0 1 970
box -8 -3 16 105
use FILL  FILL_8996
timestamp 1677677812
transform 1 0 944 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_489
timestamp 1677677812
transform 1 0 952 0 1 970
box -8 -3 104 105
use FILL  FILL_8998
timestamp 1677677812
transform 1 0 1048 0 1 970
box -8 -3 16 105
use FILL  FILL_8999
timestamp 1677677812
transform 1 0 1056 0 1 970
box -8 -3 16 105
use FILL  FILL_9000
timestamp 1677677812
transform 1 0 1064 0 1 970
box -8 -3 16 105
use FILL  FILL_9001
timestamp 1677677812
transform 1 0 1072 0 1 970
box -8 -3 16 105
use FILL  FILL_9013
timestamp 1677677812
transform 1 0 1080 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7089
timestamp 1677677812
transform 1 0 1132 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_336
timestamp 1677677812
transform 1 0 1088 0 1 970
box -8 -3 46 105
use FILL  FILL_9015
timestamp 1677677812
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_9016
timestamp 1677677812
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_9017
timestamp 1677677812
transform 1 0 1144 0 1 970
box -8 -3 16 105
use FILL  FILL_9018
timestamp 1677677812
transform 1 0 1152 0 1 970
box -8 -3 16 105
use FILL  FILL_9023
timestamp 1677677812
transform 1 0 1160 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_90
timestamp 1677677812
transform 1 0 1168 0 1 970
box -8 -3 32 105
use FILL  FILL_9025
timestamp 1677677812
transform 1 0 1192 0 1 970
box -8 -3 16 105
use FILL  FILL_9027
timestamp 1677677812
transform 1 0 1200 0 1 970
box -8 -3 16 105
use FILL  FILL_9029
timestamp 1677677812
transform 1 0 1208 0 1 970
box -8 -3 16 105
use FILL  FILL_9030
timestamp 1677677812
transform 1 0 1216 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_337
timestamp 1677677812
transform -1 0 1264 0 1 970
box -8 -3 46 105
use FILL  FILL_9031
timestamp 1677677812
transform 1 0 1264 0 1 970
box -8 -3 16 105
use FILL  FILL_9035
timestamp 1677677812
transform 1 0 1272 0 1 970
box -8 -3 16 105
use FILL  FILL_9037
timestamp 1677677812
transform 1 0 1280 0 1 970
box -8 -3 16 105
use FILL  FILL_9039
timestamp 1677677812
transform 1 0 1288 0 1 970
box -8 -3 16 105
use FILL  FILL_9040
timestamp 1677677812
transform 1 0 1296 0 1 970
box -8 -3 16 105
use FILL  FILL_9041
timestamp 1677677812
transform 1 0 1304 0 1 970
box -8 -3 16 105
use FILL  FILL_9042
timestamp 1677677812
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_9043
timestamp 1677677812
transform 1 0 1320 0 1 970
box -8 -3 16 105
use FILL  FILL_9044
timestamp 1677677812
transform 1 0 1328 0 1 970
box -8 -3 16 105
use FILL  FILL_9045
timestamp 1677677812
transform 1 0 1336 0 1 970
box -8 -3 16 105
use FILL  FILL_9046
timestamp 1677677812
transform 1 0 1344 0 1 970
box -8 -3 16 105
use FILL  FILL_9047
timestamp 1677677812
transform 1 0 1352 0 1 970
box -8 -3 16 105
use FILL  FILL_9048
timestamp 1677677812
transform 1 0 1360 0 1 970
box -8 -3 16 105
use FILL  FILL_9049
timestamp 1677677812
transform 1 0 1368 0 1 970
box -8 -3 16 105
use FILL  FILL_9050
timestamp 1677677812
transform 1 0 1376 0 1 970
box -8 -3 16 105
use FILL  FILL_9051
timestamp 1677677812
transform 1 0 1384 0 1 970
box -8 -3 16 105
use FILL  FILL_9052
timestamp 1677677812
transform 1 0 1392 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_338
timestamp 1677677812
transform 1 0 1400 0 1 970
box -8 -3 46 105
use FILL  FILL_9053
timestamp 1677677812
transform 1 0 1440 0 1 970
box -8 -3 16 105
use FILL  FILL_9054
timestamp 1677677812
transform 1 0 1448 0 1 970
box -8 -3 16 105
use FILL  FILL_9057
timestamp 1677677812
transform 1 0 1456 0 1 970
box -8 -3 16 105
use FILL  FILL_9059
timestamp 1677677812
transform 1 0 1464 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_491
timestamp 1677677812
transform -1 0 1568 0 1 970
box -8 -3 104 105
use FILL  FILL_9060
timestamp 1677677812
transform 1 0 1568 0 1 970
box -8 -3 16 105
use INVX2  INVX2_575
timestamp 1677677812
transform -1 0 1592 0 1 970
box -9 -3 26 105
use FILL  FILL_9061
timestamp 1677677812
transform 1 0 1592 0 1 970
box -8 -3 16 105
use FILL  FILL_9062
timestamp 1677677812
transform 1 0 1600 0 1 970
box -8 -3 16 105
use FILL  FILL_9063
timestamp 1677677812
transform 1 0 1608 0 1 970
box -8 -3 16 105
use FILL  FILL_9078
timestamp 1677677812
transform 1 0 1616 0 1 970
box -8 -3 16 105
use FILL  FILL_9080
timestamp 1677677812
transform 1 0 1624 0 1 970
box -8 -3 16 105
use FILL  FILL_9081
timestamp 1677677812
transform 1 0 1632 0 1 970
box -8 -3 16 105
use BUFX2  BUFX2_107
timestamp 1677677812
transform 1 0 1640 0 1 970
box -5 -3 28 105
use FILL  FILL_9082
timestamp 1677677812
transform 1 0 1664 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_339
timestamp 1677677812
transform 1 0 1672 0 1 970
box -8 -3 46 105
use FILL  FILL_9083
timestamp 1677677812
transform 1 0 1712 0 1 970
box -8 -3 16 105
use FILL  FILL_9084
timestamp 1677677812
transform 1 0 1720 0 1 970
box -8 -3 16 105
use FILL  FILL_9085
timestamp 1677677812
transform 1 0 1728 0 1 970
box -8 -3 16 105
use FILL  FILL_9086
timestamp 1677677812
transform 1 0 1736 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_340
timestamp 1677677812
transform -1 0 1784 0 1 970
box -8 -3 46 105
use FILL  FILL_9087
timestamp 1677677812
transform 1 0 1784 0 1 970
box -8 -3 16 105
use FILL  FILL_9099
timestamp 1677677812
transform 1 0 1792 0 1 970
box -8 -3 16 105
use INVX2  INVX2_577
timestamp 1677677812
transform 1 0 1800 0 1 970
box -9 -3 26 105
use FILL  FILL_9100
timestamp 1677677812
transform 1 0 1816 0 1 970
box -8 -3 16 105
use FILL  FILL_9101
timestamp 1677677812
transform 1 0 1824 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_492
timestamp 1677677812
transform -1 0 1928 0 1 970
box -8 -3 104 105
use FILL  FILL_9102
timestamp 1677677812
transform 1 0 1928 0 1 970
box -8 -3 16 105
use FILL  FILL_9103
timestamp 1677677812
transform 1 0 1936 0 1 970
box -8 -3 16 105
use FILL  FILL_9104
timestamp 1677677812
transform 1 0 1944 0 1 970
box -8 -3 16 105
use FILL  FILL_9105
timestamp 1677677812
transform 1 0 1952 0 1 970
box -8 -3 16 105
use FILL  FILL_9106
timestamp 1677677812
transform 1 0 1960 0 1 970
box -8 -3 16 105
use FILL  FILL_9107
timestamp 1677677812
transform 1 0 1968 0 1 970
box -8 -3 16 105
use FILL  FILL_9108
timestamp 1677677812
transform 1 0 1976 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_341
timestamp 1677677812
transform -1 0 2024 0 1 970
box -8 -3 46 105
use FILL  FILL_9109
timestamp 1677677812
transform 1 0 2024 0 1 970
box -8 -3 16 105
use FILL  FILL_9110
timestamp 1677677812
transform 1 0 2032 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_493
timestamp 1677677812
transform -1 0 2136 0 1 970
box -8 -3 104 105
use FILL  FILL_9111
timestamp 1677677812
transform 1 0 2136 0 1 970
box -8 -3 16 105
use FILL  FILL_9120
timestamp 1677677812
transform 1 0 2144 0 1 970
box -8 -3 16 105
use FILL  FILL_9121
timestamp 1677677812
transform 1 0 2152 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_69
timestamp 1677677812
transform -1 0 2192 0 1 970
box -8 -3 40 105
use FILL  FILL_9122
timestamp 1677677812
transform 1 0 2192 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7090
timestamp 1677677812
transform 1 0 2228 0 1 975
box -3 -3 3 3
use INVX2  INVX2_578
timestamp 1677677812
transform 1 0 2200 0 1 970
box -9 -3 26 105
use M3_M2  M3_M2_7091
timestamp 1677677812
transform 1 0 2252 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_497
timestamp 1677677812
transform -1 0 2312 0 1 970
box -8 -3 104 105
use FILL  FILL_9126
timestamp 1677677812
transform 1 0 2312 0 1 970
box -8 -3 16 105
use FILL  FILL_9127
timestamp 1677677812
transform 1 0 2320 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_155
timestamp 1677677812
transform -1 0 2360 0 1 970
box -8 -3 34 105
use INVX2  INVX2_579
timestamp 1677677812
transform 1 0 2360 0 1 970
box -9 -3 26 105
use FILL  FILL_9128
timestamp 1677677812
transform 1 0 2376 0 1 970
box -8 -3 16 105
use FILL  FILL_9129
timestamp 1677677812
transform 1 0 2384 0 1 970
box -8 -3 16 105
use FILL  FILL_9130
timestamp 1677677812
transform 1 0 2392 0 1 970
box -8 -3 16 105
use FILL  FILL_9131
timestamp 1677677812
transform 1 0 2400 0 1 970
box -8 -3 16 105
use FILL  FILL_9132
timestamp 1677677812
transform 1 0 2408 0 1 970
box -8 -3 16 105
use FILL  FILL_9133
timestamp 1677677812
transform 1 0 2416 0 1 970
box -8 -3 16 105
use FILL  FILL_9134
timestamp 1677677812
transform 1 0 2424 0 1 970
box -8 -3 16 105
use FILL  FILL_9135
timestamp 1677677812
transform 1 0 2432 0 1 970
box -8 -3 16 105
use FILL  FILL_9136
timestamp 1677677812
transform 1 0 2440 0 1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_13
timestamp 1677677812
transform -1 0 2480 0 1 970
box -7 -3 39 105
use FILL  FILL_9137
timestamp 1677677812
transform 1 0 2480 0 1 970
box -8 -3 16 105
use INVX2  INVX2_582
timestamp 1677677812
transform -1 0 2504 0 1 970
box -9 -3 26 105
use XOR2X1  XOR2X1_2
timestamp 1677677812
transform -1 0 2560 0 1 970
box -8 -3 64 105
use FILL  FILL_9144
timestamp 1677677812
transform 1 0 2560 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7092
timestamp 1677677812
transform 1 0 2580 0 1 975
box -3 -3 3 3
use XOR2X1  XOR2X1_3
timestamp 1677677812
transform 1 0 2568 0 1 970
box -8 -3 64 105
use M3_M2  M3_M2_7093
timestamp 1677677812
transform 1 0 2644 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_498
timestamp 1677677812
transform -1 0 2720 0 1 970
box -8 -3 104 105
use FILL  FILL_9149
timestamp 1677677812
transform 1 0 2720 0 1 970
box -8 -3 16 105
use FILL  FILL_9150
timestamp 1677677812
transform 1 0 2728 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7094
timestamp 1677677812
transform 1 0 2844 0 1 975
box -3 -3 3 3
use FAX1  FAX1_17
timestamp 1677677812
transform 1 0 2736 0 1 970
box -5 -3 126 105
use FILL  FILL_9155
timestamp 1677677812
transform 1 0 2856 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7095
timestamp 1677677812
transform 1 0 2988 0 1 975
box -3 -3 3 3
use FAX1  FAX1_18
timestamp 1677677812
transform -1 0 2984 0 1 970
box -5 -3 126 105
use FILL  FILL_9156
timestamp 1677677812
transform 1 0 2984 0 1 970
box -8 -3 16 105
use FILL  FILL_9174
timestamp 1677677812
transform 1 0 2992 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_24
timestamp 1677677812
transform 1 0 3000 0 1 970
box -8 -3 32 105
use NAND2X1  NAND2X1_25
timestamp 1677677812
transform 1 0 3024 0 1 970
box -8 -3 32 105
use FILL  FILL_9175
timestamp 1677677812
transform 1 0 3048 0 1 970
box -8 -3 16 105
use FILL  FILL_9181
timestamp 1677677812
transform 1 0 3056 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_157
timestamp 1677677812
transform -1 0 3096 0 1 970
box -8 -3 34 105
use AOI21X1  AOI21X1_14
timestamp 1677677812
transform -1 0 3128 0 1 970
box -7 -3 39 105
use FILL  FILL_9182
timestamp 1677677812
transform 1 0 3128 0 1 970
box -8 -3 16 105
use FILL  FILL_9183
timestamp 1677677812
transform 1 0 3136 0 1 970
box -8 -3 16 105
use FILL  FILL_9184
timestamp 1677677812
transform 1 0 3144 0 1 970
box -8 -3 16 105
use FILL  FILL_9185
timestamp 1677677812
transform 1 0 3152 0 1 970
box -8 -3 16 105
use FILL  FILL_9186
timestamp 1677677812
transform 1 0 3160 0 1 970
box -8 -3 16 105
use INVX2  INVX2_584
timestamp 1677677812
transform -1 0 3184 0 1 970
box -9 -3 26 105
use FILL  FILL_9187
timestamp 1677677812
transform 1 0 3184 0 1 970
box -8 -3 16 105
use FILL  FILL_9188
timestamp 1677677812
transform 1 0 3192 0 1 970
box -8 -3 16 105
use FILL  FILL_9195
timestamp 1677677812
transform 1 0 3200 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7096
timestamp 1677677812
transform 1 0 3244 0 1 975
box -3 -3 3 3
use AOI22X1  AOI22X1_343
timestamp 1677677812
transform -1 0 3248 0 1 970
box -8 -3 46 105
use FILL  FILL_9196
timestamp 1677677812
transform 1 0 3248 0 1 970
box -8 -3 16 105
use FILL  FILL_9197
timestamp 1677677812
transform 1 0 3256 0 1 970
box -8 -3 16 105
use FILL  FILL_9198
timestamp 1677677812
transform 1 0 3264 0 1 970
box -8 -3 16 105
use FILL  FILL_9203
timestamp 1677677812
transform 1 0 3272 0 1 970
box -8 -3 16 105
use FILL  FILL_9205
timestamp 1677677812
transform 1 0 3280 0 1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_345
timestamp 1677677812
transform 1 0 3288 0 1 970
box -8 -3 46 105
use FILL  FILL_9207
timestamp 1677677812
transform 1 0 3328 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7097
timestamp 1677677812
transform 1 0 3348 0 1 975
box -3 -3 3 3
use FILL  FILL_9208
timestamp 1677677812
transform 1 0 3336 0 1 970
box -8 -3 16 105
use FILL  FILL_9209
timestamp 1677677812
transform 1 0 3344 0 1 970
box -8 -3 16 105
use FAX1  FAX1_20
timestamp 1677677812
transform 1 0 3352 0 1 970
box -5 -3 126 105
use FILL  FILL_9210
timestamp 1677677812
transform 1 0 3472 0 1 970
box -8 -3 16 105
use FILL  FILL_9211
timestamp 1677677812
transform 1 0 3480 0 1 970
box -8 -3 16 105
use INVX2  INVX2_585
timestamp 1677677812
transform 1 0 3488 0 1 970
box -9 -3 26 105
use INVX2  INVX2_586
timestamp 1677677812
transform 1 0 3504 0 1 970
box -9 -3 26 105
use FILL  FILL_9212
timestamp 1677677812
transform 1 0 3520 0 1 970
box -8 -3 16 105
use FILL  FILL_9223
timestamp 1677677812
transform 1 0 3528 0 1 970
box -8 -3 16 105
use FILL  FILL_9224
timestamp 1677677812
transform 1 0 3536 0 1 970
box -8 -3 16 105
use FILL  FILL_9225
timestamp 1677677812
transform 1 0 3544 0 1 970
box -8 -3 16 105
use AND2X2  AND2X2_54
timestamp 1677677812
transform 1 0 3552 0 1 970
box -8 -3 40 105
use FILL  FILL_9226
timestamp 1677677812
transform 1 0 3584 0 1 970
box -8 -3 16 105
use FILL  FILL_9227
timestamp 1677677812
transform 1 0 3592 0 1 970
box -8 -3 16 105
use FILL  FILL_9228
timestamp 1677677812
transform 1 0 3600 0 1 970
box -8 -3 16 105
use FILL  FILL_9229
timestamp 1677677812
transform 1 0 3608 0 1 970
box -8 -3 16 105
use FILL  FILL_9230
timestamp 1677677812
transform 1 0 3616 0 1 970
box -8 -3 16 105
use FILL  FILL_9231
timestamp 1677677812
transform 1 0 3624 0 1 970
box -8 -3 16 105
use FILL  FILL_9232
timestamp 1677677812
transform 1 0 3632 0 1 970
box -8 -3 16 105
use FILL  FILL_9233
timestamp 1677677812
transform 1 0 3640 0 1 970
box -8 -3 16 105
use FILL  FILL_9234
timestamp 1677677812
transform 1 0 3648 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_342
timestamp 1677677812
transform 1 0 3656 0 1 970
box -8 -3 46 105
use FILL  FILL_9235
timestamp 1677677812
transform 1 0 3696 0 1 970
box -8 -3 16 105
use FILL  FILL_9236
timestamp 1677677812
transform 1 0 3704 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7098
timestamp 1677677812
transform 1 0 3724 0 1 975
box -3 -3 3 3
use FILL  FILL_9237
timestamp 1677677812
transform 1 0 3712 0 1 970
box -8 -3 16 105
use FILL  FILL_9238
timestamp 1677677812
transform 1 0 3720 0 1 970
box -8 -3 16 105
use FILL  FILL_9247
timestamp 1677677812
transform 1 0 3728 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7099
timestamp 1677677812
transform 1 0 3772 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_343
timestamp 1677677812
transform 1 0 3736 0 1 970
box -8 -3 46 105
use FILL  FILL_9248
timestamp 1677677812
transform 1 0 3776 0 1 970
box -8 -3 16 105
use FILL  FILL_9249
timestamp 1677677812
transform 1 0 3784 0 1 970
box -8 -3 16 105
use FILL  FILL_9250
timestamp 1677677812
transform 1 0 3792 0 1 970
box -8 -3 16 105
use FILL  FILL_9251
timestamp 1677677812
transform 1 0 3800 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7100
timestamp 1677677812
transform 1 0 3852 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_500
timestamp 1677677812
transform -1 0 3904 0 1 970
box -8 -3 104 105
use FILL  FILL_9252
timestamp 1677677812
transform 1 0 3904 0 1 970
box -8 -3 16 105
use FILL  FILL_9253
timestamp 1677677812
transform 1 0 3912 0 1 970
box -8 -3 16 105
use FILL  FILL_9254
timestamp 1677677812
transform 1 0 3920 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_344
timestamp 1677677812
transform 1 0 3928 0 1 970
box -8 -3 46 105
use FILL  FILL_9255
timestamp 1677677812
transform 1 0 3968 0 1 970
box -8 -3 16 105
use FILL  FILL_9256
timestamp 1677677812
transform 1 0 3976 0 1 970
box -8 -3 16 105
use FILL  FILL_9257
timestamp 1677677812
transform 1 0 3984 0 1 970
box -8 -3 16 105
use FILL  FILL_9258
timestamp 1677677812
transform 1 0 3992 0 1 970
box -8 -3 16 105
use FILL  FILL_9259
timestamp 1677677812
transform 1 0 4000 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_345
timestamp 1677677812
transform -1 0 4048 0 1 970
box -8 -3 46 105
use FILL  FILL_9260
timestamp 1677677812
transform 1 0 4048 0 1 970
box -8 -3 16 105
use FILL  FILL_9261
timestamp 1677677812
transform 1 0 4056 0 1 970
box -8 -3 16 105
use FILL  FILL_9262
timestamp 1677677812
transform 1 0 4064 0 1 970
box -8 -3 16 105
use FILL  FILL_9263
timestamp 1677677812
transform 1 0 4072 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_346
timestamp 1677677812
transform -1 0 4120 0 1 970
box -8 -3 46 105
use FILL  FILL_9264
timestamp 1677677812
transform 1 0 4120 0 1 970
box -8 -3 16 105
use FILL  FILL_9287
timestamp 1677677812
transform 1 0 4128 0 1 970
box -8 -3 16 105
use FILL  FILL_9289
timestamp 1677677812
transform 1 0 4136 0 1 970
box -8 -3 16 105
use FILL  FILL_9291
timestamp 1677677812
transform 1 0 4144 0 1 970
box -8 -3 16 105
use FILL  FILL_9293
timestamp 1677677812
transform 1 0 4152 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_347
timestamp 1677677812
transform -1 0 4200 0 1 970
box -8 -3 46 105
use FILL  FILL_9294
timestamp 1677677812
transform 1 0 4200 0 1 970
box -8 -3 16 105
use FILL  FILL_9298
timestamp 1677677812
transform 1 0 4208 0 1 970
box -8 -3 16 105
use FILL  FILL_9300
timestamp 1677677812
transform 1 0 4216 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_348
timestamp 1677677812
transform 1 0 4224 0 1 970
box -8 -3 46 105
use FILL  FILL_9301
timestamp 1677677812
transform 1 0 4264 0 1 970
box -8 -3 16 105
use FILL  FILL_9305
timestamp 1677677812
transform 1 0 4272 0 1 970
box -8 -3 16 105
use FILL  FILL_9306
timestamp 1677677812
transform 1 0 4280 0 1 970
box -8 -3 16 105
use FILL  FILL_9307
timestamp 1677677812
transform 1 0 4288 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_349
timestamp 1677677812
transform -1 0 4336 0 1 970
box -8 -3 46 105
use FILL  FILL_9308
timestamp 1677677812
transform 1 0 4336 0 1 970
box -8 -3 16 105
use FILL  FILL_9309
timestamp 1677677812
transform 1 0 4344 0 1 970
box -8 -3 16 105
use FILL  FILL_9310
timestamp 1677677812
transform 1 0 4352 0 1 970
box -8 -3 16 105
use FILL  FILL_9311
timestamp 1677677812
transform 1 0 4360 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_350
timestamp 1677677812
transform 1 0 4368 0 1 970
box -8 -3 46 105
use FILL  FILL_9312
timestamp 1677677812
transform 1 0 4408 0 1 970
box -8 -3 16 105
use FILL  FILL_9313
timestamp 1677677812
transform 1 0 4416 0 1 970
box -8 -3 16 105
use FILL  FILL_9314
timestamp 1677677812
transform 1 0 4424 0 1 970
box -8 -3 16 105
use FILL  FILL_9315
timestamp 1677677812
transform 1 0 4432 0 1 970
box -8 -3 16 105
use FILL  FILL_9316
timestamp 1677677812
transform 1 0 4440 0 1 970
box -8 -3 16 105
use INVX2  INVX2_588
timestamp 1677677812
transform -1 0 4464 0 1 970
box -9 -3 26 105
use FILL  FILL_9317
timestamp 1677677812
transform 1 0 4464 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7101
timestamp 1677677812
transform 1 0 4484 0 1 975
box -3 -3 3 3
use FILL  FILL_9318
timestamp 1677677812
transform 1 0 4472 0 1 970
box -8 -3 16 105
use FILL  FILL_9319
timestamp 1677677812
transform 1 0 4480 0 1 970
box -8 -3 16 105
use FILL  FILL_9320
timestamp 1677677812
transform 1 0 4488 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_167
timestamp 1677677812
transform -1 0 4528 0 1 970
box -8 -3 34 105
use FILL  FILL_9321
timestamp 1677677812
transform 1 0 4528 0 1 970
box -8 -3 16 105
use FILL  FILL_9334
timestamp 1677677812
transform 1 0 4536 0 1 970
box -8 -3 16 105
use FILL  FILL_9336
timestamp 1677677812
transform 1 0 4544 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_352
timestamp 1677677812
transform -1 0 4592 0 1 970
box -8 -3 46 105
use FILL  FILL_9337
timestamp 1677677812
transform 1 0 4592 0 1 970
box -8 -3 16 105
use FILL  FILL_9340
timestamp 1677677812
transform 1 0 4600 0 1 970
box -8 -3 16 105
use FILL  FILL_9342
timestamp 1677677812
transform 1 0 4608 0 1 970
box -8 -3 16 105
use FILL  FILL_9344
timestamp 1677677812
transform 1 0 4616 0 1 970
box -8 -3 16 105
use FILL  FILL_9346
timestamp 1677677812
transform 1 0 4624 0 1 970
box -8 -3 16 105
use FILL  FILL_9347
timestamp 1677677812
transform 1 0 4632 0 1 970
box -8 -3 16 105
use FILL  FILL_9348
timestamp 1677677812
transform 1 0 4640 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_354
timestamp 1677677812
transform -1 0 4688 0 1 970
box -8 -3 46 105
use FILL  FILL_9349
timestamp 1677677812
transform 1 0 4688 0 1 970
box -8 -3 16 105
use FILL  FILL_9350
timestamp 1677677812
transform 1 0 4696 0 1 970
box -8 -3 16 105
use FILL  FILL_9351
timestamp 1677677812
transform 1 0 4704 0 1 970
box -8 -3 16 105
use FILL  FILL_9352
timestamp 1677677812
transform 1 0 4712 0 1 970
box -8 -3 16 105
use FILL  FILL_9353
timestamp 1677677812
transform 1 0 4720 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_7102
timestamp 1677677812
transform 1 0 4740 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_7103
timestamp 1677677812
transform 1 0 4756 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_355
timestamp 1677677812
transform -1 0 4768 0 1 970
box -8 -3 46 105
use FILL  FILL_9354
timestamp 1677677812
transform 1 0 4768 0 1 970
box -8 -3 16 105
use FILL  FILL_9355
timestamp 1677677812
transform 1 0 4776 0 1 970
box -8 -3 16 105
use FILL  FILL_9356
timestamp 1677677812
transform 1 0 4784 0 1 970
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_75
timestamp 1677677812
transform 1 0 4819 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_7104
timestamp 1677677812
transform 1 0 188 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7943
timestamp 1677677812
transform 1 0 92 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7166
timestamp 1677677812
transform 1 0 172 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7178
timestamp 1677677812
transform 1 0 92 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7944
timestamp 1677677812
transform 1 0 196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8045
timestamp 1677677812
transform 1 0 140 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8046
timestamp 1677677812
transform 1 0 172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8047
timestamp 1677677812
transform 1 0 180 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8048
timestamp 1677677812
transform 1 0 188 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7204
timestamp 1677677812
transform 1 0 140 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7205
timestamp 1677677812
transform 1 0 180 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7206
timestamp 1677677812
transform 1 0 196 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7241
timestamp 1677677812
transform 1 0 188 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7105
timestamp 1677677812
transform 1 0 236 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7945
timestamp 1677677812
transform 1 0 212 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7167
timestamp 1677677812
transform 1 0 220 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7946
timestamp 1677677812
transform 1 0 228 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7947
timestamp 1677677812
transform 1 0 236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8049
timestamp 1677677812
transform 1 0 220 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7207
timestamp 1677677812
transform 1 0 220 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8050
timestamp 1677677812
transform 1 0 244 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7948
timestamp 1677677812
transform 1 0 252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7949
timestamp 1677677812
transform 1 0 292 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7179
timestamp 1677677812
transform 1 0 292 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8051
timestamp 1677677812
transform 1 0 340 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8052
timestamp 1677677812
transform 1 0 372 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8053
timestamp 1677677812
transform 1 0 380 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7208
timestamp 1677677812
transform 1 0 340 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7209
timestamp 1677677812
transform 1 0 380 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7950
timestamp 1677677812
transform 1 0 404 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7951
timestamp 1677677812
transform 1 0 412 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8054
timestamp 1677677812
transform 1 0 420 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7952
timestamp 1677677812
transform 1 0 444 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8055
timestamp 1677677812
transform 1 0 468 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8056
timestamp 1677677812
transform 1 0 556 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7210
timestamp 1677677812
transform 1 0 556 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7953
timestamp 1677677812
transform 1 0 580 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7954
timestamp 1677677812
transform 1 0 596 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8057
timestamp 1677677812
transform 1 0 572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8058
timestamp 1677677812
transform 1 0 588 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7211
timestamp 1677677812
transform 1 0 596 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7242
timestamp 1677677812
transform 1 0 572 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8059
timestamp 1677677812
transform 1 0 620 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8060
timestamp 1677677812
transform 1 0 636 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7126
timestamp 1677677812
transform 1 0 660 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7955
timestamp 1677677812
transform 1 0 660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8061
timestamp 1677677812
transform 1 0 652 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8062
timestamp 1677677812
transform 1 0 668 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7243
timestamp 1677677812
transform 1 0 668 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7141
timestamp 1677677812
transform 1 0 716 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7956
timestamp 1677677812
transform 1 0 716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7957
timestamp 1677677812
transform 1 0 732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8063
timestamp 1677677812
transform 1 0 780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8064
timestamp 1677677812
transform 1 0 812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8065
timestamp 1677677812
transform 1 0 820 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7212
timestamp 1677677812
transform 1 0 780 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7244
timestamp 1677677812
transform 1 0 804 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7288
timestamp 1677677812
transform 1 0 740 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7213
timestamp 1677677812
transform 1 0 820 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7245
timestamp 1677677812
transform 1 0 828 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7142
timestamp 1677677812
transform 1 0 860 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7958
timestamp 1677677812
transform 1 0 852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7959
timestamp 1677677812
transform 1 0 860 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7143
timestamp 1677677812
transform 1 0 876 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8066
timestamp 1677677812
transform 1 0 868 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7246
timestamp 1677677812
transform 1 0 868 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7106
timestamp 1677677812
transform 1 0 924 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7144
timestamp 1677677812
transform 1 0 932 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7960
timestamp 1677677812
transform 1 0 908 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7961
timestamp 1677677812
transform 1 0 932 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8067
timestamp 1677677812
transform 1 0 916 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8068
timestamp 1677677812
transform 1 0 932 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7214
timestamp 1677677812
transform 1 0 916 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7272
timestamp 1677677812
transform 1 0 932 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7107
timestamp 1677677812
transform 1 0 964 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8069
timestamp 1677677812
transform 1 0 972 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7962
timestamp 1677677812
transform 1 0 980 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7215
timestamp 1677677812
transform 1 0 980 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7127
timestamp 1677677812
transform 1 0 1012 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7937
timestamp 1677677812
transform 1 0 1012 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_7963
timestamp 1677677812
transform 1 0 1036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7964
timestamp 1677677812
transform 1 0 1100 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8070
timestamp 1677677812
transform 1 0 1108 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8071
timestamp 1677677812
transform 1 0 1116 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8072
timestamp 1677677812
transform 1 0 1132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8073
timestamp 1677677812
transform 1 0 1148 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7216
timestamp 1677677812
transform 1 0 1108 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7247
timestamp 1677677812
transform 1 0 1100 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7273
timestamp 1677677812
transform 1 0 1116 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7274
timestamp 1677677812
transform 1 0 1148 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7965
timestamp 1677677812
transform 1 0 1164 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7180
timestamp 1677677812
transform 1 0 1164 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8150
timestamp 1677677812
transform 1 0 1164 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7289
timestamp 1677677812
transform 1 0 1164 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7966
timestamp 1677677812
transform 1 0 1188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7967
timestamp 1677677812
transform 1 0 1196 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7181
timestamp 1677677812
transform 1 0 1196 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7248
timestamp 1677677812
transform 1 0 1188 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7108
timestamp 1677677812
transform 1 0 1220 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8074
timestamp 1677677812
transform 1 0 1212 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7249
timestamp 1677677812
transform 1 0 1212 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7968
timestamp 1677677812
transform 1 0 1236 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8075
timestamp 1677677812
transform 1 0 1228 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7217
timestamp 1677677812
transform 1 0 1236 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7275
timestamp 1677677812
transform 1 0 1244 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8076
timestamp 1677677812
transform 1 0 1260 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7128
timestamp 1677677812
transform 1 0 1284 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7969
timestamp 1677677812
transform 1 0 1284 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7145
timestamp 1677677812
transform 1 0 1300 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7146
timestamp 1677677812
transform 1 0 1364 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7970
timestamp 1677677812
transform 1 0 1300 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7168
timestamp 1677677812
transform 1 0 1388 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7147
timestamp 1677677812
transform 1 0 1420 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7971
timestamp 1677677812
transform 1 0 1396 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8077
timestamp 1677677812
transform 1 0 1324 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7182
timestamp 1677677812
transform 1 0 1348 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8078
timestamp 1677677812
transform 1 0 1380 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8079
timestamp 1677677812
transform 1 0 1388 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8080
timestamp 1677677812
transform 1 0 1404 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8081
timestamp 1677677812
transform 1 0 1420 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7250
timestamp 1677677812
transform 1 0 1340 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7251
timestamp 1677677812
transform 1 0 1372 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7276
timestamp 1677677812
transform 1 0 1332 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7218
timestamp 1677677812
transform 1 0 1404 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7252
timestamp 1677677812
transform 1 0 1420 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7129
timestamp 1677677812
transform 1 0 1436 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7148
timestamp 1677677812
transform 1 0 1452 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7972
timestamp 1677677812
transform 1 0 1436 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7169
timestamp 1677677812
transform 1 0 1444 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7973
timestamp 1677677812
transform 1 0 1452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8082
timestamp 1677677812
transform 1 0 1444 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7219
timestamp 1677677812
transform 1 0 1436 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8178
timestamp 1677677812
transform 1 0 1428 0 1 885
box -2 -2 2 2
use M3_M2  M3_M2_7253
timestamp 1677677812
transform 1 0 1452 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7974
timestamp 1677677812
transform 1 0 1532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8083
timestamp 1677677812
transform 1 0 1524 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7183
timestamp 1677677812
transform 1 0 1532 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8084
timestamp 1677677812
transform 1 0 1604 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7109
timestamp 1677677812
transform 1 0 1652 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7130
timestamp 1677677812
transform 1 0 1644 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7975
timestamp 1677677812
transform 1 0 1636 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7976
timestamp 1677677812
transform 1 0 1652 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8085
timestamp 1677677812
transform 1 0 1628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8086
timestamp 1677677812
transform 1 0 1644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8087
timestamp 1677677812
transform 1 0 1660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8088
timestamp 1677677812
transform 1 0 1668 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7220
timestamp 1677677812
transform 1 0 1668 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7131
timestamp 1677677812
transform 1 0 1684 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7132
timestamp 1677677812
transform 1 0 1700 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7977
timestamp 1677677812
transform 1 0 1700 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7978
timestamp 1677677812
transform 1 0 1708 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7979
timestamp 1677677812
transform 1 0 1724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7980
timestamp 1677677812
transform 1 0 1740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8089
timestamp 1677677812
transform 1 0 1732 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7221
timestamp 1677677812
transform 1 0 1708 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7254
timestamp 1677677812
transform 1 0 1732 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8090
timestamp 1677677812
transform 1 0 1748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7981
timestamp 1677677812
transform 1 0 1884 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8091
timestamp 1677677812
transform 1 0 1836 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8092
timestamp 1677677812
transform 1 0 1900 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7222
timestamp 1677677812
transform 1 0 1900 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7110
timestamp 1677677812
transform 1 0 1964 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7111
timestamp 1677677812
transform 1 0 2012 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7112
timestamp 1677677812
transform 1 0 2052 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7113
timestamp 1677677812
transform 1 0 2084 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7982
timestamp 1677677812
transform 1 0 1996 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7133
timestamp 1677677812
transform 1 0 2100 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_7983
timestamp 1677677812
transform 1 0 2092 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8093
timestamp 1677677812
transform 1 0 1964 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8094
timestamp 1677677812
transform 1 0 2012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8095
timestamp 1677677812
transform 1 0 2068 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7290
timestamp 1677677812
transform 1 0 2028 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8151
timestamp 1677677812
transform 1 0 2108 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7255
timestamp 1677677812
transform 1 0 2108 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7134
timestamp 1677677812
transform 1 0 2132 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8152
timestamp 1677677812
transform 1 0 2156 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7223
timestamp 1677677812
transform 1 0 2164 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8153
timestamp 1677677812
transform 1 0 2180 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8173
timestamp 1677677812
transform 1 0 2164 0 1 905
box -2 -2 2 2
use M2_M1  M2_M1_8154
timestamp 1677677812
transform 1 0 2196 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8174
timestamp 1677677812
transform 1 0 2188 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_7277
timestamp 1677677812
transform 1 0 2188 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7291
timestamp 1677677812
transform 1 0 2180 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7114
timestamp 1677677812
transform 1 0 2228 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7224
timestamp 1677677812
transform 1 0 2220 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8175
timestamp 1677677812
transform 1 0 2220 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_7225
timestamp 1677677812
transform 1 0 2236 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8176
timestamp 1677677812
transform 1 0 2236 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_7115
timestamp 1677677812
transform 1 0 2300 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7984
timestamp 1677677812
transform 1 0 2284 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7985
timestamp 1677677812
transform 1 0 2292 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7986
timestamp 1677677812
transform 1 0 2308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8096
timestamp 1677677812
transform 1 0 2260 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8097
timestamp 1677677812
transform 1 0 2268 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7184
timestamp 1677677812
transform 1 0 2276 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7185
timestamp 1677677812
transform 1 0 2308 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8098
timestamp 1677677812
transform 1 0 2332 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7226
timestamp 1677677812
transform 1 0 2292 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8155
timestamp 1677677812
transform 1 0 2308 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7292
timestamp 1677677812
transform 1 0 2284 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7256
timestamp 1677677812
transform 1 0 2308 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7257
timestamp 1677677812
transform 1 0 2324 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7293
timestamp 1677677812
transform 1 0 2316 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7938
timestamp 1677677812
transform 1 0 2364 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_7987
timestamp 1677677812
transform 1 0 2348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7988
timestamp 1677677812
transform 1 0 2356 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7989
timestamp 1677677812
transform 1 0 2468 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8099
timestamp 1677677812
transform 1 0 2452 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7227
timestamp 1677677812
transform 1 0 2468 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8100
timestamp 1677677812
transform 1 0 2484 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8101
timestamp 1677677812
transform 1 0 2492 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7258
timestamp 1677677812
transform 1 0 2484 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7990
timestamp 1677677812
transform 1 0 2508 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7228
timestamp 1677677812
transform 1 0 2508 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7991
timestamp 1677677812
transform 1 0 2524 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7294
timestamp 1677677812
transform 1 0 2524 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8102
timestamp 1677677812
transform 1 0 2540 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7186
timestamp 1677677812
transform 1 0 2548 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8103
timestamp 1677677812
transform 1 0 2556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8104
timestamp 1677677812
transform 1 0 2564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_7992
timestamp 1677677812
transform 1 0 2580 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7278
timestamp 1677677812
transform 1 0 2588 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_7993
timestamp 1677677812
transform 1 0 2620 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7116
timestamp 1677677812
transform 1 0 2652 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7117
timestamp 1677677812
transform 1 0 2676 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_7994
timestamp 1677677812
transform 1 0 2716 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8105
timestamp 1677677812
transform 1 0 2612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8106
timestamp 1677677812
transform 1 0 2628 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8107
timestamp 1677677812
transform 1 0 2636 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8108
timestamp 1677677812
transform 1 0 2692 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7229
timestamp 1677677812
transform 1 0 2612 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7259
timestamp 1677677812
transform 1 0 2636 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_7995
timestamp 1677677812
transform 1 0 2732 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7187
timestamp 1677677812
transform 1 0 2732 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_7939
timestamp 1677677812
transform 1 0 2852 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7170
timestamp 1677677812
transform 1 0 2756 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7171
timestamp 1677677812
transform 1 0 2852 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_7996
timestamp 1677677812
transform 1 0 2860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_7997
timestamp 1677677812
transform 1 0 2868 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8109
timestamp 1677677812
transform 1 0 2748 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8110
timestamp 1677677812
transform 1 0 2764 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7295
timestamp 1677677812
transform 1 0 2852 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7118
timestamp 1677677812
transform 1 0 2980 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8156
timestamp 1677677812
transform 1 0 3012 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_7940
timestamp 1677677812
transform 1 0 3028 0 1 945
box -2 -2 2 2
use M2_M1  M2_M1_7998
timestamp 1677677812
transform 1 0 3068 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7230
timestamp 1677677812
transform 1 0 3068 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_7941
timestamp 1677677812
transform 1 0 3076 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7172
timestamp 1677677812
transform 1 0 3084 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8111
timestamp 1677677812
transform 1 0 3076 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8112
timestamp 1677677812
transform 1 0 3084 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7260
timestamp 1677677812
transform 1 0 3076 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8113
timestamp 1677677812
transform 1 0 3108 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7173
timestamp 1677677812
transform 1 0 3124 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8157
timestamp 1677677812
transform 1 0 3116 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7261
timestamp 1677677812
transform 1 0 3116 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7135
timestamp 1677677812
transform 1 0 3164 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7149
timestamp 1677677812
transform 1 0 3156 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_7999
timestamp 1677677812
transform 1 0 3156 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7174
timestamp 1677677812
transform 1 0 3164 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8114
timestamp 1677677812
transform 1 0 3148 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7188
timestamp 1677677812
transform 1 0 3156 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7119
timestamp 1677677812
transform 1 0 3188 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8115
timestamp 1677677812
transform 1 0 3180 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7231
timestamp 1677677812
transform 1 0 3148 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8158
timestamp 1677677812
transform 1 0 3164 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8177
timestamp 1677677812
transform 1 0 3172 0 1 905
box -2 -2 2 2
use M3_M2  M3_M2_7150
timestamp 1677677812
transform 1 0 3220 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8000
timestamp 1677677812
transform 1 0 3220 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8116
timestamp 1677677812
transform 1 0 3212 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7189
timestamp 1677677812
transform 1 0 3220 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8159
timestamp 1677677812
transform 1 0 3220 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7136
timestamp 1677677812
transform 1 0 3236 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7151
timestamp 1677677812
transform 1 0 3260 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8001
timestamp 1677677812
transform 1 0 3252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8002
timestamp 1677677812
transform 1 0 3260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8117
timestamp 1677677812
transform 1 0 3244 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7232
timestamp 1677677812
transform 1 0 3268 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8118
timestamp 1677677812
transform 1 0 3292 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7262
timestamp 1677677812
transform 1 0 3292 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7190
timestamp 1677677812
transform 1 0 3308 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7120
timestamp 1677677812
transform 1 0 3324 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7152
timestamp 1677677812
transform 1 0 3324 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7175
timestamp 1677677812
transform 1 0 3340 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8003
timestamp 1677677812
transform 1 0 3348 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8119
timestamp 1677677812
transform 1 0 3324 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7191
timestamp 1677677812
transform 1 0 3332 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8120
timestamp 1677677812
transform 1 0 3340 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7296
timestamp 1677677812
transform 1 0 3324 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8004
timestamp 1677677812
transform 1 0 3372 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8121
timestamp 1677677812
transform 1 0 3372 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7279
timestamp 1677677812
transform 1 0 3372 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7297
timestamp 1677677812
transform 1 0 3364 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_7942
timestamp 1677677812
transform 1 0 3388 0 1 945
box -2 -2 2 2
use M3_M2  M3_M2_7153
timestamp 1677677812
transform 1 0 3508 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8005
timestamp 1677677812
transform 1 0 3492 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8006
timestamp 1677677812
transform 1 0 3500 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7192
timestamp 1677677812
transform 1 0 3388 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8122
timestamp 1677677812
transform 1 0 3476 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8123
timestamp 1677677812
transform 1 0 3484 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7280
timestamp 1677677812
transform 1 0 3484 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7233
timestamp 1677677812
transform 1 0 3500 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7298
timestamp 1677677812
transform 1 0 3396 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7299
timestamp 1677677812
transform 1 0 3492 0 1 885
box -3 -3 3 3
use M2_M1  M2_M1_8007
timestamp 1677677812
transform 1 0 3532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8124
timestamp 1677677812
transform 1 0 3540 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8125
timestamp 1677677812
transform 1 0 3572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8008
timestamp 1677677812
transform 1 0 3580 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7176
timestamp 1677677812
transform 1 0 3596 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_8009
timestamp 1677677812
transform 1 0 3604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8126
timestamp 1677677812
transform 1 0 3596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8127
timestamp 1677677812
transform 1 0 3612 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8128
timestamp 1677677812
transform 1 0 3644 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8160
timestamp 1677677812
transform 1 0 3628 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8010
timestamp 1677677812
transform 1 0 3660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8011
timestamp 1677677812
transform 1 0 3668 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7234
timestamp 1677677812
transform 1 0 3660 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7177
timestamp 1677677812
transform 1 0 3684 0 1 935
box -3 -3 3 3
use M3_M2  M3_M2_7121
timestamp 1677677812
transform 1 0 3708 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7154
timestamp 1677677812
transform 1 0 3700 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8129
timestamp 1677677812
transform 1 0 3700 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7193
timestamp 1677677812
transform 1 0 3716 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8161
timestamp 1677677812
transform 1 0 3716 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8012
timestamp 1677677812
transform 1 0 3724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8013
timestamp 1677677812
transform 1 0 3732 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7155
timestamp 1677677812
transform 1 0 3756 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8130
timestamp 1677677812
transform 1 0 3740 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7194
timestamp 1677677812
transform 1 0 3756 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8162
timestamp 1677677812
transform 1 0 3756 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8131
timestamp 1677677812
transform 1 0 3780 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8132
timestamp 1677677812
transform 1 0 3804 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7263
timestamp 1677677812
transform 1 0 3804 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7122
timestamp 1677677812
transform 1 0 3860 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8014
timestamp 1677677812
transform 1 0 3852 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8015
timestamp 1677677812
transform 1 0 3860 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8163
timestamp 1677677812
transform 1 0 3900 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8016
timestamp 1677677812
transform 1 0 3924 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8017
timestamp 1677677812
transform 1 0 3948 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7156
timestamp 1677677812
transform 1 0 3980 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8018
timestamp 1677677812
transform 1 0 3972 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8133
timestamp 1677677812
transform 1 0 3980 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7195
timestamp 1677677812
transform 1 0 3996 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8164
timestamp 1677677812
transform 1 0 3996 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7264
timestamp 1677677812
transform 1 0 3996 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8134
timestamp 1677677812
transform 1 0 4012 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7157
timestamp 1677677812
transform 1 0 4028 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_7137
timestamp 1677677812
transform 1 0 4044 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7158
timestamp 1677677812
transform 1 0 4060 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8019
timestamp 1677677812
transform 1 0 4044 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8020
timestamp 1677677812
transform 1 0 4052 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8135
timestamp 1677677812
transform 1 0 4060 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8165
timestamp 1677677812
transform 1 0 4076 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7159
timestamp 1677677812
transform 1 0 4100 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8136
timestamp 1677677812
transform 1 0 4092 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7281
timestamp 1677677812
transform 1 0 4092 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8137
timestamp 1677677812
transform 1 0 4132 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7265
timestamp 1677677812
transform 1 0 4124 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7300
timestamp 1677677812
transform 1 0 4124 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7160
timestamp 1677677812
transform 1 0 4148 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8021
timestamp 1677677812
transform 1 0 4148 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7196
timestamp 1677677812
transform 1 0 4156 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8138
timestamp 1677677812
transform 1 0 4164 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8166
timestamp 1677677812
transform 1 0 4180 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7266
timestamp 1677677812
transform 1 0 4164 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7267
timestamp 1677677812
transform 1 0 4180 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7161
timestamp 1677677812
transform 1 0 4196 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8022
timestamp 1677677812
transform 1 0 4188 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8023
timestamp 1677677812
transform 1 0 4196 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8167
timestamp 1677677812
transform 1 0 4196 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7282
timestamp 1677677812
transform 1 0 4196 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7268
timestamp 1677677812
transform 1 0 4212 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_8024
timestamp 1677677812
transform 1 0 4252 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8025
timestamp 1677677812
transform 1 0 4260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8139
timestamp 1677677812
transform 1 0 4244 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7197
timestamp 1677677812
transform 1 0 4260 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7198
timestamp 1677677812
transform 1 0 4276 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8168
timestamp 1677677812
transform 1 0 4284 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7269
timestamp 1677677812
transform 1 0 4284 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7123
timestamp 1677677812
transform 1 0 4324 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7162
timestamp 1677677812
transform 1 0 4332 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8026
timestamp 1677677812
transform 1 0 4308 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8027
timestamp 1677677812
transform 1 0 4316 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8028
timestamp 1677677812
transform 1 0 4324 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8169
timestamp 1677677812
transform 1 0 4316 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7283
timestamp 1677677812
transform 1 0 4316 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8029
timestamp 1677677812
transform 1 0 4364 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7199
timestamp 1677677812
transform 1 0 4364 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8170
timestamp 1677677812
transform 1 0 4372 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7270
timestamp 1677677812
transform 1 0 4372 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7124
timestamp 1677677812
transform 1 0 4396 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_7138
timestamp 1677677812
transform 1 0 4396 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8030
timestamp 1677677812
transform 1 0 4388 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8031
timestamp 1677677812
transform 1 0 4396 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7139
timestamp 1677677812
transform 1 0 4460 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_7163
timestamp 1677677812
transform 1 0 4460 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8032
timestamp 1677677812
transform 1 0 4428 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8033
timestamp 1677677812
transform 1 0 4436 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8034
timestamp 1677677812
transform 1 0 4452 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8035
timestamp 1677677812
transform 1 0 4468 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7200
timestamp 1677677812
transform 1 0 4412 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8140
timestamp 1677677812
transform 1 0 4428 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7201
timestamp 1677677812
transform 1 0 4436 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_8141
timestamp 1677677812
transform 1 0 4444 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8142
timestamp 1677677812
transform 1 0 4460 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7235
timestamp 1677677812
transform 1 0 4428 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7236
timestamp 1677677812
transform 1 0 4452 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_8036
timestamp 1677677812
transform 1 0 4484 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8171
timestamp 1677677812
transform 1 0 4484 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_7284
timestamp 1677677812
transform 1 0 4484 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7237
timestamp 1677677812
transform 1 0 4508 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7285
timestamp 1677677812
transform 1 0 4516 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_7164
timestamp 1677677812
transform 1 0 4548 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8037
timestamp 1677677812
transform 1 0 4540 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7202
timestamp 1677677812
transform 1 0 4540 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7165
timestamp 1677677812
transform 1 0 4572 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_8038
timestamp 1677677812
transform 1 0 4556 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8039
timestamp 1677677812
transform 1 0 4572 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8143
timestamp 1677677812
transform 1 0 4548 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7140
timestamp 1677677812
transform 1 0 4596 0 1 955
box -3 -3 3 3
use M2_M1  M2_M1_8144
timestamp 1677677812
transform 1 0 4564 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8145
timestamp 1677677812
transform 1 0 4580 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7203
timestamp 1677677812
transform 1 0 4588 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_7238
timestamp 1677677812
transform 1 0 4564 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7286
timestamp 1677677812
transform 1 0 4556 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8172
timestamp 1677677812
transform 1 0 4596 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_8040
timestamp 1677677812
transform 1 0 4604 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8041
timestamp 1677677812
transform 1 0 4612 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_7301
timestamp 1677677812
transform 1 0 4596 0 1 885
box -3 -3 3 3
use M3_M2  M3_M2_7271
timestamp 1677677812
transform 1 0 4612 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_7125
timestamp 1677677812
transform 1 0 4660 0 1 965
box -3 -3 3 3
use M2_M1  M2_M1_8042
timestamp 1677677812
transform 1 0 4660 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8146
timestamp 1677677812
transform 1 0 4668 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7287
timestamp 1677677812
transform 1 0 4676 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_8043
timestamp 1677677812
transform 1 0 4692 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8044
timestamp 1677677812
transform 1 0 4788 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_8147
timestamp 1677677812
transform 1 0 4740 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8148
timestamp 1677677812
transform 1 0 4772 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_8149
timestamp 1677677812
transform 1 0 4796 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_7239
timestamp 1677677812
transform 1 0 4772 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_7240
timestamp 1677677812
transform 1 0 4788 0 1 915
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_76
timestamp 1677677812
transform 1 0 24 0 1 870
box -10 -3 10 3
use FILL  FILL_8944
timestamp 1677677812
transform 1 0 72 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_483
timestamp 1677677812
transform 1 0 80 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_566
timestamp 1677677812
transform -1 0 192 0 -1 970
box -9 -3 26 105
use FILL  FILL_8945
timestamp 1677677812
transform 1 0 192 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_331
timestamp 1677677812
transform 1 0 200 0 -1 970
box -8 -3 46 105
use FILL  FILL_8946
timestamp 1677677812
transform 1 0 240 0 -1 970
box -8 -3 16 105
use FILL  FILL_8947
timestamp 1677677812
transform 1 0 248 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_567
timestamp 1677677812
transform 1 0 256 0 -1 970
box -9 -3 26 105
use FILL  FILL_8948
timestamp 1677677812
transform 1 0 272 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_484
timestamp 1677677812
transform 1 0 280 0 -1 970
box -8 -3 104 105
use FILL  FILL_8949
timestamp 1677677812
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_8950
timestamp 1677677812
transform 1 0 384 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_568
timestamp 1677677812
transform -1 0 408 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_569
timestamp 1677677812
transform 1 0 408 0 -1 970
box -9 -3 26 105
use FILL  FILL_8951
timestamp 1677677812
transform 1 0 424 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_486
timestamp 1677677812
transform 1 0 432 0 -1 970
box -8 -3 104 105
use FILL  FILL_8955
timestamp 1677677812
transform 1 0 528 0 -1 970
box -8 -3 16 105
use FILL  FILL_8956
timestamp 1677677812
transform 1 0 536 0 -1 970
box -8 -3 16 105
use FILL  FILL_8957
timestamp 1677677812
transform 1 0 544 0 -1 970
box -8 -3 16 105
use FILL  FILL_8958
timestamp 1677677812
transform 1 0 552 0 -1 970
box -8 -3 16 105
use FILL  FILL_8959
timestamp 1677677812
transform 1 0 560 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_333
timestamp 1677677812
transform 1 0 568 0 -1 970
box -8 -3 46 105
use FILL  FILL_8967
timestamp 1677677812
transform 1 0 608 0 -1 970
box -8 -3 16 105
use FILL  FILL_8968
timestamp 1677677812
transform 1 0 616 0 -1 970
box -8 -3 16 105
use FILL  FILL_8969
timestamp 1677677812
transform 1 0 624 0 -1 970
box -8 -3 16 105
use FILL  FILL_8970
timestamp 1677677812
transform 1 0 632 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_336
timestamp 1677677812
transform 1 0 640 0 -1 970
box -8 -3 46 105
use FILL  FILL_8971
timestamp 1677677812
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_8972
timestamp 1677677812
transform 1 0 688 0 -1 970
box -8 -3 16 105
use FILL  FILL_8973
timestamp 1677677812
transform 1 0 696 0 -1 970
box -8 -3 16 105
use FILL  FILL_8975
timestamp 1677677812
transform 1 0 704 0 -1 970
box -8 -3 16 105
use FILL  FILL_8977
timestamp 1677677812
transform 1 0 712 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_488
timestamp 1677677812
transform 1 0 720 0 -1 970
box -8 -3 104 105
use FILL  FILL_8980
timestamp 1677677812
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_8981
timestamp 1677677812
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_8983
timestamp 1677677812
transform 1 0 832 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_572
timestamp 1677677812
transform -1 0 856 0 -1 970
box -9 -3 26 105
use FILL  FILL_8985
timestamp 1677677812
transform 1 0 856 0 -1 970
box -8 -3 16 105
use FILL  FILL_8987
timestamp 1677677812
transform 1 0 864 0 -1 970
box -8 -3 16 105
use FILL  FILL_8992
timestamp 1677677812
transform 1 0 872 0 -1 970
box -8 -3 16 105
use FILL  FILL_8993
timestamp 1677677812
transform 1 0 880 0 -1 970
box -8 -3 16 105
use FILL  FILL_8994
timestamp 1677677812
transform 1 0 888 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_335
timestamp 1677677812
transform -1 0 936 0 -1 970
box -8 -3 46 105
use FILL  FILL_8995
timestamp 1677677812
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_8997
timestamp 1677677812
transform 1 0 944 0 -1 970
box -8 -3 16 105
use FILL  FILL_9002
timestamp 1677677812
transform 1 0 952 0 -1 970
box -8 -3 16 105
use FILL  FILL_9003
timestamp 1677677812
transform 1 0 960 0 -1 970
box -8 -3 16 105
use FILL  FILL_9004
timestamp 1677677812
transform 1 0 968 0 -1 970
box -8 -3 16 105
use FILL  FILL_9005
timestamp 1677677812
transform 1 0 976 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_573
timestamp 1677677812
transform 1 0 984 0 -1 970
box -9 -3 26 105
use FILL  FILL_9006
timestamp 1677677812
transform 1 0 1000 0 -1 970
box -8 -3 16 105
use FILL  FILL_9007
timestamp 1677677812
transform 1 0 1008 0 -1 970
box -8 -3 16 105
use FILL  FILL_9008
timestamp 1677677812
transform 1 0 1016 0 -1 970
box -8 -3 16 105
use FILL  FILL_9009
timestamp 1677677812
transform 1 0 1024 0 -1 970
box -8 -3 16 105
use FILL  FILL_9010
timestamp 1677677812
transform 1 0 1032 0 -1 970
box -8 -3 16 105
use FILL  FILL_9011
timestamp 1677677812
transform 1 0 1040 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_89
timestamp 1677677812
transform 1 0 1048 0 -1 970
box -8 -3 32 105
use FILL  FILL_9012
timestamp 1677677812
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_9014
timestamp 1677677812
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use FILL  FILL_9019
timestamp 1677677812
transform 1 0 1088 0 -1 970
box -8 -3 16 105
use FILL  FILL_9020
timestamp 1677677812
transform 1 0 1096 0 -1 970
box -8 -3 16 105
use FILL  FILL_9021
timestamp 1677677812
transform 1 0 1104 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_337
timestamp 1677677812
transform 1 0 1112 0 -1 970
box -8 -3 46 105
use FILL  FILL_9022
timestamp 1677677812
transform 1 0 1152 0 -1 970
box -8 -3 16 105
use FILL  FILL_9024
timestamp 1677677812
transform 1 0 1160 0 -1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_91
timestamp 1677677812
transform 1 0 1168 0 -1 970
box -8 -3 32 105
use FILL  FILL_9026
timestamp 1677677812
transform 1 0 1192 0 -1 970
box -8 -3 16 105
use FILL  FILL_9028
timestamp 1677677812
transform 1 0 1200 0 -1 970
box -8 -3 16 105
use FILL  FILL_9032
timestamp 1677677812
transform 1 0 1208 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_338
timestamp 1677677812
transform -1 0 1256 0 -1 970
box -8 -3 46 105
use FILL  FILL_9033
timestamp 1677677812
transform 1 0 1256 0 -1 970
box -8 -3 16 105
use FILL  FILL_9034
timestamp 1677677812
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_9036
timestamp 1677677812
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_9038
timestamp 1677677812
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7302
timestamp 1677677812
transform 1 0 1300 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_490
timestamp 1677677812
transform 1 0 1288 0 -1 970
box -8 -3 104 105
use AOI22X1  AOI22X1_339
timestamp 1677677812
transform -1 0 1424 0 -1 970
box -8 -3 46 105
use FILL  FILL_9055
timestamp 1677677812
transform 1 0 1424 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_574
timestamp 1677677812
transform 1 0 1432 0 -1 970
box -9 -3 26 105
use FILL  FILL_9056
timestamp 1677677812
transform 1 0 1448 0 -1 970
box -8 -3 16 105
use FILL  FILL_9058
timestamp 1677677812
transform 1 0 1456 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7303
timestamp 1677677812
transform 1 0 1476 0 1 875
box -3 -3 3 3
use FILL  FILL_9064
timestamp 1677677812
transform 1 0 1464 0 -1 970
box -8 -3 16 105
use FILL  FILL_9065
timestamp 1677677812
transform 1 0 1472 0 -1 970
box -8 -3 16 105
use FILL  FILL_9066
timestamp 1677677812
transform 1 0 1480 0 -1 970
box -8 -3 16 105
use FILL  FILL_9067
timestamp 1677677812
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use FILL  FILL_9068
timestamp 1677677812
transform 1 0 1496 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_576
timestamp 1677677812
transform 1 0 1504 0 -1 970
box -9 -3 26 105
use FILL  FILL_9069
timestamp 1677677812
transform 1 0 1520 0 -1 970
box -8 -3 16 105
use FILL  FILL_9070
timestamp 1677677812
transform 1 0 1528 0 -1 970
box -8 -3 16 105
use FILL  FILL_9071
timestamp 1677677812
transform 1 0 1536 0 -1 970
box -8 -3 16 105
use FILL  FILL_9072
timestamp 1677677812
transform 1 0 1544 0 -1 970
box -8 -3 16 105
use FILL  FILL_9073
timestamp 1677677812
transform 1 0 1552 0 -1 970
box -8 -3 16 105
use FILL  FILL_9074
timestamp 1677677812
transform 1 0 1560 0 -1 970
box -8 -3 16 105
use FILL  FILL_9075
timestamp 1677677812
transform 1 0 1568 0 -1 970
box -8 -3 16 105
use FILL  FILL_9076
timestamp 1677677812
transform 1 0 1576 0 -1 970
box -8 -3 16 105
use BUFX2  BUFX2_106
timestamp 1677677812
transform -1 0 1608 0 -1 970
box -5 -3 28 105
use FILL  FILL_9077
timestamp 1677677812
transform 1 0 1608 0 -1 970
box -8 -3 16 105
use FILL  FILL_9079
timestamp 1677677812
transform 1 0 1616 0 -1 970
box -8 -3 16 105
use FILL  FILL_9088
timestamp 1677677812
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_340
timestamp 1677677812
transform -1 0 1672 0 -1 970
box -8 -3 46 105
use FILL  FILL_9089
timestamp 1677677812
transform 1 0 1672 0 -1 970
box -8 -3 16 105
use FILL  FILL_9090
timestamp 1677677812
transform 1 0 1680 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7304
timestamp 1677677812
transform 1 0 1700 0 1 875
box -3 -3 3 3
use FILL  FILL_9091
timestamp 1677677812
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_9092
timestamp 1677677812
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_341
timestamp 1677677812
transform 1 0 1704 0 -1 970
box -8 -3 46 105
use FILL  FILL_9093
timestamp 1677677812
transform 1 0 1744 0 -1 970
box -8 -3 16 105
use FILL  FILL_9094
timestamp 1677677812
transform 1 0 1752 0 -1 970
box -8 -3 16 105
use FILL  FILL_9095
timestamp 1677677812
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_9096
timestamp 1677677812
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use FILL  FILL_9097
timestamp 1677677812
transform 1 0 1776 0 -1 970
box -8 -3 16 105
use FILL  FILL_9098
timestamp 1677677812
transform 1 0 1784 0 -1 970
box -8 -3 16 105
use FILL  FILL_9112
timestamp 1677677812
transform 1 0 1792 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_494
timestamp 1677677812
transform -1 0 1896 0 -1 970
box -8 -3 104 105
use FILL  FILL_9113
timestamp 1677677812
transform 1 0 1896 0 -1 970
box -8 -3 16 105
use FILL  FILL_9114
timestamp 1677677812
transform 1 0 1904 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7305
timestamp 1677677812
transform 1 0 1972 0 1 875
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_495
timestamp 1677677812
transform -1 0 2008 0 -1 970
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_496
timestamp 1677677812
transform -1 0 2104 0 -1 970
box -8 -3 104 105
use FILL  FILL_9115
timestamp 1677677812
transform 1 0 2104 0 -1 970
box -8 -3 16 105
use FILL  FILL_9116
timestamp 1677677812
transform 1 0 2112 0 -1 970
box -8 -3 16 105
use FILL  FILL_9117
timestamp 1677677812
transform 1 0 2120 0 -1 970
box -8 -3 16 105
use FILL  FILL_9118
timestamp 1677677812
transform 1 0 2128 0 -1 970
box -8 -3 16 105
use FILL  FILL_9119
timestamp 1677677812
transform 1 0 2136 0 -1 970
box -8 -3 16 105
use FILL  FILL_9123
timestamp 1677677812
transform 1 0 2144 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_70
timestamp 1677677812
transform -1 0 2184 0 -1 970
box -8 -3 40 105
use FILL  FILL_9124
timestamp 1677677812
transform 1 0 2184 0 -1 970
box -8 -3 16 105
use FILL  FILL_9125
timestamp 1677677812
transform 1 0 2192 0 -1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_71
timestamp 1677677812
transform 1 0 2200 0 -1 970
box -8 -3 40 105
use FILL  FILL_9138
timestamp 1677677812
transform 1 0 2232 0 -1 970
box -8 -3 16 105
use FILL  FILL_9139
timestamp 1677677812
transform 1 0 2240 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_580
timestamp 1677677812
transform 1 0 2248 0 -1 970
box -9 -3 26 105
use INVX2  INVX2_581
timestamp 1677677812
transform -1 0 2280 0 -1 970
box -9 -3 26 105
use FILL  FILL_9140
timestamp 1677677812
transform 1 0 2280 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_23
timestamp 1677677812
transform 1 0 2288 0 -1 970
box -8 -3 32 105
use OAI21X1  OAI21X1_156
timestamp 1677677812
transform -1 0 2344 0 -1 970
box -8 -3 34 105
use FILL  FILL_9141
timestamp 1677677812
transform 1 0 2344 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7306
timestamp 1677677812
transform 1 0 2420 0 1 875
box -3 -3 3 3
use M3_M2  M3_M2_7307
timestamp 1677677812
transform 1 0 2476 0 1 875
box -3 -3 3 3
use FAX1  FAX1_16
timestamp 1677677812
transform -1 0 2472 0 -1 970
box -5 -3 126 105
use FILL  FILL_9142
timestamp 1677677812
transform 1 0 2472 0 -1 970
box -8 -3 16 105
use FILL  FILL_9143
timestamp 1677677812
transform 1 0 2480 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_583
timestamp 1677677812
transform -1 0 2504 0 -1 970
box -9 -3 26 105
use FILL  FILL_9145
timestamp 1677677812
transform 1 0 2504 0 -1 970
box -8 -3 16 105
use FILL  FILL_9146
timestamp 1677677812
transform 1 0 2512 0 -1 970
box -8 -3 16 105
use FILL  FILL_9147
timestamp 1677677812
transform 1 0 2520 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_53
timestamp 1677677812
transform 1 0 2528 0 -1 970
box -8 -3 40 105
use FILL  FILL_9148
timestamp 1677677812
transform 1 0 2560 0 -1 970
box -8 -3 16 105
use FILL  FILL_9151
timestamp 1677677812
transform 1 0 2568 0 -1 970
box -8 -3 16 105
use FILL  FILL_9152
timestamp 1677677812
transform 1 0 2576 0 -1 970
box -8 -3 16 105
use FILL  FILL_9153
timestamp 1677677812
transform 1 0 2584 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_342
timestamp 1677677812
transform 1 0 2592 0 -1 970
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_499
timestamp 1677677812
transform -1 0 2728 0 -1 970
box -8 -3 104 105
use FILL  FILL_9154
timestamp 1677677812
transform 1 0 2728 0 -1 970
box -8 -3 16 105
use FILL  FILL_9157
timestamp 1677677812
transform 1 0 2736 0 -1 970
box -8 -3 16 105
use FAX1  FAX1_19
timestamp 1677677812
transform 1 0 2744 0 -1 970
box -5 -3 126 105
use FILL  FILL_9158
timestamp 1677677812
transform 1 0 2864 0 -1 970
box -8 -3 16 105
use FILL  FILL_9159
timestamp 1677677812
transform 1 0 2872 0 -1 970
box -8 -3 16 105
use FILL  FILL_9160
timestamp 1677677812
transform 1 0 2880 0 -1 970
box -8 -3 16 105
use FILL  FILL_9161
timestamp 1677677812
transform 1 0 2888 0 -1 970
box -8 -3 16 105
use FILL  FILL_9162
timestamp 1677677812
transform 1 0 2896 0 -1 970
box -8 -3 16 105
use FILL  FILL_9163
timestamp 1677677812
transform 1 0 2904 0 -1 970
box -8 -3 16 105
use FILL  FILL_9164
timestamp 1677677812
transform 1 0 2912 0 -1 970
box -8 -3 16 105
use FILL  FILL_9165
timestamp 1677677812
transform 1 0 2920 0 -1 970
box -8 -3 16 105
use FILL  FILL_9166
timestamp 1677677812
transform 1 0 2928 0 -1 970
box -8 -3 16 105
use FILL  FILL_9167
timestamp 1677677812
transform 1 0 2936 0 -1 970
box -8 -3 16 105
use FILL  FILL_9168
timestamp 1677677812
transform 1 0 2944 0 -1 970
box -8 -3 16 105
use FILL  FILL_9169
timestamp 1677677812
transform 1 0 2952 0 -1 970
box -8 -3 16 105
use FILL  FILL_9170
timestamp 1677677812
transform 1 0 2960 0 -1 970
box -8 -3 16 105
use FILL  FILL_9171
timestamp 1677677812
transform 1 0 2968 0 -1 970
box -8 -3 16 105
use FILL  FILL_9172
timestamp 1677677812
transform 1 0 2976 0 -1 970
box -8 -3 16 105
use FILL  FILL_9173
timestamp 1677677812
transform 1 0 2984 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_26
timestamp 1677677812
transform 1 0 2992 0 -1 970
box -8 -3 32 105
use FILL  FILL_9176
timestamp 1677677812
transform 1 0 3016 0 -1 970
box -8 -3 16 105
use FILL  FILL_9177
timestamp 1677677812
transform 1 0 3024 0 -1 970
box -8 -3 16 105
use FILL  FILL_9178
timestamp 1677677812
transform 1 0 3032 0 -1 970
box -8 -3 16 105
use FILL  FILL_9179
timestamp 1677677812
transform 1 0 3040 0 -1 970
box -8 -3 16 105
use FILL  FILL_9180
timestamp 1677677812
transform 1 0 3048 0 -1 970
box -8 -3 16 105
use FILL  FILL_9189
timestamp 1677677812
transform 1 0 3056 0 -1 970
box -8 -3 16 105
use FILL  FILL_9190
timestamp 1677677812
transform 1 0 3064 0 -1 970
box -8 -3 16 105
use FILL  FILL_9191
timestamp 1677677812
transform 1 0 3072 0 -1 970
box -8 -3 16 105
use AOI21X1  AOI21X1_15
timestamp 1677677812
transform 1 0 3080 0 -1 970
box -7 -3 39 105
use FILL  FILL_9192
timestamp 1677677812
transform 1 0 3112 0 -1 970
box -8 -3 16 105
use FILL  FILL_9193
timestamp 1677677812
transform 1 0 3120 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_158
timestamp 1677677812
transform -1 0 3160 0 -1 970
box -8 -3 34 105
use NAND3X1  NAND3X1_72
timestamp 1677677812
transform -1 0 3192 0 -1 970
box -8 -3 40 105
use FILL  FILL_9194
timestamp 1677677812
transform 1 0 3192 0 -1 970
box -8 -3 16 105
use FILL  FILL_9199
timestamp 1677677812
transform 1 0 3200 0 -1 970
box -8 -3 16 105
use FILL  FILL_9200
timestamp 1677677812
transform 1 0 3208 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7308
timestamp 1677677812
transform 1 0 3228 0 1 875
box -3 -3 3 3
use FILL  FILL_9201
timestamp 1677677812
transform 1 0 3216 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_344
timestamp 1677677812
transform -1 0 3264 0 -1 970
box -8 -3 46 105
use FILL  FILL_9202
timestamp 1677677812
transform 1 0 3264 0 -1 970
box -8 -3 16 105
use FILL  FILL_9204
timestamp 1677677812
transform 1 0 3272 0 -1 970
box -8 -3 16 105
use FILL  FILL_9206
timestamp 1677677812
transform 1 0 3280 0 -1 970
box -8 -3 16 105
use FILL  FILL_9213
timestamp 1677677812
transform 1 0 3288 0 -1 970
box -8 -3 16 105
use FILL  FILL_9214
timestamp 1677677812
transform 1 0 3296 0 -1 970
box -8 -3 16 105
use FILL  FILL_9215
timestamp 1677677812
transform 1 0 3304 0 -1 970
box -8 -3 16 105
use FILL  FILL_9216
timestamp 1677677812
transform 1 0 3312 0 -1 970
box -8 -3 16 105
use AOI22X1  AOI22X1_346
timestamp 1677677812
transform -1 0 3360 0 -1 970
box -8 -3 46 105
use FILL  FILL_9217
timestamp 1677677812
transform 1 0 3360 0 -1 970
box -8 -3 16 105
use FILL  FILL_9218
timestamp 1677677812
transform 1 0 3368 0 -1 970
box -8 -3 16 105
use FAX1  FAX1_21
timestamp 1677677812
transform -1 0 3496 0 -1 970
box -5 -3 126 105
use FILL  FILL_9219
timestamp 1677677812
transform 1 0 3496 0 -1 970
box -8 -3 16 105
use FILL  FILL_9220
timestamp 1677677812
transform 1 0 3504 0 -1 970
box -8 -3 16 105
use FILL  FILL_9221
timestamp 1677677812
transform 1 0 3512 0 -1 970
box -8 -3 16 105
use FILL  FILL_9222
timestamp 1677677812
transform 1 0 3520 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_55
timestamp 1677677812
transform 1 0 3528 0 -1 970
box -8 -3 40 105
use FILL  FILL_9239
timestamp 1677677812
transform 1 0 3560 0 -1 970
box -8 -3 16 105
use FILL  FILL_9240
timestamp 1677677812
transform 1 0 3568 0 -1 970
box -8 -3 16 105
use FILL  FILL_9241
timestamp 1677677812
transform 1 0 3576 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_587
timestamp 1677677812
transform 1 0 3584 0 -1 970
box -9 -3 26 105
use M3_M2  M3_M2_7309
timestamp 1677677812
transform 1 0 3628 0 1 875
box -3 -3 3 3
use OAI21X1  OAI21X1_159
timestamp 1677677812
transform 1 0 3600 0 -1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_27
timestamp 1677677812
transform -1 0 3656 0 -1 970
box -8 -3 32 105
use FILL  FILL_9242
timestamp 1677677812
transform 1 0 3656 0 -1 970
box -8 -3 16 105
use FILL  FILL_9243
timestamp 1677677812
transform 1 0 3664 0 -1 970
box -8 -3 16 105
use FILL  FILL_9244
timestamp 1677677812
transform 1 0 3672 0 -1 970
box -8 -3 16 105
use FILL  FILL_9245
timestamp 1677677812
transform 1 0 3680 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_160
timestamp 1677677812
transform 1 0 3688 0 -1 970
box -8 -3 34 105
use FILL  FILL_9246
timestamp 1677677812
transform 1 0 3720 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_161
timestamp 1677677812
transform 1 0 3728 0 -1 970
box -8 -3 34 105
use FILL  FILL_9265
timestamp 1677677812
transform 1 0 3760 0 -1 970
box -8 -3 16 105
use FILL  FILL_9266
timestamp 1677677812
transform 1 0 3768 0 -1 970
box -8 -3 16 105
use FILL  FILL_9267
timestamp 1677677812
transform 1 0 3776 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_28
timestamp 1677677812
transform -1 0 3808 0 -1 970
box -8 -3 32 105
use FILL  FILL_9268
timestamp 1677677812
transform 1 0 3808 0 -1 970
box -8 -3 16 105
use FILL  FILL_9269
timestamp 1677677812
transform 1 0 3816 0 -1 970
box -8 -3 16 105
use FILL  FILL_9270
timestamp 1677677812
transform 1 0 3824 0 -1 970
box -8 -3 16 105
use FILL  FILL_9271
timestamp 1677677812
transform 1 0 3832 0 -1 970
box -8 -3 16 105
use FILL  FILL_9272
timestamp 1677677812
transform 1 0 3840 0 -1 970
box -8 -3 16 105
use FILL  FILL_9273
timestamp 1677677812
transform 1 0 3848 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_29
timestamp 1677677812
transform 1 0 3856 0 -1 970
box -8 -3 32 105
use FILL  FILL_9274
timestamp 1677677812
transform 1 0 3880 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7310
timestamp 1677677812
transform 1 0 3900 0 1 875
box -3 -3 3 3
use FILL  FILL_9275
timestamp 1677677812
transform 1 0 3888 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_162
timestamp 1677677812
transform -1 0 3928 0 -1 970
box -8 -3 34 105
use FILL  FILL_9276
timestamp 1677677812
transform 1 0 3928 0 -1 970
box -8 -3 16 105
use FILL  FILL_9277
timestamp 1677677812
transform 1 0 3936 0 -1 970
box -8 -3 16 105
use FILL  FILL_9278
timestamp 1677677812
transform 1 0 3944 0 -1 970
box -8 -3 16 105
use FILL  FILL_9279
timestamp 1677677812
transform 1 0 3952 0 -1 970
box -8 -3 16 105
use FILL  FILL_9280
timestamp 1677677812
transform 1 0 3960 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_163
timestamp 1677677812
transform 1 0 3968 0 -1 970
box -8 -3 34 105
use FILL  FILL_9281
timestamp 1677677812
transform 1 0 4000 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_30
timestamp 1677677812
transform -1 0 4032 0 -1 970
box -8 -3 32 105
use FILL  FILL_9282
timestamp 1677677812
transform 1 0 4032 0 -1 970
box -8 -3 16 105
use FILL  FILL_9283
timestamp 1677677812
transform 1 0 4040 0 -1 970
box -8 -3 16 105
use M3_M2  M3_M2_7311
timestamp 1677677812
transform 1 0 4076 0 1 875
box -3 -3 3 3
use OAI21X1  OAI21X1_164
timestamp 1677677812
transform 1 0 4048 0 -1 970
box -8 -3 34 105
use FILL  FILL_9284
timestamp 1677677812
transform 1 0 4080 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_31
timestamp 1677677812
transform -1 0 4112 0 -1 970
box -8 -3 32 105
use FILL  FILL_9285
timestamp 1677677812
transform 1 0 4112 0 -1 970
box -8 -3 16 105
use FILL  FILL_9286
timestamp 1677677812
transform 1 0 4120 0 -1 970
box -8 -3 16 105
use FILL  FILL_9288
timestamp 1677677812
transform 1 0 4128 0 -1 970
box -8 -3 16 105
use FILL  FILL_9290
timestamp 1677677812
transform 1 0 4136 0 -1 970
box -8 -3 16 105
use FILL  FILL_9292
timestamp 1677677812
transform 1 0 4144 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_165
timestamp 1677677812
transform 1 0 4152 0 -1 970
box -8 -3 34 105
use FILL  FILL_9295
timestamp 1677677812
transform 1 0 4184 0 -1 970
box -8 -3 16 105
use FILL  FILL_9296
timestamp 1677677812
transform 1 0 4192 0 -1 970
box -8 -3 16 105
use FILL  FILL_9297
timestamp 1677677812
transform 1 0 4200 0 -1 970
box -8 -3 16 105
use FILL  FILL_9299
timestamp 1677677812
transform 1 0 4208 0 -1 970
box -8 -3 16 105
use FILL  FILL_9302
timestamp 1677677812
transform 1 0 4216 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_166
timestamp 1677677812
transform -1 0 4256 0 -1 970
box -8 -3 34 105
use FILL  FILL_9303
timestamp 1677677812
transform 1 0 4256 0 -1 970
box -8 -3 16 105
use FILL  FILL_9304
timestamp 1677677812
transform 1 0 4264 0 -1 970
box -8 -3 16 105
use FILL  FILL_9322
timestamp 1677677812
transform 1 0 4272 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_168
timestamp 1677677812
transform -1 0 4312 0 -1 970
box -8 -3 34 105
use FILL  FILL_9323
timestamp 1677677812
transform 1 0 4312 0 -1 970
box -8 -3 16 105
use FILL  FILL_9324
timestamp 1677677812
transform 1 0 4320 0 -1 970
box -8 -3 16 105
use FILL  FILL_9325
timestamp 1677677812
transform 1 0 4328 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_169
timestamp 1677677812
transform -1 0 4368 0 -1 970
box -8 -3 34 105
use FILL  FILL_9326
timestamp 1677677812
transform 1 0 4368 0 -1 970
box -8 -3 16 105
use FILL  FILL_9327
timestamp 1677677812
transform 1 0 4376 0 -1 970
box -8 -3 16 105
use FILL  FILL_9328
timestamp 1677677812
transform 1 0 4384 0 -1 970
box -8 -3 16 105
use FILL  FILL_9329
timestamp 1677677812
transform 1 0 4392 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_170
timestamp 1677677812
transform -1 0 4432 0 -1 970
box -8 -3 34 105
use OAI22X1  OAI22X1_351
timestamp 1677677812
transform -1 0 4472 0 -1 970
box -8 -3 46 105
use FILL  FILL_9330
timestamp 1677677812
transform 1 0 4472 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_171
timestamp 1677677812
transform -1 0 4512 0 -1 970
box -8 -3 34 105
use FILL  FILL_9331
timestamp 1677677812
transform 1 0 4512 0 -1 970
box -8 -3 16 105
use FILL  FILL_9332
timestamp 1677677812
transform 1 0 4520 0 -1 970
box -8 -3 16 105
use FILL  FILL_9333
timestamp 1677677812
transform 1 0 4528 0 -1 970
box -8 -3 16 105
use FILL  FILL_9335
timestamp 1677677812
transform 1 0 4536 0 -1 970
box -8 -3 16 105
use FILL  FILL_9338
timestamp 1677677812
transform 1 0 4544 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_353
timestamp 1677677812
transform 1 0 4552 0 -1 970
box -8 -3 46 105
use FILL  FILL_9339
timestamp 1677677812
transform 1 0 4592 0 -1 970
box -8 -3 16 105
use FILL  FILL_9341
timestamp 1677677812
transform 1 0 4600 0 -1 970
box -8 -3 16 105
use FILL  FILL_9343
timestamp 1677677812
transform 1 0 4608 0 -1 970
box -8 -3 16 105
use FILL  FILL_9345
timestamp 1677677812
transform 1 0 4616 0 -1 970
box -8 -3 16 105
use FILL  FILL_9357
timestamp 1677677812
transform 1 0 4624 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_172
timestamp 1677677812
transform -1 0 4664 0 -1 970
box -8 -3 34 105
use FILL  FILL_9358
timestamp 1677677812
transform 1 0 4664 0 -1 970
box -8 -3 16 105
use FILL  FILL_9359
timestamp 1677677812
transform 1 0 4672 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_501
timestamp 1677677812
transform 1 0 4680 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_589
timestamp 1677677812
transform -1 0 4792 0 -1 970
box -9 -3 26 105
use top_level_VIA0  top_level_VIA0_77
timestamp 1677677812
transform 1 0 4843 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_7361
timestamp 1677677812
transform 1 0 132 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7362
timestamp 1677677812
transform 1 0 172 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8187
timestamp 1677677812
transform 1 0 132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8188
timestamp 1677677812
transform 1 0 164 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8189
timestamp 1677677812
transform 1 0 172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8312
timestamp 1677677812
transform 1 0 84 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7447
timestamp 1677677812
transform 1 0 164 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7363
timestamp 1677677812
transform 1 0 204 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8313
timestamp 1677677812
transform 1 0 204 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8314
timestamp 1677677812
transform 1 0 212 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7331
timestamp 1677677812
transform 1 0 236 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7364
timestamp 1677677812
transform 1 0 244 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8190
timestamp 1677677812
transform 1 0 220 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8191
timestamp 1677677812
transform 1 0 228 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7402
timestamp 1677677812
transform 1 0 236 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8192
timestamp 1677677812
transform 1 0 244 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7403
timestamp 1677677812
transform 1 0 252 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7332
timestamp 1677677812
transform 1 0 268 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8193
timestamp 1677677812
transform 1 0 260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8194
timestamp 1677677812
transform 1 0 268 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8315
timestamp 1677677812
transform 1 0 228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8316
timestamp 1677677812
transform 1 0 252 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7448
timestamp 1677677812
transform 1 0 228 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7428
timestamp 1677677812
transform 1 0 260 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8317
timestamp 1677677812
transform 1 0 276 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7429
timestamp 1677677812
transform 1 0 324 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8195
timestamp 1677677812
transform 1 0 364 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7404
timestamp 1677677812
transform 1 0 372 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8318
timestamp 1677677812
transform 1 0 372 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8196
timestamp 1677677812
transform 1 0 404 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8319
timestamp 1677677812
transform 1 0 412 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7333
timestamp 1677677812
transform 1 0 436 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8197
timestamp 1677677812
transform 1 0 436 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7365
timestamp 1677677812
transform 1 0 500 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7366
timestamp 1677677812
transform 1 0 540 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8198
timestamp 1677677812
transform 1 0 500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8199
timestamp 1677677812
transform 1 0 532 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8200
timestamp 1677677812
transform 1 0 540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8320
timestamp 1677677812
transform 1 0 452 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7430
timestamp 1677677812
transform 1 0 532 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7367
timestamp 1677677812
transform 1 0 556 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8321
timestamp 1677677812
transform 1 0 548 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8322
timestamp 1677677812
transform 1 0 556 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7431
timestamp 1677677812
transform 1 0 572 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7334
timestamp 1677677812
transform 1 0 588 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7368
timestamp 1677677812
transform 1 0 604 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8201
timestamp 1677677812
transform 1 0 580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8202
timestamp 1677677812
transform 1 0 588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8203
timestamp 1677677812
transform 1 0 604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8204
timestamp 1677677812
transform 1 0 620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8323
timestamp 1677677812
transform 1 0 588 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7369
timestamp 1677677812
transform 1 0 652 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7405
timestamp 1677677812
transform 1 0 644 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8205
timestamp 1677677812
transform 1 0 652 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7406
timestamp 1677677812
transform 1 0 660 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8324
timestamp 1677677812
transform 1 0 636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8325
timestamp 1677677812
transform 1 0 644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8326
timestamp 1677677812
transform 1 0 660 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8327
timestamp 1677677812
transform 1 0 676 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7449
timestamp 1677677812
transform 1 0 636 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8328
timestamp 1677677812
transform 1 0 692 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7482
timestamp 1677677812
transform 1 0 684 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7316
timestamp 1677677812
transform 1 0 748 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_7370
timestamp 1677677812
transform 1 0 748 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8206
timestamp 1677677812
transform 1 0 708 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8207
timestamp 1677677812
transform 1 0 716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8208
timestamp 1677677812
transform 1 0 748 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8329
timestamp 1677677812
transform 1 0 724 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8330
timestamp 1677677812
transform 1 0 740 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7450
timestamp 1677677812
transform 1 0 724 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8209
timestamp 1677677812
transform 1 0 764 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8210
timestamp 1677677812
transform 1 0 812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8331
timestamp 1677677812
transform 1 0 780 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8332
timestamp 1677677812
transform 1 0 788 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7451
timestamp 1677677812
transform 1 0 780 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7432
timestamp 1677677812
transform 1 0 796 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8333
timestamp 1677677812
transform 1 0 804 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7433
timestamp 1677677812
transform 1 0 812 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8211
timestamp 1677677812
transform 1 0 828 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7452
timestamp 1677677812
transform 1 0 820 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7483
timestamp 1677677812
transform 1 0 804 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8212
timestamp 1677677812
transform 1 0 852 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8334
timestamp 1677677812
transform 1 0 836 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8335
timestamp 1677677812
transform 1 0 844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8336
timestamp 1677677812
transform 1 0 860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8337
timestamp 1677677812
transform 1 0 868 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7453
timestamp 1677677812
transform 1 0 844 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7484
timestamp 1677677812
transform 1 0 836 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7485
timestamp 1677677812
transform 1 0 860 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7371
timestamp 1677677812
transform 1 0 884 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8213
timestamp 1677677812
transform 1 0 884 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7454
timestamp 1677677812
transform 1 0 892 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8214
timestamp 1677677812
transform 1 0 908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8215
timestamp 1677677812
transform 1 0 916 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8216
timestamp 1677677812
transform 1 0 972 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8338
timestamp 1677677812
transform 1 0 996 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7434
timestamp 1677677812
transform 1 0 1012 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8430
timestamp 1677677812
transform 1 0 1012 0 1 795
box -2 -2 2 2
use M2_M1  M2_M1_8217
timestamp 1677677812
transform 1 0 1060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8339
timestamp 1677677812
transform 1 0 1052 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7407
timestamp 1677677812
transform 1 0 1068 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8340
timestamp 1677677812
transform 1 0 1068 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7455
timestamp 1677677812
transform 1 0 1068 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7372
timestamp 1677677812
transform 1 0 1084 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7373
timestamp 1677677812
transform 1 0 1124 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8218
timestamp 1677677812
transform 1 0 1084 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8219
timestamp 1677677812
transform 1 0 1124 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7408
timestamp 1677677812
transform 1 0 1132 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8341
timestamp 1677677812
transform 1 0 1100 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8220
timestamp 1677677812
transform 1 0 1196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8342
timestamp 1677677812
transform 1 0 1188 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7335
timestamp 1677677812
transform 1 0 1212 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8221
timestamp 1677677812
transform 1 0 1212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8222
timestamp 1677677812
transform 1 0 1228 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8223
timestamp 1677677812
transform 1 0 1244 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7486
timestamp 1677677812
transform 1 0 1236 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8343
timestamp 1677677812
transform 1 0 1260 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7435
timestamp 1677677812
transform 1 0 1268 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8344
timestamp 1677677812
transform 1 0 1276 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8345
timestamp 1677677812
transform 1 0 1284 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7456
timestamp 1677677812
transform 1 0 1260 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8431
timestamp 1677677812
transform 1 0 1268 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7457
timestamp 1677677812
transform 1 0 1284 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7487
timestamp 1677677812
transform 1 0 1284 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7312
timestamp 1677677812
transform 1 0 1316 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_8346
timestamp 1677677812
transform 1 0 1308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8224
timestamp 1677677812
transform 1 0 1316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8225
timestamp 1677677812
transform 1 0 1332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8226
timestamp 1677677812
transform 1 0 1348 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8347
timestamp 1677677812
transform 1 0 1340 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7320
timestamp 1677677812
transform 1 0 1436 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7336
timestamp 1677677812
transform 1 0 1436 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8227
timestamp 1677677812
transform 1 0 1396 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8228
timestamp 1677677812
transform 1 0 1444 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8348
timestamp 1677677812
transform 1 0 1476 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7337
timestamp 1677677812
transform 1 0 1580 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7374
timestamp 1677677812
transform 1 0 1548 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7375
timestamp 1677677812
transform 1 0 1588 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8229
timestamp 1677677812
transform 1 0 1548 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8230
timestamp 1677677812
transform 1 0 1580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8231
timestamp 1677677812
transform 1 0 1588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8349
timestamp 1677677812
transform 1 0 1500 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7458
timestamp 1677677812
transform 1 0 1500 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7459
timestamp 1677677812
transform 1 0 1532 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8232
timestamp 1677677812
transform 1 0 1628 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7321
timestamp 1677677812
transform 1 0 1676 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7338
timestamp 1677677812
transform 1 0 1644 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7339
timestamp 1677677812
transform 1 0 1668 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8233
timestamp 1677677812
transform 1 0 1652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8234
timestamp 1677677812
transform 1 0 1668 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8235
timestamp 1677677812
transform 1 0 1676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8350
timestamp 1677677812
transform 1 0 1636 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8351
timestamp 1677677812
transform 1 0 1644 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8352
timestamp 1677677812
transform 1 0 1660 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7488
timestamp 1677677812
transform 1 0 1628 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7489
timestamp 1677677812
transform 1 0 1652 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8353
timestamp 1677677812
transform 1 0 1708 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7313
timestamp 1677677812
transform 1 0 1724 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_8236
timestamp 1677677812
transform 1 0 1732 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7409
timestamp 1677677812
transform 1 0 1740 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8237
timestamp 1677677812
transform 1 0 1756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8354
timestamp 1677677812
transform 1 0 1740 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8355
timestamp 1677677812
transform 1 0 1748 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7322
timestamp 1677677812
transform 1 0 1844 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7376
timestamp 1677677812
transform 1 0 1788 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7377
timestamp 1677677812
transform 1 0 1828 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8238
timestamp 1677677812
transform 1 0 1788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8239
timestamp 1677677812
transform 1 0 1796 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7410
timestamp 1677677812
transform 1 0 1804 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8240
timestamp 1677677812
transform 1 0 1828 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8356
timestamp 1677677812
transform 1 0 1876 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7323
timestamp 1677677812
transform 1 0 1940 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8241
timestamp 1677677812
transform 1 0 1908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8242
timestamp 1677677812
transform 1 0 1924 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7411
timestamp 1677677812
transform 1 0 1932 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8243
timestamp 1677677812
transform 1 0 1940 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8357
timestamp 1677677812
transform 1 0 1900 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7436
timestamp 1677677812
transform 1 0 1908 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7412
timestamp 1677677812
transform 1 0 1948 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8244
timestamp 1677677812
transform 1 0 1956 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8245
timestamp 1677677812
transform 1 0 1964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8358
timestamp 1677677812
transform 1 0 1932 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8359
timestamp 1677677812
transform 1 0 1940 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8246
timestamp 1677677812
transform 1 0 1980 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8360
timestamp 1677677812
transform 1 0 1972 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7437
timestamp 1677677812
transform 1 0 1980 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7340
timestamp 1677677812
transform 1 0 2028 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7378
timestamp 1677677812
transform 1 0 2012 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8247
timestamp 1677677812
transform 1 0 2012 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7413
timestamp 1677677812
transform 1 0 2020 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7379
timestamp 1677677812
transform 1 0 2036 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8248
timestamp 1677677812
transform 1 0 2028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8361
timestamp 1677677812
transform 1 0 2020 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8249
timestamp 1677677812
transform 1 0 2044 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8362
timestamp 1677677812
transform 1 0 2036 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7341
timestamp 1677677812
transform 1 0 2076 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8250
timestamp 1677677812
transform 1 0 2124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8251
timestamp 1677677812
transform 1 0 2180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8252
timestamp 1677677812
transform 1 0 2188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8363
timestamp 1677677812
transform 1 0 2100 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8364
timestamp 1677677812
transform 1 0 2196 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7490
timestamp 1677677812
transform 1 0 2196 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7317
timestamp 1677677812
transform 1 0 2236 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8253
timestamp 1677677812
transform 1 0 2276 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7438
timestamp 1677677812
transform 1 0 2212 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7414
timestamp 1677677812
transform 1 0 2308 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7342
timestamp 1677677812
transform 1 0 2332 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8180
timestamp 1677677812
transform 1 0 2332 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8254
timestamp 1677677812
transform 1 0 2316 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8255
timestamp 1677677812
transform 1 0 2324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8365
timestamp 1677677812
transform 1 0 2228 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8366
timestamp 1677677812
transform 1 0 2316 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7491
timestamp 1677677812
transform 1 0 2300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7415
timestamp 1677677812
transform 1 0 2332 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7343
timestamp 1677677812
transform 1 0 2372 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7416
timestamp 1677677812
transform 1 0 2380 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7344
timestamp 1677677812
transform 1 0 2436 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7345
timestamp 1677677812
transform 1 0 2492 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8256
timestamp 1677677812
transform 1 0 2540 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8367
timestamp 1677677812
transform 1 0 2444 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7439
timestamp 1677677812
transform 1 0 2508 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8368
timestamp 1677677812
transform 1 0 2556 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8432
timestamp 1677677812
transform 1 0 2452 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7492
timestamp 1677677812
transform 1 0 2556 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7380
timestamp 1677677812
transform 1 0 2580 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8257
timestamp 1677677812
transform 1 0 2580 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8258
timestamp 1677677812
transform 1 0 2588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8259
timestamp 1677677812
transform 1 0 2604 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8369
timestamp 1677677812
transform 1 0 2572 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8370
timestamp 1677677812
transform 1 0 2588 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8371
timestamp 1677677812
transform 1 0 2612 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7346
timestamp 1677677812
transform 1 0 2628 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7381
timestamp 1677677812
transform 1 0 2628 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8260
timestamp 1677677812
transform 1 0 2628 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8372
timestamp 1677677812
transform 1 0 2636 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7382
timestamp 1677677812
transform 1 0 2700 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8261
timestamp 1677677812
transform 1 0 2700 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8373
timestamp 1677677812
transform 1 0 2724 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7324
timestamp 1677677812
transform 1 0 2748 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7347
timestamp 1677677812
transform 1 0 2740 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7383
timestamp 1677677812
transform 1 0 2748 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8262
timestamp 1677677812
transform 1 0 2740 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7493
timestamp 1677677812
transform 1 0 2732 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7325
timestamp 1677677812
transform 1 0 2852 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7384
timestamp 1677677812
transform 1 0 2812 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8263
timestamp 1677677812
transform 1 0 2812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8264
timestamp 1677677812
transform 1 0 2852 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7417
timestamp 1677677812
transform 1 0 2860 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8265
timestamp 1677677812
transform 1 0 2876 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7418
timestamp 1677677812
transform 1 0 2900 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8374
timestamp 1677677812
transform 1 0 2836 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8375
timestamp 1677677812
transform 1 0 2852 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7494
timestamp 1677677812
transform 1 0 2836 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7495
timestamp 1677677812
transform 1 0 2852 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7385
timestamp 1677677812
transform 1 0 2980 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8376
timestamp 1677677812
transform 1 0 2972 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8377
timestamp 1677677812
transform 1 0 2980 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7460
timestamp 1677677812
transform 1 0 2948 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8433
timestamp 1677677812
transform 1 0 2964 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_7461
timestamp 1677677812
transform 1 0 3028 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8181
timestamp 1677677812
transform 1 0 3044 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7386
timestamp 1677677812
transform 1 0 3060 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7419
timestamp 1677677812
transform 1 0 3052 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8266
timestamp 1677677812
transform 1 0 3060 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8267
timestamp 1677677812
transform 1 0 3068 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8378
timestamp 1677677812
transform 1 0 3052 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7496
timestamp 1677677812
transform 1 0 3052 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8182
timestamp 1677677812
transform 1 0 3092 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8179
timestamp 1677677812
transform 1 0 3108 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_7387
timestamp 1677677812
transform 1 0 3116 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8268
timestamp 1677677812
transform 1 0 3116 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7348
timestamp 1677677812
transform 1 0 3188 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8183
timestamp 1677677812
transform 1 0 3188 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7388
timestamp 1677677812
transform 1 0 3196 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8269
timestamp 1677677812
transform 1 0 3196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8270
timestamp 1677677812
transform 1 0 3212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8379
timestamp 1677677812
transform 1 0 3204 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7440
timestamp 1677677812
transform 1 0 3220 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8380
timestamp 1677677812
transform 1 0 3228 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7462
timestamp 1677677812
transform 1 0 3204 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7326
timestamp 1677677812
transform 1 0 3260 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7327
timestamp 1677677812
transform 1 0 3276 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_7349
timestamp 1677677812
transform 1 0 3276 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8271
timestamp 1677677812
transform 1 0 3260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8272
timestamp 1677677812
transform 1 0 3276 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7441
timestamp 1677677812
transform 1 0 3260 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8381
timestamp 1677677812
transform 1 0 3268 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8382
timestamp 1677677812
transform 1 0 3284 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8383
timestamp 1677677812
transform 1 0 3292 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7463
timestamp 1677677812
transform 1 0 3284 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7497
timestamp 1677677812
transform 1 0 3300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7464
timestamp 1677677812
transform 1 0 3316 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7389
timestamp 1677677812
transform 1 0 3356 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8273
timestamp 1677677812
transform 1 0 3332 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8274
timestamp 1677677812
transform 1 0 3356 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8384
timestamp 1677677812
transform 1 0 3332 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7465
timestamp 1677677812
transform 1 0 3332 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8385
timestamp 1677677812
transform 1 0 3380 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8386
timestamp 1677677812
transform 1 0 3388 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7498
timestamp 1677677812
transform 1 0 3356 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7466
timestamp 1677677812
transform 1 0 3388 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7328
timestamp 1677677812
transform 1 0 3420 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8275
timestamp 1677677812
transform 1 0 3420 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8276
timestamp 1677677812
transform 1 0 3476 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7420
timestamp 1677677812
transform 1 0 3492 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8277
timestamp 1677677812
transform 1 0 3500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8387
timestamp 1677677812
transform 1 0 3508 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8184
timestamp 1677677812
transform 1 0 3532 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7421
timestamp 1677677812
transform 1 0 3532 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8278
timestamp 1677677812
transform 1 0 3540 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7422
timestamp 1677677812
transform 1 0 3548 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8388
timestamp 1677677812
transform 1 0 3532 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7467
timestamp 1677677812
transform 1 0 3516 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7468
timestamp 1677677812
transform 1 0 3532 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8389
timestamp 1677677812
transform 1 0 3572 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7318
timestamp 1677677812
transform 1 0 3588 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8279
timestamp 1677677812
transform 1 0 3588 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8390
timestamp 1677677812
transform 1 0 3628 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7319
timestamp 1677677812
transform 1 0 3644 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_8280
timestamp 1677677812
transform 1 0 3652 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7469
timestamp 1677677812
transform 1 0 3668 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7350
timestamp 1677677812
transform 1 0 3692 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7390
timestamp 1677677812
transform 1 0 3692 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8281
timestamp 1677677812
transform 1 0 3684 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8282
timestamp 1677677812
transform 1 0 3700 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7351
timestamp 1677677812
transform 1 0 3740 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8185
timestamp 1677677812
transform 1 0 3724 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_8283
timestamp 1677677812
transform 1 0 3716 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8391
timestamp 1677677812
transform 1 0 3692 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8392
timestamp 1677677812
transform 1 0 3708 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7470
timestamp 1677677812
transform 1 0 3692 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7391
timestamp 1677677812
transform 1 0 3732 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8284
timestamp 1677677812
transform 1 0 3748 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7314
timestamp 1677677812
transform 1 0 3780 0 1 865
box -3 -3 3 3
use M2_M1  M2_M1_8285
timestamp 1677677812
transform 1 0 3812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8393
timestamp 1677677812
transform 1 0 3780 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8394
timestamp 1677677812
transform 1 0 3788 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8395
timestamp 1677677812
transform 1 0 3804 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7471
timestamp 1677677812
transform 1 0 3788 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7472
timestamp 1677677812
transform 1 0 3804 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7499
timestamp 1677677812
transform 1 0 3820 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8286
timestamp 1677677812
transform 1 0 3836 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7500
timestamp 1677677812
transform 1 0 3836 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7352
timestamp 1677677812
transform 1 0 3876 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7392
timestamp 1677677812
transform 1 0 3892 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8287
timestamp 1677677812
transform 1 0 3876 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8288
timestamp 1677677812
transform 1 0 3892 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8396
timestamp 1677677812
transform 1 0 3860 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8397
timestamp 1677677812
transform 1 0 3868 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8398
timestamp 1677677812
transform 1 0 3884 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7473
timestamp 1677677812
transform 1 0 3868 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7501
timestamp 1677677812
transform 1 0 3860 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7353
timestamp 1677677812
transform 1 0 3908 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8289
timestamp 1677677812
transform 1 0 3908 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8399
timestamp 1677677812
transform 1 0 3908 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7474
timestamp 1677677812
transform 1 0 3900 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7502
timestamp 1677677812
transform 1 0 3908 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7475
timestamp 1677677812
transform 1 0 3924 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7393
timestamp 1677677812
transform 1 0 3964 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8290
timestamp 1677677812
transform 1 0 3964 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8400
timestamp 1677677812
transform 1 0 3940 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7442
timestamp 1677677812
transform 1 0 3948 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8401
timestamp 1677677812
transform 1 0 3956 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7329
timestamp 1677677812
transform 1 0 4012 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8402
timestamp 1677677812
transform 1 0 4004 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7394
timestamp 1677677812
transform 1 0 4028 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8291
timestamp 1677677812
transform 1 0 4028 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8403
timestamp 1677677812
transform 1 0 4036 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7443
timestamp 1677677812
transform 1 0 4044 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8404
timestamp 1677677812
transform 1 0 4052 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7354
timestamp 1677677812
transform 1 0 4084 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8405
timestamp 1677677812
transform 1 0 4076 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8292
timestamp 1677677812
transform 1 0 4084 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8406
timestamp 1677677812
transform 1 0 4084 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7355
timestamp 1677677812
transform 1 0 4116 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7395
timestamp 1677677812
transform 1 0 4100 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8293
timestamp 1677677812
transform 1 0 4100 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8294
timestamp 1677677812
transform 1 0 4116 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8295
timestamp 1677677812
transform 1 0 4124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8407
timestamp 1677677812
transform 1 0 4108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8408
timestamp 1677677812
transform 1 0 4124 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8409
timestamp 1677677812
transform 1 0 4156 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8296
timestamp 1677677812
transform 1 0 4172 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8186
timestamp 1677677812
transform 1 0 4188 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_7396
timestamp 1677677812
transform 1 0 4204 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7423
timestamp 1677677812
transform 1 0 4196 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_7397
timestamp 1677677812
transform 1 0 4252 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7424
timestamp 1677677812
transform 1 0 4252 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8297
timestamp 1677677812
transform 1 0 4260 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8410
timestamp 1677677812
transform 1 0 4236 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8411
timestamp 1677677812
transform 1 0 4252 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8412
timestamp 1677677812
transform 1 0 4268 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7356
timestamp 1677677812
transform 1 0 4284 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8298
timestamp 1677677812
transform 1 0 4284 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7357
timestamp 1677677812
transform 1 0 4332 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7425
timestamp 1677677812
transform 1 0 4308 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8299
timestamp 1677677812
transform 1 0 4332 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7398
timestamp 1677677812
transform 1 0 4348 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8413
timestamp 1677677812
transform 1 0 4308 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8414
timestamp 1677677812
transform 1 0 4324 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8415
timestamp 1677677812
transform 1 0 4340 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7476
timestamp 1677677812
transform 1 0 4308 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7503
timestamp 1677677812
transform 1 0 4300 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7504
timestamp 1677677812
transform 1 0 4324 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7505
timestamp 1677677812
transform 1 0 4340 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8416
timestamp 1677677812
transform 1 0 4356 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7477
timestamp 1677677812
transform 1 0 4356 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8300
timestamp 1677677812
transform 1 0 4380 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8301
timestamp 1677677812
transform 1 0 4396 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7330
timestamp 1677677812
transform 1 0 4412 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_8302
timestamp 1677677812
transform 1 0 4412 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8417
timestamp 1677677812
transform 1 0 4388 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8418
timestamp 1677677812
transform 1 0 4404 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7506
timestamp 1677677812
transform 1 0 4404 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7399
timestamp 1677677812
transform 1 0 4420 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7358
timestamp 1677677812
transform 1 0 4468 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8303
timestamp 1677677812
transform 1 0 4452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8304
timestamp 1677677812
transform 1 0 4468 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8419
timestamp 1677677812
transform 1 0 4444 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7444
timestamp 1677677812
transform 1 0 4452 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_8420
timestamp 1677677812
transform 1 0 4460 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8421
timestamp 1677677812
transform 1 0 4476 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8422
timestamp 1677677812
transform 1 0 4484 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7478
timestamp 1677677812
transform 1 0 4444 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7315
timestamp 1677677812
transform 1 0 4492 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_7359
timestamp 1677677812
transform 1 0 4492 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_7479
timestamp 1677677812
transform 1 0 4484 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7507
timestamp 1677677812
transform 1 0 4476 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7400
timestamp 1677677812
transform 1 0 4532 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_8305
timestamp 1677677812
transform 1 0 4508 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8306
timestamp 1677677812
transform 1 0 4516 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8307
timestamp 1677677812
transform 1 0 4532 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_7445
timestamp 1677677812
transform 1 0 4508 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7426
timestamp 1677677812
transform 1 0 4540 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8423
timestamp 1677677812
transform 1 0 4524 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8424
timestamp 1677677812
transform 1 0 4540 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7508
timestamp 1677677812
transform 1 0 4540 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7401
timestamp 1677677812
transform 1 0 4564 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_7427
timestamp 1677677812
transform 1 0 4580 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_8425
timestamp 1677677812
transform 1 0 4604 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7360
timestamp 1677677812
transform 1 0 4636 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_8308
timestamp 1677677812
transform 1 0 4636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8309
timestamp 1677677812
transform 1 0 4652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8426
timestamp 1677677812
transform 1 0 4628 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_8427
timestamp 1677677812
transform 1 0 4644 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7480
timestamp 1677677812
transform 1 0 4620 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_7509
timestamp 1677677812
transform 1 0 4620 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_7446
timestamp 1677677812
transform 1 0 4652 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_7481
timestamp 1677677812
transform 1 0 4644 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_8428
timestamp 1677677812
transform 1 0 4676 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_7510
timestamp 1677677812
transform 1 0 4676 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_8310
timestamp 1677677812
transform 1 0 4732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8311
timestamp 1677677812
transform 1 0 4788 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_8429
timestamp 1677677812
transform 1 0 4708 0 1 805
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_78
timestamp 1677677812
transform 1 0 48 0 1 770
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_502
timestamp 1677677812
transform 1 0 72 0 1 770
box -8 -3 104 105
use FILL  FILL_9360
timestamp 1677677812
transform 1 0 168 0 1 770
box -8 -3 16 105
use INVX2  INVX2_590
timestamp 1677677812
transform -1 0 192 0 1 770
box -9 -3 26 105
use FILL  FILL_9361
timestamp 1677677812
transform 1 0 192 0 1 770
box -8 -3 16 105
use FILL  FILL_9364
timestamp 1677677812
transform 1 0 200 0 1 770
box -8 -3 16 105
use INVX2  INVX2_592
timestamp 1677677812
transform 1 0 208 0 1 770
box -9 -3 26 105
use AOI22X1  AOI22X1_347
timestamp 1677677812
transform -1 0 264 0 1 770
box -8 -3 46 105
use FILL  FILL_9366
timestamp 1677677812
transform 1 0 264 0 1 770
box -8 -3 16 105
use FILL  FILL_9367
timestamp 1677677812
transform 1 0 272 0 1 770
box -8 -3 16 105
use FILL  FILL_9372
timestamp 1677677812
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_9374
timestamp 1677677812
transform 1 0 288 0 1 770
box -8 -3 16 105
use FILL  FILL_9375
timestamp 1677677812
transform 1 0 296 0 1 770
box -8 -3 16 105
use FILL  FILL_9376
timestamp 1677677812
transform 1 0 304 0 1 770
box -8 -3 16 105
use FILL  FILL_9377
timestamp 1677677812
transform 1 0 312 0 1 770
box -8 -3 16 105
use FILL  FILL_9378
timestamp 1677677812
transform 1 0 320 0 1 770
box -8 -3 16 105
use FILL  FILL_9379
timestamp 1677677812
transform 1 0 328 0 1 770
box -8 -3 16 105
use FILL  FILL_9380
timestamp 1677677812
transform 1 0 336 0 1 770
box -8 -3 16 105
use FILL  FILL_9381
timestamp 1677677812
transform 1 0 344 0 1 770
box -8 -3 16 105
use FILL  FILL_9382
timestamp 1677677812
transform 1 0 352 0 1 770
box -8 -3 16 105
use FILL  FILL_9383
timestamp 1677677812
transform 1 0 360 0 1 770
box -8 -3 16 105
use FILL  FILL_9384
timestamp 1677677812
transform 1 0 368 0 1 770
box -8 -3 16 105
use FILL  FILL_9385
timestamp 1677677812
transform 1 0 376 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_348
timestamp 1677677812
transform -1 0 424 0 1 770
box -8 -3 46 105
use FILL  FILL_9386
timestamp 1677677812
transform 1 0 424 0 1 770
box -8 -3 16 105
use FILL  FILL_9387
timestamp 1677677812
transform 1 0 432 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_504
timestamp 1677677812
transform 1 0 440 0 1 770
box -8 -3 104 105
use INVX2  INVX2_593
timestamp 1677677812
transform -1 0 552 0 1 770
box -9 -3 26 105
use INVX2  INVX2_594
timestamp 1677677812
transform 1 0 552 0 1 770
box -9 -3 26 105
use FILL  FILL_9388
timestamp 1677677812
transform 1 0 568 0 1 770
box -8 -3 16 105
use FILL  FILL_9389
timestamp 1677677812
transform 1 0 576 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_351
timestamp 1677677812
transform 1 0 584 0 1 770
box -8 -3 46 105
use FILL  FILL_9401
timestamp 1677677812
transform 1 0 624 0 1 770
box -8 -3 16 105
use FILL  FILL_9402
timestamp 1677677812
transform 1 0 632 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_357
timestamp 1677677812
transform -1 0 680 0 1 770
box -8 -3 46 105
use FILL  FILL_9403
timestamp 1677677812
transform 1 0 680 0 1 770
box -8 -3 16 105
use BUFX2  BUFX2_108
timestamp 1677677812
transform -1 0 712 0 1 770
box -5 -3 28 105
use FILL  FILL_9404
timestamp 1677677812
transform 1 0 712 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7511
timestamp 1677677812
transform 1 0 748 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_358
timestamp 1677677812
transform 1 0 720 0 1 770
box -8 -3 46 105
use FILL  FILL_9405
timestamp 1677677812
transform 1 0 760 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7512
timestamp 1677677812
transform 1 0 780 0 1 775
box -3 -3 3 3
use FILL  FILL_9412
timestamp 1677677812
transform 1 0 768 0 1 770
box -8 -3 16 105
use FILL  FILL_9413
timestamp 1677677812
transform 1 0 776 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_359
timestamp 1677677812
transform 1 0 784 0 1 770
box -8 -3 46 105
use FILL  FILL_9414
timestamp 1677677812
transform 1 0 824 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_352
timestamp 1677677812
transform -1 0 872 0 1 770
box -8 -3 46 105
use FILL  FILL_9415
timestamp 1677677812
transform 1 0 872 0 1 770
box -8 -3 16 105
use FILL  FILL_9416
timestamp 1677677812
transform 1 0 880 0 1 770
box -8 -3 16 105
use FILL  FILL_9417
timestamp 1677677812
transform 1 0 888 0 1 770
box -8 -3 16 105
use INVX2  INVX2_598
timestamp 1677677812
transform 1 0 896 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_507
timestamp 1677677812
transform -1 0 1008 0 1 770
box -8 -3 104 105
use FILL  FILL_9418
timestamp 1677677812
transform 1 0 1008 0 1 770
box -8 -3 16 105
use FILL  FILL_9424
timestamp 1677677812
transform 1 0 1016 0 1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_92
timestamp 1677677812
transform 1 0 1024 0 1 770
box -8 -3 32 105
use FILL  FILL_9425
timestamp 1677677812
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_9428
timestamp 1677677812
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_9429
timestamp 1677677812
transform 1 0 1064 0 1 770
box -8 -3 16 105
use INVX2  INVX2_601
timestamp 1677677812
transform 1 0 1072 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_509
timestamp 1677677812
transform 1 0 1088 0 1 770
box -8 -3 104 105
use FILL  FILL_9430
timestamp 1677677812
transform 1 0 1184 0 1 770
box -8 -3 16 105
use FILL  FILL_9443
timestamp 1677677812
transform 1 0 1192 0 1 770
box -8 -3 16 105
use FILL  FILL_9445
timestamp 1677677812
transform 1 0 1200 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_354
timestamp 1677677812
transform 1 0 1208 0 1 770
box -8 -3 46 105
use FILL  FILL_9447
timestamp 1677677812
transform 1 0 1248 0 1 770
box -8 -3 16 105
use FILL  FILL_9449
timestamp 1677677812
transform 1 0 1256 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7513
timestamp 1677677812
transform 1 0 1276 0 1 775
box -3 -3 3 3
use NOR2X1  NOR2X1_95
timestamp 1677677812
transform 1 0 1264 0 1 770
box -8 -3 32 105
use FILL  FILL_9451
timestamp 1677677812
transform 1 0 1288 0 1 770
box -8 -3 16 105
use FILL  FILL_9452
timestamp 1677677812
transform 1 0 1296 0 1 770
box -8 -3 16 105
use FILL  FILL_9453
timestamp 1677677812
transform 1 0 1304 0 1 770
box -8 -3 16 105
use FILL  FILL_9454
timestamp 1677677812
transform 1 0 1312 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7514
timestamp 1677677812
transform 1 0 1332 0 1 775
box -3 -3 3 3
use OAI22X1  OAI22X1_361
timestamp 1677677812
transform -1 0 1360 0 1 770
box -8 -3 46 105
use FILL  FILL_9455
timestamp 1677677812
transform 1 0 1360 0 1 770
box -8 -3 16 105
use FILL  FILL_9456
timestamp 1677677812
transform 1 0 1368 0 1 770
box -8 -3 16 105
use FILL  FILL_9457
timestamp 1677677812
transform 1 0 1376 0 1 770
box -8 -3 16 105
use FILL  FILL_9458
timestamp 1677677812
transform 1 0 1384 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_510
timestamp 1677677812
transform -1 0 1488 0 1 770
box -8 -3 104 105
use M3_M2  M3_M2_7515
timestamp 1677677812
transform 1 0 1508 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_7516
timestamp 1677677812
transform 1 0 1540 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_511
timestamp 1677677812
transform 1 0 1488 0 1 770
box -8 -3 104 105
use INVX2  INVX2_603
timestamp 1677677812
transform -1 0 1600 0 1 770
box -9 -3 26 105
use FILL  FILL_9459
timestamp 1677677812
transform 1 0 1600 0 1 770
box -8 -3 16 105
use FILL  FILL_9460
timestamp 1677677812
transform 1 0 1608 0 1 770
box -8 -3 16 105
use FILL  FILL_9461
timestamp 1677677812
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_9462
timestamp 1677677812
transform 1 0 1624 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_356
timestamp 1677677812
transform -1 0 1672 0 1 770
box -8 -3 46 105
use FILL  FILL_9463
timestamp 1677677812
transform 1 0 1672 0 1 770
box -8 -3 16 105
use FILL  FILL_9464
timestamp 1677677812
transform 1 0 1680 0 1 770
box -8 -3 16 105
use FILL  FILL_9465
timestamp 1677677812
transform 1 0 1688 0 1 770
box -8 -3 16 105
use FILL  FILL_9466
timestamp 1677677812
transform 1 0 1696 0 1 770
box -8 -3 16 105
use FILL  FILL_9467
timestamp 1677677812
transform 1 0 1704 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_357
timestamp 1677677812
transform 1 0 1712 0 1 770
box -8 -3 46 105
use FILL  FILL_9468
timestamp 1677677812
transform 1 0 1752 0 1 770
box -8 -3 16 105
use FILL  FILL_9469
timestamp 1677677812
transform 1 0 1760 0 1 770
box -8 -3 16 105
use FILL  FILL_9470
timestamp 1677677812
transform 1 0 1768 0 1 770
box -8 -3 16 105
use INVX2  INVX2_604
timestamp 1677677812
transform 1 0 1776 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_512
timestamp 1677677812
transform -1 0 1888 0 1 770
box -8 -3 104 105
use FILL  FILL_9471
timestamp 1677677812
transform 1 0 1888 0 1 770
box -8 -3 16 105
use FILL  FILL_9472
timestamp 1677677812
transform 1 0 1896 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_358
timestamp 1677677812
transform -1 0 1944 0 1 770
box -8 -3 46 105
use FILL  FILL_9473
timestamp 1677677812
transform 1 0 1944 0 1 770
box -8 -3 16 105
use INVX2  INVX2_605
timestamp 1677677812
transform 1 0 1952 0 1 770
box -9 -3 26 105
use FILL  FILL_9474
timestamp 1677677812
transform 1 0 1968 0 1 770
box -8 -3 16 105
use FILL  FILL_9495
timestamp 1677677812
transform 1 0 1976 0 1 770
box -8 -3 16 105
use FILL  FILL_9497
timestamp 1677677812
transform 1 0 1984 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_361
timestamp 1677677812
transform -1 0 2032 0 1 770
box -8 -3 46 105
use FILL  FILL_9498
timestamp 1677677812
transform 1 0 2032 0 1 770
box -8 -3 16 105
use FILL  FILL_9506
timestamp 1677677812
transform 1 0 2040 0 1 770
box -8 -3 16 105
use FILL  FILL_9508
timestamp 1677677812
transform 1 0 2048 0 1 770
box -8 -3 16 105
use INVX2  INVX2_609
timestamp 1677677812
transform 1 0 2056 0 1 770
box -9 -3 26 105
use FILL  FILL_9510
timestamp 1677677812
transform 1 0 2072 0 1 770
box -8 -3 16 105
use FILL  FILL_9514
timestamp 1677677812
transform 1 0 2080 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_517
timestamp 1677677812
transform 1 0 2088 0 1 770
box -8 -3 104 105
use FILL  FILL_9515
timestamp 1677677812
transform 1 0 2184 0 1 770
box -8 -3 16 105
use FILL  FILL_9516
timestamp 1677677812
transform 1 0 2192 0 1 770
box -8 -3 16 105
use INVX2  INVX2_610
timestamp 1677677812
transform 1 0 2200 0 1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_518
timestamp 1677677812
transform 1 0 2216 0 1 770
box -8 -3 104 105
use NAND2X1  NAND2X1_32
timestamp 1677677812
transform 1 0 2312 0 1 770
box -8 -3 32 105
use FILL  FILL_9517
timestamp 1677677812
transform 1 0 2336 0 1 770
box -8 -3 16 105
use FILL  FILL_9523
timestamp 1677677812
transform 1 0 2344 0 1 770
box -8 -3 16 105
use FILL  FILL_9525
timestamp 1677677812
transform 1 0 2352 0 1 770
box -8 -3 16 105
use FILL  FILL_9527
timestamp 1677677812
transform 1 0 2360 0 1 770
box -8 -3 16 105
use FILL  FILL_9529
timestamp 1677677812
transform 1 0 2368 0 1 770
box -8 -3 16 105
use FILL  FILL_9531
timestamp 1677677812
transform 1 0 2376 0 1 770
box -8 -3 16 105
use FILL  FILL_9533
timestamp 1677677812
transform 1 0 2384 0 1 770
box -8 -3 16 105
use FILL  FILL_9535
timestamp 1677677812
transform 1 0 2392 0 1 770
box -8 -3 16 105
use FILL  FILL_9537
timestamp 1677677812
transform 1 0 2400 0 1 770
box -8 -3 16 105
use FILL  FILL_9539
timestamp 1677677812
transform 1 0 2408 0 1 770
box -8 -3 16 105
use FILL  FILL_9540
timestamp 1677677812
transform 1 0 2416 0 1 770
box -8 -3 16 105
use FILL  FILL_9541
timestamp 1677677812
transform 1 0 2424 0 1 770
box -8 -3 16 105
use FILL  FILL_9542
timestamp 1677677812
transform 1 0 2432 0 1 770
box -8 -3 16 105
use FAX1  FAX1_22
timestamp 1677677812
transform -1 0 2560 0 1 770
box -5 -3 126 105
use FILL  FILL_9543
timestamp 1677677812
transform 1 0 2560 0 1 770
box -8 -3 16 105
use FILL  FILL_9544
timestamp 1677677812
transform 1 0 2568 0 1 770
box -8 -3 16 105
use FILL  FILL_9545
timestamp 1677677812
transform 1 0 2576 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_362
timestamp 1677677812
transform 1 0 2584 0 1 770
box -8 -3 46 105
use FILL  FILL_9546
timestamp 1677677812
transform 1 0 2624 0 1 770
box -8 -3 16 105
use FILL  FILL_9547
timestamp 1677677812
transform 1 0 2632 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_521
timestamp 1677677812
transform -1 0 2736 0 1 770
box -8 -3 104 105
use FILL  FILL_9548
timestamp 1677677812
transform 1 0 2736 0 1 770
box -8 -3 16 105
use FILL  FILL_9549
timestamp 1677677812
transform 1 0 2744 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_522
timestamp 1677677812
transform -1 0 2848 0 1 770
box -8 -3 104 105
use FILL  FILL_9550
timestamp 1677677812
transform 1 0 2848 0 1 770
box -8 -3 16 105
use FAX1  FAX1_23
timestamp 1677677812
transform 1 0 2856 0 1 770
box -5 -3 126 105
use FILL  FILL_9572
timestamp 1677677812
transform 1 0 2976 0 1 770
box -8 -3 16 105
use FILL  FILL_9573
timestamp 1677677812
transform 1 0 2984 0 1 770
box -8 -3 16 105
use FILL  FILL_9574
timestamp 1677677812
transform 1 0 2992 0 1 770
box -8 -3 16 105
use FILL  FILL_9575
timestamp 1677677812
transform 1 0 3000 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_33
timestamp 1677677812
transform 1 0 3008 0 1 770
box -8 -3 32 105
use FILL  FILL_9576
timestamp 1677677812
transform 1 0 3032 0 1 770
box -8 -3 16 105
use FILL  FILL_9577
timestamp 1677677812
transform 1 0 3040 0 1 770
box -8 -3 16 105
use FILL  FILL_9578
timestamp 1677677812
transform 1 0 3048 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_7517
timestamp 1677677812
transform 1 0 3068 0 1 775
box -3 -3 3 3
use INVX2  INVX2_612
timestamp 1677677812
transform 1 0 3056 0 1 770
box -9 -3 26 105
use FILL  FILL_9579
timestamp 1677677812
transform 1 0 3072 0 1 770
box -8 -3 16 105
use FILL  FILL_9593
timestamp 1677677812
transform 1 0 3080 0 1 770
box -8 -3 16 105
use FILL  FILL_9595
timestamp 1677677812
transform 1 0 3088 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_73
timestamp 1677677812
transform -1 0 3128 0 1 770
box -8 -3 40 105
use FILL  FILL_9596
timestamp 1677677812
transform 1 0 3128 0 1 770
box -8 -3 16 105
use FILL  FILL_9599
timestamp 1677677812
transform 1 0 3136 0 1 770
box -8 -3 16 105
use FILL  FILL_9601
timestamp 1677677812
transform 1 0 3144 0 1 770
box -8 -3 16 105
use FILL  FILL_9603
timestamp 1677677812
transform 1 0 3152 0 1 770
box -8 -3 16 105
use FILL  FILL_9604
timestamp 1677677812
transform 1 0 3160 0 1 770
box -8 -3 16 105
use FILL  FILL_9605
timestamp 1677677812
transform 1 0 3168 0 1 770
box -8 -3 16 105
use FILL  FILL_9606
timestamp 1677677812
transform 1 0 3176 0 1 770
box -8 -3 16 105
use FILL  FILL_9607
timestamp 1677677812
transform 1 0 3184 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_364
timestamp 1677677812
transform -1 0 3232 0 1 770
box -8 -3 46 105
use M3_M2  M3_M2_7518
timestamp 1677677812
transform 1 0 3244 0 1 775
box -3 -3 3 3
use FILL  FILL_9608
timestamp 1677677812
transform 1 0 3232 0 1 770
box -8 -3 16 105
use FILL  FILL_9609
timestamp 1677677812
transform 1 0 3240 0 1 770
box -8 -3 16 105
use FILL  FILL_9610
timestamp 1677677812
transform 1 0 3248 0 1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_365
timestamp 1677677812
transform 1 0 3256 0 1 770
box -8 -3 46 105
use FILL  FILL_9614
timestamp 1677677812
transform 1 0 3296 0 1 770
box -8 -3 16 105
use FILL  FILL_9615
timestamp 1677677812
transform 1 0 3304 0 1 770
box -8 -3 16 105
use FILL  FILL_9616
timestamp 1677677812
transform 1 0 3312 0 1 770
box -8 -3 16 105
use FILL  FILL_9617
timestamp 1677677812
transform 1 0 3320 0 1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_4
timestamp 1677677812
transform 1 0 3328 0 1 770
box -8 -3 64 105
use FILL  FILL_9618
timestamp 1677677812
transform 1 0 3384 0 1 770
box -8 -3 16 105
use FILL  FILL_9619
timestamp 1677677812
transform 1 0 3392 0 1 770
box -8 -3 16 105
use FILL  FILL_9620
timestamp 1677677812
transform 1 0 3400 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_59
timestamp 1677677812
transform 1 0 3408 0 1 770
box -8 -3 40 105
use FILL  FILL_9621
timestamp 1677677812
transform 1 0 3440 0 1 770
box -8 -3 16 105
use FILL  FILL_9622
timestamp 1677677812
transform 1 0 3448 0 1 770
box -8 -3 16 105
use FILL  FILL_9623
timestamp 1677677812
transform 1 0 3456 0 1 770
box -8 -3 16 105
use FILL  FILL_9624
timestamp 1677677812
transform 1 0 3464 0 1 770
box -8 -3 16 105
use FILL  FILL_9625
timestamp 1677677812
transform 1 0 3472 0 1 770
box -8 -3 16 105
use FILL  FILL_9626
timestamp 1677677812
transform 1 0 3480 0 1 770
box -8 -3 16 105
use FILL  FILL_9627
timestamp 1677677812
transform 1 0 3488 0 1 770
box -8 -3 16 105
use FILL  FILL_9628
timestamp 1677677812
transform 1 0 3496 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_36
timestamp 1677677812
transform 1 0 3504 0 1 770
box -8 -3 32 105
use AND2X2  AND2X2_60
timestamp 1677677812
transform 1 0 3528 0 1 770
box -8 -3 40 105
use FILL  FILL_9629
timestamp 1677677812
transform 1 0 3560 0 1 770
box -8 -3 16 105
use FILL  FILL_9635
timestamp 1677677812
transform 1 0 3568 0 1 770
box -8 -3 16 105
use FILL  FILL_9637
timestamp 1677677812
transform 1 0 3576 0 1 770
box -8 -3 16 105
use FILL  FILL_9639
timestamp 1677677812
transform 1 0 3584 0 1 770
box -8 -3 16 105
use FILL  FILL_9641
timestamp 1677677812
transform 1 0 3592 0 1 770
box -8 -3 16 105
use INVX2  INVX2_615
timestamp 1677677812
transform 1 0 3600 0 1 770
box -9 -3 26 105
use FILL  FILL_9642
timestamp 1677677812
transform 1 0 3616 0 1 770
box -8 -3 16 105
use FILL  FILL_9645
timestamp 1677677812
transform 1 0 3624 0 1 770
box -8 -3 16 105
use FILL  FILL_9646
timestamp 1677677812
transform 1 0 3632 0 1 770
box -8 -3 16 105
use FILL  FILL_9647
timestamp 1677677812
transform 1 0 3640 0 1 770
box -8 -3 16 105
use FILL  FILL_9648
timestamp 1677677812
transform 1 0 3648 0 1 770
box -8 -3 16 105
use FILL  FILL_9649
timestamp 1677677812
transform 1 0 3656 0 1 770
box -8 -3 16 105
use FILL  FILL_9650
timestamp 1677677812
transform 1 0 3664 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_364
timestamp 1677677812
transform 1 0 3672 0 1 770
box -8 -3 46 105
use FILL  FILL_9652
timestamp 1677677812
transform 1 0 3712 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_38
timestamp 1677677812
transform -1 0 3744 0 1 770
box -8 -3 32 105
use FILL  FILL_9653
timestamp 1677677812
transform 1 0 3744 0 1 770
box -8 -3 16 105
use FILL  FILL_9654
timestamp 1677677812
transform 1 0 3752 0 1 770
box -8 -3 16 105
use FILL  FILL_9655
timestamp 1677677812
transform 1 0 3760 0 1 770
box -8 -3 16 105
use FILL  FILL_9656
timestamp 1677677812
transform 1 0 3768 0 1 770
box -8 -3 16 105
use FILL  FILL_9657
timestamp 1677677812
transform 1 0 3776 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_366
timestamp 1677677812
transform 1 0 3784 0 1 770
box -8 -3 46 105
use FILL  FILL_9667
timestamp 1677677812
transform 1 0 3824 0 1 770
box -8 -3 16 105
use FILL  FILL_9668
timestamp 1677677812
transform 1 0 3832 0 1 770
box -8 -3 16 105
use FILL  FILL_9669
timestamp 1677677812
transform 1 0 3840 0 1 770
box -8 -3 16 105
use FILL  FILL_9670
timestamp 1677677812
transform 1 0 3848 0 1 770
box -8 -3 16 105
use FILL  FILL_9675
timestamp 1677677812
transform 1 0 3856 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_368
timestamp 1677677812
transform 1 0 3864 0 1 770
box -8 -3 46 105
use FILL  FILL_9677
timestamp 1677677812
transform 1 0 3904 0 1 770
box -8 -3 16 105
use FILL  FILL_9684
timestamp 1677677812
transform 1 0 3912 0 1 770
box -8 -3 16 105
use FILL  FILL_9686
timestamp 1677677812
transform 1 0 3920 0 1 770
box -8 -3 16 105
use FILL  FILL_9688
timestamp 1677677812
transform 1 0 3928 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_369
timestamp 1677677812
transform 1 0 3936 0 1 770
box -8 -3 46 105
use FILL  FILL_9690
timestamp 1677677812
transform 1 0 3976 0 1 770
box -8 -3 16 105
use FILL  FILL_9697
timestamp 1677677812
transform 1 0 3984 0 1 770
box -8 -3 16 105
use FILL  FILL_9699
timestamp 1677677812
transform 1 0 3992 0 1 770
box -8 -3 16 105
use FILL  FILL_9701
timestamp 1677677812
transform 1 0 4000 0 1 770
box -8 -3 16 105
use FILL  FILL_9703
timestamp 1677677812
transform 1 0 4008 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_370
timestamp 1677677812
transform -1 0 4056 0 1 770
box -8 -3 46 105
use FILL  FILL_9704
timestamp 1677677812
transform 1 0 4056 0 1 770
box -8 -3 16 105
use FILL  FILL_9712
timestamp 1677677812
transform 1 0 4064 0 1 770
box -8 -3 16 105
use FILL  FILL_9714
timestamp 1677677812
transform 1 0 4072 0 1 770
box -8 -3 16 105
use FILL  FILL_9716
timestamp 1677677812
transform 1 0 4080 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_371
timestamp 1677677812
transform -1 0 4128 0 1 770
box -8 -3 46 105
use FILL  FILL_9717
timestamp 1677677812
transform 1 0 4128 0 1 770
box -8 -3 16 105
use FILL  FILL_9725
timestamp 1677677812
transform 1 0 4136 0 1 770
box -8 -3 16 105
use FILL  FILL_9727
timestamp 1677677812
transform 1 0 4144 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_39
timestamp 1677677812
transform 1 0 4152 0 1 770
box -8 -3 32 105
use FILL  FILL_9729
timestamp 1677677812
transform 1 0 4176 0 1 770
box -8 -3 16 105
use FILL  FILL_9730
timestamp 1677677812
transform 1 0 4184 0 1 770
box -8 -3 16 105
use FILL  FILL_9731
timestamp 1677677812
transform 1 0 4192 0 1 770
box -8 -3 16 105
use FILL  FILL_9732
timestamp 1677677812
transform 1 0 4200 0 1 770
box -8 -3 16 105
use FILL  FILL_9735
timestamp 1677677812
transform 1 0 4208 0 1 770
box -8 -3 16 105
use FILL  FILL_9737
timestamp 1677677812
transform 1 0 4216 0 1 770
box -8 -3 16 105
use FILL  FILL_9739
timestamp 1677677812
transform 1 0 4224 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_373
timestamp 1677677812
transform 1 0 4232 0 1 770
box -8 -3 46 105
use FILL  FILL_9741
timestamp 1677677812
transform 1 0 4272 0 1 770
box -8 -3 16 105
use FILL  FILL_9742
timestamp 1677677812
transform 1 0 4280 0 1 770
box -8 -3 16 105
use FILL  FILL_9743
timestamp 1677677812
transform 1 0 4288 0 1 770
box -8 -3 16 105
use FILL  FILL_9744
timestamp 1677677812
transform 1 0 4296 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_375
timestamp 1677677812
transform 1 0 4304 0 1 770
box -8 -3 46 105
use FILL  FILL_9749
timestamp 1677677812
transform 1 0 4344 0 1 770
box -8 -3 16 105
use FILL  FILL_9750
timestamp 1677677812
transform 1 0 4352 0 1 770
box -8 -3 16 105
use FILL  FILL_9751
timestamp 1677677812
transform 1 0 4360 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_376
timestamp 1677677812
transform 1 0 4368 0 1 770
box -8 -3 46 105
use FILL  FILL_9752
timestamp 1677677812
transform 1 0 4408 0 1 770
box -8 -3 16 105
use FILL  FILL_9753
timestamp 1677677812
transform 1 0 4416 0 1 770
box -8 -3 16 105
use FILL  FILL_9754
timestamp 1677677812
transform 1 0 4424 0 1 770
box -8 -3 16 105
use FILL  FILL_9755
timestamp 1677677812
transform 1 0 4432 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_377
timestamp 1677677812
transform 1 0 4440 0 1 770
box -8 -3 46 105
use FILL  FILL_9756
timestamp 1677677812
transform 1 0 4480 0 1 770
box -8 -3 16 105
use FILL  FILL_9757
timestamp 1677677812
transform 1 0 4488 0 1 770
box -8 -3 16 105
use FILL  FILL_9758
timestamp 1677677812
transform 1 0 4496 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_378
timestamp 1677677812
transform 1 0 4504 0 1 770
box -8 -3 46 105
use FILL  FILL_9759
timestamp 1677677812
transform 1 0 4544 0 1 770
box -8 -3 16 105
use FILL  FILL_9776
timestamp 1677677812
transform 1 0 4552 0 1 770
box -8 -3 16 105
use FILL  FILL_9778
timestamp 1677677812
transform 1 0 4560 0 1 770
box -8 -3 16 105
use FILL  FILL_9780
timestamp 1677677812
transform 1 0 4568 0 1 770
box -8 -3 16 105
use FILL  FILL_9781
timestamp 1677677812
transform 1 0 4576 0 1 770
box -8 -3 16 105
use FILL  FILL_9782
timestamp 1677677812
transform 1 0 4584 0 1 770
box -8 -3 16 105
use FILL  FILL_9783
timestamp 1677677812
transform 1 0 4592 0 1 770
box -8 -3 16 105
use FILL  FILL_9784
timestamp 1677677812
transform 1 0 4600 0 1 770
box -8 -3 16 105
use FILL  FILL_9785
timestamp 1677677812
transform 1 0 4608 0 1 770
box -8 -3 16 105
use FILL  FILL_9787
timestamp 1677677812
transform 1 0 4616 0 1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_383
timestamp 1677677812
transform -1 0 4664 0 1 770
box -8 -3 46 105
use FILL  FILL_9788
timestamp 1677677812
transform 1 0 4664 0 1 770
box -8 -3 16 105
use FILL  FILL_9789
timestamp 1677677812
transform 1 0 4672 0 1 770
box -8 -3 16 105
use FILL  FILL_9790
timestamp 1677677812
transform 1 0 4680 0 1 770
box -8 -3 16 105
use FILL  FILL_9795
timestamp 1677677812
transform 1 0 4688 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_526
timestamp 1677677812
transform 1 0 4696 0 1 770
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_79
timestamp 1677677812
transform 1 0 4819 0 1 770
box -10 -3 10 3
use M2_M1  M2_M1_8439
timestamp 1677677812
transform 1 0 92 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7578
timestamp 1677677812
transform 1 0 172 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8546
timestamp 1677677812
transform 1 0 140 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8547
timestamp 1677677812
transform 1 0 172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8548
timestamp 1677677812
transform 1 0 180 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7624
timestamp 1677677812
transform 1 0 140 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7625
timestamp 1677677812
transform 1 0 180 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8440
timestamp 1677677812
transform 1 0 220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8441
timestamp 1677677812
transform 1 0 228 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8549
timestamp 1677677812
transform 1 0 212 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7706
timestamp 1677677812
transform 1 0 220 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7533
timestamp 1677677812
transform 1 0 252 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7546
timestamp 1677677812
transform 1 0 244 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8442
timestamp 1677677812
transform 1 0 252 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7579
timestamp 1677677812
transform 1 0 260 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8443
timestamp 1677677812
transform 1 0 268 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8550
timestamp 1677677812
transform 1 0 260 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8444
timestamp 1677677812
transform 1 0 300 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7580
timestamp 1677677812
transform 1 0 332 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8551
timestamp 1677677812
transform 1 0 348 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8552
timestamp 1677677812
transform 1 0 380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8553
timestamp 1677677812
transform 1 0 388 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7626
timestamp 1677677812
transform 1 0 348 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7627
timestamp 1677677812
transform 1 0 388 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7676
timestamp 1677677812
transform 1 0 380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7707
timestamp 1677677812
transform 1 0 308 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7547
timestamp 1677677812
transform 1 0 452 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7519
timestamp 1677677812
transform 1 0 476 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8445
timestamp 1677677812
transform 1 0 428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8446
timestamp 1677677812
transform 1 0 436 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8447
timestamp 1677677812
transform 1 0 452 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8448
timestamp 1677677812
transform 1 0 460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8449
timestamp 1677677812
transform 1 0 468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8554
timestamp 1677677812
transform 1 0 428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8555
timestamp 1677677812
transform 1 0 444 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7628
timestamp 1677677812
transform 1 0 444 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7677
timestamp 1677677812
transform 1 0 436 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7629
timestamp 1677677812
transform 1 0 468 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7520
timestamp 1677677812
transform 1 0 532 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7581
timestamp 1677677812
transform 1 0 524 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8556
timestamp 1677677812
transform 1 0 516 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8557
timestamp 1677677812
transform 1 0 524 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7630
timestamp 1677677812
transform 1 0 524 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7548
timestamp 1677677812
transform 1 0 548 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7549
timestamp 1677677812
transform 1 0 588 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8450
timestamp 1677677812
transform 1 0 548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8451
timestamp 1677677812
transform 1 0 572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8558
timestamp 1677677812
transform 1 0 556 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7582
timestamp 1677677812
transform 1 0 580 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8452
timestamp 1677677812
transform 1 0 588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8453
timestamp 1677677812
transform 1 0 604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8559
timestamp 1677677812
transform 1 0 620 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7521
timestamp 1677677812
transform 1 0 636 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8454
timestamp 1677677812
transform 1 0 636 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7583
timestamp 1677677812
transform 1 0 660 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8560
timestamp 1677677812
transform 1 0 660 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8561
timestamp 1677677812
transform 1 0 724 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8562
timestamp 1677677812
transform 1 0 732 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7678
timestamp 1677677812
transform 1 0 676 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8455
timestamp 1677677812
transform 1 0 748 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7522
timestamp 1677677812
transform 1 0 788 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8456
timestamp 1677677812
transform 1 0 764 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8457
timestamp 1677677812
transform 1 0 772 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8458
timestamp 1677677812
transform 1 0 788 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8563
timestamp 1677677812
transform 1 0 796 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8564
timestamp 1677677812
transform 1 0 812 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7631
timestamp 1677677812
transform 1 0 812 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7550
timestamp 1677677812
transform 1 0 828 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8459
timestamp 1677677812
transform 1 0 828 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7551
timestamp 1677677812
transform 1 0 868 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8460
timestamp 1677677812
transform 1 0 844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8461
timestamp 1677677812
transform 1 0 860 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8462
timestamp 1677677812
transform 1 0 884 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8463
timestamp 1677677812
transform 1 0 892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8565
timestamp 1677677812
transform 1 0 836 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7679
timestamp 1677677812
transform 1 0 828 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7604
timestamp 1677677812
transform 1 0 844 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8566
timestamp 1677677812
transform 1 0 852 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8567
timestamp 1677677812
transform 1 0 868 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7605
timestamp 1677677812
transform 1 0 876 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8568
timestamp 1677677812
transform 1 0 884 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7632
timestamp 1677677812
transform 1 0 860 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7680
timestamp 1677677812
transform 1 0 860 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7692
timestamp 1677677812
transform 1 0 836 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7584
timestamp 1677677812
transform 1 0 908 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7585
timestamp 1677677812
transform 1 0 940 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8464
timestamp 1677677812
transform 1 0 988 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8569
timestamp 1677677812
transform 1 0 908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8570
timestamp 1677677812
transform 1 0 940 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7633
timestamp 1677677812
transform 1 0 908 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7534
timestamp 1677677812
transform 1 0 1012 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8434
timestamp 1677677812
transform 1 0 1012 0 1 745
box -2 -2 2 2
use M3_M2  M3_M2_7523
timestamp 1677677812
transform 1 0 1036 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8435
timestamp 1677677812
transform 1 0 1036 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_8465
timestamp 1677677812
transform 1 0 1028 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7552
timestamp 1677677812
transform 1 0 1052 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8571
timestamp 1677677812
transform 1 0 1052 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7634
timestamp 1677677812
transform 1 0 1052 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8466
timestamp 1677677812
transform 1 0 1068 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7635
timestamp 1677677812
transform 1 0 1076 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7535
timestamp 1677677812
transform 1 0 1100 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8572
timestamp 1677677812
transform 1 0 1116 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8573
timestamp 1677677812
transform 1 0 1124 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8574
timestamp 1677677812
transform 1 0 1180 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7606
timestamp 1677677812
transform 1 0 1188 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7693
timestamp 1677677812
transform 1 0 1180 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7524
timestamp 1677677812
transform 1 0 1244 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8467
timestamp 1677677812
transform 1 0 1212 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8468
timestamp 1677677812
transform 1 0 1220 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8469
timestamp 1677677812
transform 1 0 1236 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8470
timestamp 1677677812
transform 1 0 1244 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7607
timestamp 1677677812
transform 1 0 1220 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8575
timestamp 1677677812
transform 1 0 1228 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8576
timestamp 1677677812
transform 1 0 1244 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7525
timestamp 1677677812
transform 1 0 1260 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8577
timestamp 1677677812
transform 1 0 1260 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7536
timestamp 1677677812
transform 1 0 1364 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7537
timestamp 1677677812
transform 1 0 1380 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8471
timestamp 1677677812
transform 1 0 1380 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8578
timestamp 1677677812
transform 1 0 1292 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8579
timestamp 1677677812
transform 1 0 1300 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8580
timestamp 1677677812
transform 1 0 1332 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7636
timestamp 1677677812
transform 1 0 1292 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7637
timestamp 1677677812
transform 1 0 1332 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8581
timestamp 1677677812
transform 1 0 1396 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8472
timestamp 1677677812
transform 1 0 1508 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8582
timestamp 1677677812
transform 1 0 1476 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7694
timestamp 1677677812
transform 1 0 1444 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8473
timestamp 1677677812
transform 1 0 1532 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7538
timestamp 1677677812
transform 1 0 1628 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7539
timestamp 1677677812
transform 1 0 1660 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8474
timestamp 1677677812
transform 1 0 1628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8475
timestamp 1677677812
transform 1 0 1644 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7586
timestamp 1677677812
transform 1 0 1652 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8583
timestamp 1677677812
transform 1 0 1556 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8584
timestamp 1677677812
transform 1 0 1612 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8585
timestamp 1677677812
transform 1 0 1620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8586
timestamp 1677677812
transform 1 0 1636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8587
timestamp 1677677812
transform 1 0 1652 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7638
timestamp 1677677812
transform 1 0 1612 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7639
timestamp 1677677812
transform 1 0 1644 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7695
timestamp 1677677812
transform 1 0 1620 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7553
timestamp 1677677812
transform 1 0 1692 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8476
timestamp 1677677812
transform 1 0 1692 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7587
timestamp 1677677812
transform 1 0 1708 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8588
timestamp 1677677812
transform 1 0 1684 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8589
timestamp 1677677812
transform 1 0 1700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8590
timestamp 1677677812
transform 1 0 1708 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7640
timestamp 1677677812
transform 1 0 1684 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7641
timestamp 1677677812
transform 1 0 1708 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7540
timestamp 1677677812
transform 1 0 1740 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7554
timestamp 1677677812
transform 1 0 1732 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8477
timestamp 1677677812
transform 1 0 1732 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8478
timestamp 1677677812
transform 1 0 1740 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7541
timestamp 1677677812
transform 1 0 1844 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8479
timestamp 1677677812
transform 1 0 1844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8591
timestamp 1677677812
transform 1 0 1756 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8592
timestamp 1677677812
transform 1 0 1764 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8593
timestamp 1677677812
transform 1 0 1820 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7642
timestamp 1677677812
transform 1 0 1756 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7643
timestamp 1677677812
transform 1 0 1772 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7555
timestamp 1677677812
transform 1 0 1860 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7542
timestamp 1677677812
transform 1 0 1876 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7543
timestamp 1677677812
transform 1 0 1892 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8480
timestamp 1677677812
transform 1 0 1884 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7644
timestamp 1677677812
transform 1 0 1884 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7556
timestamp 1677677812
transform 1 0 1900 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8481
timestamp 1677677812
transform 1 0 1900 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8594
timestamp 1677677812
transform 1 0 1908 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8595
timestamp 1677677812
transform 1 0 1916 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7708
timestamp 1677677812
transform 1 0 1916 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8482
timestamp 1677677812
transform 1 0 1948 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8596
timestamp 1677677812
transform 1 0 1940 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8597
timestamp 1677677812
transform 1 0 1956 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7645
timestamp 1677677812
transform 1 0 1940 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7646
timestamp 1677677812
transform 1 0 1964 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7696
timestamp 1677677812
transform 1 0 1956 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7709
timestamp 1677677812
transform 1 0 1964 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8660
timestamp 1677677812
transform 1 0 2060 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8598
timestamp 1677677812
transform 1 0 2076 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8661
timestamp 1677677812
transform 1 0 2076 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7557
timestamp 1677677812
transform 1 0 2100 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7558
timestamp 1677677812
transform 1 0 2172 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8483
timestamp 1677677812
transform 1 0 2172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8599
timestamp 1677677812
transform 1 0 2140 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7608
timestamp 1677677812
transform 1 0 2148 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7647
timestamp 1677677812
transform 1 0 2172 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7559
timestamp 1677677812
transform 1 0 2228 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7560
timestamp 1677677812
transform 1 0 2276 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8484
timestamp 1677677812
transform 1 0 2276 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8600
timestamp 1677677812
transform 1 0 2196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8601
timestamp 1677677812
transform 1 0 2252 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7609
timestamp 1677677812
transform 1 0 2276 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7648
timestamp 1677677812
transform 1 0 2252 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8485
timestamp 1677677812
transform 1 0 2292 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7649
timestamp 1677677812
transform 1 0 2292 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8662
timestamp 1677677812
transform 1 0 2308 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7697
timestamp 1677677812
transform 1 0 2300 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7588
timestamp 1677677812
transform 1 0 2348 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8663
timestamp 1677677812
transform 1 0 2356 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8602
timestamp 1677677812
transform 1 0 2372 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8486
timestamp 1677677812
transform 1 0 2404 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7650
timestamp 1677677812
transform 1 0 2404 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7561
timestamp 1677677812
transform 1 0 2420 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8436
timestamp 1677677812
transform 1 0 2436 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_8487
timestamp 1677677812
transform 1 0 2420 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7589
timestamp 1677677812
transform 1 0 2436 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8603
timestamp 1677677812
transform 1 0 2436 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8488
timestamp 1677677812
transform 1 0 2452 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7562
timestamp 1677677812
transform 1 0 2468 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8489
timestamp 1677677812
transform 1 0 2468 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8604
timestamp 1677677812
transform 1 0 2484 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7651
timestamp 1677677812
transform 1 0 2484 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7563
timestamp 1677677812
transform 1 0 2548 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8490
timestamp 1677677812
transform 1 0 2548 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8491
timestamp 1677677812
transform 1 0 2556 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7590
timestamp 1677677812
transform 1 0 2580 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8492
timestamp 1677677812
transform 1 0 2588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8605
timestamp 1677677812
transform 1 0 2564 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8606
timestamp 1677677812
transform 1 0 2580 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8607
timestamp 1677677812
transform 1 0 2588 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7652
timestamp 1677677812
transform 1 0 2588 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7564
timestamp 1677677812
transform 1 0 2604 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8493
timestamp 1677677812
transform 1 0 2612 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7591
timestamp 1677677812
transform 1 0 2620 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8494
timestamp 1677677812
transform 1 0 2628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8608
timestamp 1677677812
transform 1 0 2620 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8609
timestamp 1677677812
transform 1 0 2636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8610
timestamp 1677677812
transform 1 0 2644 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7698
timestamp 1677677812
transform 1 0 2612 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7699
timestamp 1677677812
transform 1 0 2628 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7592
timestamp 1677677812
transform 1 0 2708 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8495
timestamp 1677677812
transform 1 0 2732 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8611
timestamp 1677677812
transform 1 0 2708 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8612
timestamp 1677677812
transform 1 0 2764 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8613
timestamp 1677677812
transform 1 0 2804 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7653
timestamp 1677677812
transform 1 0 2804 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7593
timestamp 1677677812
transform 1 0 2852 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8496
timestamp 1677677812
transform 1 0 2860 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7610
timestamp 1677677812
transform 1 0 2852 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8497
timestamp 1677677812
transform 1 0 2892 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8614
timestamp 1677677812
transform 1 0 2868 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8615
timestamp 1677677812
transform 1 0 2884 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7654
timestamp 1677677812
transform 1 0 2868 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7700
timestamp 1677677812
transform 1 0 2876 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7611
timestamp 1677677812
transform 1 0 2892 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7612
timestamp 1677677812
transform 1 0 2972 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8616
timestamp 1677677812
transform 1 0 2980 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8664
timestamp 1677677812
transform 1 0 2972 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7681
timestamp 1677677812
transform 1 0 2980 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7565
timestamp 1677677812
transform 1 0 2996 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8498
timestamp 1677677812
transform 1 0 2996 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8499
timestamp 1677677812
transform 1 0 3004 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8617
timestamp 1677677812
transform 1 0 2996 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7655
timestamp 1677677812
transform 1 0 3004 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7613
timestamp 1677677812
transform 1 0 3012 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8665
timestamp 1677677812
transform 1 0 3020 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7682
timestamp 1677677812
transform 1 0 3020 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7526
timestamp 1677677812
transform 1 0 3044 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7544
timestamp 1677677812
transform 1 0 3044 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_7566
timestamp 1677677812
transform 1 0 3036 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8500
timestamp 1677677812
transform 1 0 3044 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8501
timestamp 1677677812
transform 1 0 3068 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8618
timestamp 1677677812
transform 1 0 3044 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8619
timestamp 1677677812
transform 1 0 3060 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8620
timestamp 1677677812
transform 1 0 3100 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7545
timestamp 1677677812
transform 1 0 3124 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_8437
timestamp 1677677812
transform 1 0 3124 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_8438
timestamp 1677677812
transform 1 0 3132 0 1 745
box -2 -2 2 2
use M2_M1  M2_M1_8502
timestamp 1677677812
transform 1 0 3140 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8621
timestamp 1677677812
transform 1 0 3148 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7656
timestamp 1677677812
transform 1 0 3148 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7567
timestamp 1677677812
transform 1 0 3172 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8622
timestamp 1677677812
transform 1 0 3172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8623
timestamp 1677677812
transform 1 0 3196 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8666
timestamp 1677677812
transform 1 0 3180 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_7657
timestamp 1677677812
transform 1 0 3188 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8670
timestamp 1677677812
transform 1 0 3188 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_8624
timestamp 1677677812
transform 1 0 3212 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7527
timestamp 1677677812
transform 1 0 3228 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8667
timestamp 1677677812
transform 1 0 3220 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8668
timestamp 1677677812
transform 1 0 3228 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8503
timestamp 1677677812
transform 1 0 3244 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7658
timestamp 1677677812
transform 1 0 3244 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8504
timestamp 1677677812
transform 1 0 3260 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7528
timestamp 1677677812
transform 1 0 3308 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7529
timestamp 1677677812
transform 1 0 3380 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7568
timestamp 1677677812
transform 1 0 3348 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8505
timestamp 1677677812
transform 1 0 3308 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8506
timestamp 1677677812
transform 1 0 3324 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8625
timestamp 1677677812
transform 1 0 3284 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7614
timestamp 1677677812
transform 1 0 3308 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8626
timestamp 1677677812
transform 1 0 3348 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7659
timestamp 1677677812
transform 1 0 3284 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7701
timestamp 1677677812
transform 1 0 3260 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7530
timestamp 1677677812
transform 1 0 3420 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8627
timestamp 1677677812
transform 1 0 3412 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7660
timestamp 1677677812
transform 1 0 3412 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8507
timestamp 1677677812
transform 1 0 3428 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8508
timestamp 1677677812
transform 1 0 3516 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8628
timestamp 1677677812
transform 1 0 3452 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8629
timestamp 1677677812
transform 1 0 3508 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7661
timestamp 1677677812
transform 1 0 3516 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8669
timestamp 1677677812
transform 1 0 3548 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_8630
timestamp 1677677812
transform 1 0 3580 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7702
timestamp 1677677812
transform 1 0 3580 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8509
timestamp 1677677812
transform 1 0 3588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8631
timestamp 1677677812
transform 1 0 3596 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7683
timestamp 1677677812
transform 1 0 3596 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8510
timestamp 1677677812
transform 1 0 3628 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8511
timestamp 1677677812
transform 1 0 3644 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8632
timestamp 1677677812
transform 1 0 3652 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7662
timestamp 1677677812
transform 1 0 3652 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8512
timestamp 1677677812
transform 1 0 3668 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8633
timestamp 1677677812
transform 1 0 3676 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7684
timestamp 1677677812
transform 1 0 3676 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7710
timestamp 1677677812
transform 1 0 3684 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7594
timestamp 1677677812
transform 1 0 3700 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8513
timestamp 1677677812
transform 1 0 3708 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7569
timestamp 1677677812
transform 1 0 3740 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8514
timestamp 1677677812
transform 1 0 3740 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8515
timestamp 1677677812
transform 1 0 3756 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8634
timestamp 1677677812
transform 1 0 3748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8635
timestamp 1677677812
transform 1 0 3764 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7663
timestamp 1677677812
transform 1 0 3764 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7685
timestamp 1677677812
transform 1 0 3748 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7703
timestamp 1677677812
transform 1 0 3764 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8516
timestamp 1677677812
transform 1 0 3780 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7570
timestamp 1677677812
transform 1 0 3788 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8517
timestamp 1677677812
transform 1 0 3788 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7615
timestamp 1677677812
transform 1 0 3780 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8636
timestamp 1677677812
transform 1 0 3788 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7711
timestamp 1677677812
transform 1 0 3788 0 1 685
box -3 -3 3 3
use M2_M1  M2_M1_8518
timestamp 1677677812
transform 1 0 3828 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7595
timestamp 1677677812
transform 1 0 3836 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8519
timestamp 1677677812
transform 1 0 3844 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8637
timestamp 1677677812
transform 1 0 3820 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8638
timestamp 1677677812
transform 1 0 3836 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7664
timestamp 1677677812
transform 1 0 3812 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7616
timestamp 1677677812
transform 1 0 3844 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7704
timestamp 1677677812
transform 1 0 3828 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_7596
timestamp 1677677812
transform 1 0 3892 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7665
timestamp 1677677812
transform 1 0 3892 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7686
timestamp 1677677812
transform 1 0 3908 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7705
timestamp 1677677812
transform 1 0 3916 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_8639
timestamp 1677677812
transform 1 0 3980 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7712
timestamp 1677677812
transform 1 0 3980 0 1 685
box -3 -3 3 3
use M3_M2  M3_M2_7597
timestamp 1677677812
transform 1 0 4084 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8520
timestamp 1677677812
transform 1 0 4100 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8521
timestamp 1677677812
transform 1 0 4124 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8640
timestamp 1677677812
transform 1 0 4140 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8522
timestamp 1677677812
transform 1 0 4180 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7598
timestamp 1677677812
transform 1 0 4188 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8523
timestamp 1677677812
transform 1 0 4196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8641
timestamp 1677677812
transform 1 0 4172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8642
timestamp 1677677812
transform 1 0 4188 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7617
timestamp 1677677812
transform 1 0 4196 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7666
timestamp 1677677812
transform 1 0 4188 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7687
timestamp 1677677812
transform 1 0 4172 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7599
timestamp 1677677812
transform 1 0 4212 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8643
timestamp 1677677812
transform 1 0 4212 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7600
timestamp 1677677812
transform 1 0 4228 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7531
timestamp 1677677812
transform 1 0 4284 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_7571
timestamp 1677677812
transform 1 0 4260 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8524
timestamp 1677677812
transform 1 0 4260 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7667
timestamp 1677677812
transform 1 0 4252 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7601
timestamp 1677677812
transform 1 0 4268 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7572
timestamp 1677677812
transform 1 0 4300 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8525
timestamp 1677677812
transform 1 0 4276 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8526
timestamp 1677677812
transform 1 0 4292 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8527
timestamp 1677677812
transform 1 0 4300 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8644
timestamp 1677677812
transform 1 0 4284 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7618
timestamp 1677677812
transform 1 0 4292 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8645
timestamp 1677677812
transform 1 0 4300 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7688
timestamp 1677677812
transform 1 0 4300 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7532
timestamp 1677677812
transform 1 0 4332 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_8528
timestamp 1677677812
transform 1 0 4348 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8529
timestamp 1677677812
transform 1 0 4364 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8646
timestamp 1677677812
transform 1 0 4356 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7619
timestamp 1677677812
transform 1 0 4364 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7668
timestamp 1677677812
transform 1 0 4356 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7689
timestamp 1677677812
transform 1 0 4380 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7669
timestamp 1677677812
transform 1 0 4396 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8530
timestamp 1677677812
transform 1 0 4420 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8531
timestamp 1677677812
transform 1 0 4436 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7620
timestamp 1677677812
transform 1 0 4420 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8647
timestamp 1677677812
transform 1 0 4428 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8648
timestamp 1677677812
transform 1 0 4444 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7670
timestamp 1677677812
transform 1 0 4428 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7690
timestamp 1677677812
transform 1 0 4444 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_7573
timestamp 1677677812
transform 1 0 4468 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8532
timestamp 1677677812
transform 1 0 4468 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7574
timestamp 1677677812
transform 1 0 4516 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8533
timestamp 1677677812
transform 1 0 4484 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8534
timestamp 1677677812
transform 1 0 4500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8535
timestamp 1677677812
transform 1 0 4516 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7621
timestamp 1677677812
transform 1 0 4484 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8649
timestamp 1677677812
transform 1 0 4492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8650
timestamp 1677677812
transform 1 0 4508 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8651
timestamp 1677677812
transform 1 0 4524 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7671
timestamp 1677677812
transform 1 0 4532 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7691
timestamp 1677677812
transform 1 0 4524 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_8652
timestamp 1677677812
transform 1 0 4556 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7575
timestamp 1677677812
transform 1 0 4572 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_7576
timestamp 1677677812
transform 1 0 4612 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8536
timestamp 1677677812
transform 1 0 4572 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8537
timestamp 1677677812
transform 1 0 4588 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8538
timestamp 1677677812
transform 1 0 4604 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8539
timestamp 1677677812
transform 1 0 4612 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8653
timestamp 1677677812
transform 1 0 4596 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7622
timestamp 1677677812
transform 1 0 4604 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_7672
timestamp 1677677812
transform 1 0 4580 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7673
timestamp 1677677812
transform 1 0 4596 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_7602
timestamp 1677677812
transform 1 0 4636 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_8654
timestamp 1677677812
transform 1 0 4636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8540
timestamp 1677677812
transform 1 0 4660 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_7603
timestamp 1677677812
transform 1 0 4668 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_7577
timestamp 1677677812
transform 1 0 4684 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_8541
timestamp 1677677812
transform 1 0 4676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8655
timestamp 1677677812
transform 1 0 4652 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8656
timestamp 1677677812
transform 1 0 4668 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7623
timestamp 1677677812
transform 1 0 4676 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_8542
timestamp 1677677812
transform 1 0 4692 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8657
timestamp 1677677812
transform 1 0 4708 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7674
timestamp 1677677812
transform 1 0 4708 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8543
timestamp 1677677812
transform 1 0 4732 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8544
timestamp 1677677812
transform 1 0 4748 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_8658
timestamp 1677677812
transform 1 0 4740 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_8659
timestamp 1677677812
transform 1 0 4756 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_7675
timestamp 1677677812
transform 1 0 4756 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_8545
timestamp 1677677812
transform 1 0 4788 0 1 735
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_80
timestamp 1677677812
transform 1 0 24 0 1 670
box -10 -3 10 3
use FILL  FILL_9362
timestamp 1677677812
transform 1 0 72 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_503
timestamp 1677677812
transform 1 0 80 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_591
timestamp 1677677812
transform -1 0 192 0 -1 770
box -9 -3 26 105
use FILL  FILL_9363
timestamp 1677677812
transform 1 0 192 0 -1 770
box -8 -3 16 105
use FILL  FILL_9365
timestamp 1677677812
transform 1 0 200 0 -1 770
box -8 -3 16 105
use FILL  FILL_9368
timestamp 1677677812
transform 1 0 208 0 -1 770
box -8 -3 16 105
use FILL  FILL_9369
timestamp 1677677812
transform 1 0 216 0 -1 770
box -8 -3 16 105
use FILL  FILL_9370
timestamp 1677677812
transform 1 0 224 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_356
timestamp 1677677812
transform 1 0 232 0 -1 770
box -8 -3 46 105
use FILL  FILL_9371
timestamp 1677677812
transform 1 0 272 0 -1 770
box -8 -3 16 105
use FILL  FILL_9373
timestamp 1677677812
transform 1 0 280 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_505
timestamp 1677677812
transform 1 0 288 0 -1 770
box -8 -3 104 105
use FILL  FILL_9390
timestamp 1677677812
transform 1 0 384 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_595
timestamp 1677677812
transform -1 0 408 0 -1 770
box -9 -3 26 105
use FILL  FILL_9391
timestamp 1677677812
transform 1 0 408 0 -1 770
box -8 -3 16 105
use FILL  FILL_9392
timestamp 1677677812
transform 1 0 416 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_349
timestamp 1677677812
transform -1 0 464 0 -1 770
box -8 -3 46 105
use FILL  FILL_9393
timestamp 1677677812
transform 1 0 464 0 -1 770
box -8 -3 16 105
use FILL  FILL_9394
timestamp 1677677812
transform 1 0 472 0 -1 770
box -8 -3 16 105
use FILL  FILL_9395
timestamp 1677677812
transform 1 0 480 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_596
timestamp 1677677812
transform 1 0 488 0 -1 770
box -9 -3 26 105
use FILL  FILL_9396
timestamp 1677677812
transform 1 0 504 0 -1 770
box -8 -3 16 105
use FILL  FILL_9397
timestamp 1677677812
transform 1 0 512 0 -1 770
box -8 -3 16 105
use FILL  FILL_9398
timestamp 1677677812
transform 1 0 520 0 -1 770
box -8 -3 16 105
use FILL  FILL_9399
timestamp 1677677812
transform 1 0 528 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_350
timestamp 1677677812
transform 1 0 536 0 -1 770
box -8 -3 46 105
use FILL  FILL_9400
timestamp 1677677812
transform 1 0 576 0 -1 770
box -8 -3 16 105
use FILL  FILL_9406
timestamp 1677677812
transform 1 0 584 0 -1 770
box -8 -3 16 105
use FILL  FILL_9407
timestamp 1677677812
transform 1 0 592 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_597
timestamp 1677677812
transform 1 0 600 0 -1 770
box -9 -3 26 105
use FILL  FILL_9408
timestamp 1677677812
transform 1 0 616 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_506
timestamp 1677677812
transform 1 0 624 0 -1 770
box -8 -3 104 105
use FILL  FILL_9409
timestamp 1677677812
transform 1 0 720 0 -1 770
box -8 -3 16 105
use BUFX2  BUFX2_109
timestamp 1677677812
transform 1 0 728 0 -1 770
box -5 -3 28 105
use FILL  FILL_9410
timestamp 1677677812
transform 1 0 752 0 -1 770
box -8 -3 16 105
use FILL  FILL_9411
timestamp 1677677812
transform 1 0 760 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_360
timestamp 1677677812
transform 1 0 768 0 -1 770
box -8 -3 46 105
use FILL  FILL_9419
timestamp 1677677812
transform 1 0 808 0 -1 770
box -8 -3 16 105
use FILL  FILL_9420
timestamp 1677677812
transform 1 0 816 0 -1 770
box -8 -3 16 105
use FILL  FILL_9421
timestamp 1677677812
transform 1 0 824 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_353
timestamp 1677677812
transform 1 0 832 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_599
timestamp 1677677812
transform -1 0 888 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_600
timestamp 1677677812
transform 1 0 888 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_508
timestamp 1677677812
transform -1 0 1000 0 -1 770
box -8 -3 104 105
use FILL  FILL_9422
timestamp 1677677812
transform 1 0 1000 0 -1 770
box -8 -3 16 105
use FILL  FILL_9423
timestamp 1677677812
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_93
timestamp 1677677812
transform 1 0 1016 0 -1 770
box -8 -3 32 105
use FILL  FILL_9426
timestamp 1677677812
transform 1 0 1040 0 -1 770
box -8 -3 16 105
use FILL  FILL_9427
timestamp 1677677812
transform 1 0 1048 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_94
timestamp 1677677812
transform 1 0 1056 0 -1 770
box -8 -3 32 105
use FILL  FILL_9431
timestamp 1677677812
transform 1 0 1080 0 -1 770
box -8 -3 16 105
use FILL  FILL_9432
timestamp 1677677812
transform 1 0 1088 0 -1 770
box -8 -3 16 105
use FILL  FILL_9433
timestamp 1677677812
transform 1 0 1096 0 -1 770
box -8 -3 16 105
use FILL  FILL_9434
timestamp 1677677812
transform 1 0 1104 0 -1 770
box -8 -3 16 105
use FILL  FILL_9435
timestamp 1677677812
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_9436
timestamp 1677677812
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_9437
timestamp 1677677812
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_9438
timestamp 1677677812
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_9439
timestamp 1677677812
transform 1 0 1144 0 -1 770
box -8 -3 16 105
use FILL  FILL_9440
timestamp 1677677812
transform 1 0 1152 0 -1 770
box -8 -3 16 105
use FILL  FILL_9441
timestamp 1677677812
transform 1 0 1160 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_602
timestamp 1677677812
transform -1 0 1184 0 -1 770
box -9 -3 26 105
use FILL  FILL_9442
timestamp 1677677812
transform 1 0 1184 0 -1 770
box -8 -3 16 105
use FILL  FILL_9444
timestamp 1677677812
transform 1 0 1192 0 -1 770
box -8 -3 16 105
use FILL  FILL_9446
timestamp 1677677812
transform 1 0 1200 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_355
timestamp 1677677812
transform 1 0 1208 0 -1 770
box -8 -3 46 105
use FILL  FILL_9448
timestamp 1677677812
transform 1 0 1248 0 -1 770
box -8 -3 16 105
use FILL  FILL_9450
timestamp 1677677812
transform 1 0 1256 0 -1 770
box -8 -3 16 105
use FILL  FILL_9475
timestamp 1677677812
transform 1 0 1264 0 -1 770
box -8 -3 16 105
use FILL  FILL_9476
timestamp 1677677812
transform 1 0 1272 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_606
timestamp 1677677812
transform 1 0 1280 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_513
timestamp 1677677812
transform -1 0 1392 0 -1 770
box -8 -3 104 105
use FILL  FILL_9477
timestamp 1677677812
transform 1 0 1392 0 -1 770
box -8 -3 16 105
use FILL  FILL_9478
timestamp 1677677812
transform 1 0 1400 0 -1 770
box -8 -3 16 105
use FILL  FILL_9479
timestamp 1677677812
transform 1 0 1408 0 -1 770
box -8 -3 16 105
use FILL  FILL_9480
timestamp 1677677812
transform 1 0 1416 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_514
timestamp 1677677812
transform -1 0 1520 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_515
timestamp 1677677812
transform 1 0 1520 0 -1 770
box -8 -3 104 105
use AOI22X1  AOI22X1_359
timestamp 1677677812
transform 1 0 1616 0 -1 770
box -8 -3 46 105
use FILL  FILL_9481
timestamp 1677677812
transform 1 0 1656 0 -1 770
box -8 -3 16 105
use FILL  FILL_9482
timestamp 1677677812
transform 1 0 1664 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_362
timestamp 1677677812
transform -1 0 1712 0 -1 770
box -8 -3 46 105
use FILL  FILL_9483
timestamp 1677677812
transform 1 0 1712 0 -1 770
box -8 -3 16 105
use FILL  FILL_9484
timestamp 1677677812
transform 1 0 1720 0 -1 770
box -8 -3 16 105
use FILL  FILL_9485
timestamp 1677677812
transform 1 0 1728 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_607
timestamp 1677677812
transform 1 0 1736 0 -1 770
box -9 -3 26 105
use FILL  FILL_9486
timestamp 1677677812
transform 1 0 1752 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_516
timestamp 1677677812
transform -1 0 1856 0 -1 770
box -8 -3 104 105
use FILL  FILL_9487
timestamp 1677677812
transform 1 0 1856 0 -1 770
box -8 -3 16 105
use FILL  FILL_9488
timestamp 1677677812
transform 1 0 1864 0 -1 770
box -8 -3 16 105
use FILL  FILL_9489
timestamp 1677677812
transform 1 0 1872 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_608
timestamp 1677677812
transform 1 0 1880 0 -1 770
box -9 -3 26 105
use FILL  FILL_9490
timestamp 1677677812
transform 1 0 1896 0 -1 770
box -8 -3 16 105
use FILL  FILL_9491
timestamp 1677677812
transform 1 0 1904 0 -1 770
box -8 -3 16 105
use FILL  FILL_9492
timestamp 1677677812
transform 1 0 1912 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_360
timestamp 1677677812
transform -1 0 1960 0 -1 770
box -8 -3 46 105
use FILL  FILL_9493
timestamp 1677677812
transform 1 0 1960 0 -1 770
box -8 -3 16 105
use FILL  FILL_9494
timestamp 1677677812
transform 1 0 1968 0 -1 770
box -8 -3 16 105
use FILL  FILL_9496
timestamp 1677677812
transform 1 0 1976 0 -1 770
box -8 -3 16 105
use FILL  FILL_9499
timestamp 1677677812
transform 1 0 1984 0 -1 770
box -8 -3 16 105
use FILL  FILL_9500
timestamp 1677677812
transform 1 0 1992 0 -1 770
box -8 -3 16 105
use FILL  FILL_9501
timestamp 1677677812
transform 1 0 2000 0 -1 770
box -8 -3 16 105
use FILL  FILL_9502
timestamp 1677677812
transform 1 0 2008 0 -1 770
box -8 -3 16 105
use FILL  FILL_9503
timestamp 1677677812
transform 1 0 2016 0 -1 770
box -8 -3 16 105
use FILL  FILL_9504
timestamp 1677677812
transform 1 0 2024 0 -1 770
box -8 -3 16 105
use FILL  FILL_9505
timestamp 1677677812
transform 1 0 2032 0 -1 770
box -8 -3 16 105
use FILL  FILL_9507
timestamp 1677677812
transform 1 0 2040 0 -1 770
box -8 -3 16 105
use FILL  FILL_9509
timestamp 1677677812
transform 1 0 2048 0 -1 770
box -8 -3 16 105
use FILL  FILL_9511
timestamp 1677677812
transform 1 0 2056 0 -1 770
box -8 -3 16 105
use FILL  FILL_9512
timestamp 1677677812
transform 1 0 2064 0 -1 770
box -8 -3 16 105
use FILL  FILL_9513
timestamp 1677677812
transform 1 0 2072 0 -1 770
box -8 -3 16 105
use FILL  FILL_9518
timestamp 1677677812
transform 1 0 2080 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_519
timestamp 1677677812
transform -1 0 2184 0 -1 770
box -8 -3 104 105
use FILL  FILL_9519
timestamp 1677677812
transform 1 0 2184 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_520
timestamp 1677677812
transform -1 0 2288 0 -1 770
box -8 -3 104 105
use FILL  FILL_9520
timestamp 1677677812
transform 1 0 2288 0 -1 770
box -8 -3 16 105
use FILL  FILL_9521
timestamp 1677677812
transform 1 0 2296 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_173
timestamp 1677677812
transform -1 0 2336 0 -1 770
box -8 -3 34 105
use FILL  FILL_9522
timestamp 1677677812
transform 1 0 2336 0 -1 770
box -8 -3 16 105
use FILL  FILL_9524
timestamp 1677677812
transform 1 0 2344 0 -1 770
box -8 -3 16 105
use FILL  FILL_9526
timestamp 1677677812
transform 1 0 2352 0 -1 770
box -8 -3 16 105
use FILL  FILL_9528
timestamp 1677677812
transform 1 0 2360 0 -1 770
box -8 -3 16 105
use FILL  FILL_9530
timestamp 1677677812
transform 1 0 2368 0 -1 770
box -8 -3 16 105
use FILL  FILL_9532
timestamp 1677677812
transform 1 0 2376 0 -1 770
box -8 -3 16 105
use FILL  FILL_9534
timestamp 1677677812
transform 1 0 2384 0 -1 770
box -8 -3 16 105
use FILL  FILL_9536
timestamp 1677677812
transform 1 0 2392 0 -1 770
box -8 -3 16 105
use FILL  FILL_9538
timestamp 1677677812
transform 1 0 2400 0 -1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_16
timestamp 1677677812
transform 1 0 2408 0 -1 770
box -7 -3 39 105
use FILL  FILL_9551
timestamp 1677677812
transform 1 0 2440 0 -1 770
box -8 -3 16 105
use FILL  FILL_9552
timestamp 1677677812
transform 1 0 2448 0 -1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_17
timestamp 1677677812
transform 1 0 2456 0 -1 770
box -7 -3 39 105
use FILL  FILL_9553
timestamp 1677677812
transform 1 0 2488 0 -1 770
box -8 -3 16 105
use FILL  FILL_9554
timestamp 1677677812
transform 1 0 2496 0 -1 770
box -8 -3 16 105
use FILL  FILL_9555
timestamp 1677677812
transform 1 0 2504 0 -1 770
box -8 -3 16 105
use FILL  FILL_9556
timestamp 1677677812
transform 1 0 2512 0 -1 770
box -8 -3 16 105
use FILL  FILL_9557
timestamp 1677677812
transform 1 0 2520 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_611
timestamp 1677677812
transform -1 0 2544 0 -1 770
box -9 -3 26 105
use FILL  FILL_9558
timestamp 1677677812
transform 1 0 2544 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_56
timestamp 1677677812
transform 1 0 2552 0 -1 770
box -8 -3 40 105
use FILL  FILL_9559
timestamp 1677677812
transform 1 0 2584 0 -1 770
box -8 -3 16 105
use FILL  FILL_9560
timestamp 1677677812
transform 1 0 2592 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_363
timestamp 1677677812
transform 1 0 2600 0 -1 770
box -8 -3 46 105
use FILL  FILL_9561
timestamp 1677677812
transform 1 0 2640 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_523
timestamp 1677677812
transform -1 0 2744 0 -1 770
box -8 -3 104 105
use FILL  FILL_9562
timestamp 1677677812
transform 1 0 2744 0 -1 770
box -8 -3 16 105
use FILL  FILL_9563
timestamp 1677677812
transform 1 0 2752 0 -1 770
box -8 -3 16 105
use FILL  FILL_9564
timestamp 1677677812
transform 1 0 2760 0 -1 770
box -8 -3 16 105
use FILL  FILL_9565
timestamp 1677677812
transform 1 0 2768 0 -1 770
box -8 -3 16 105
use FILL  FILL_9566
timestamp 1677677812
transform 1 0 2776 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_57
timestamp 1677677812
transform -1 0 2816 0 -1 770
box -8 -3 40 105
use FILL  FILL_9567
timestamp 1677677812
transform 1 0 2816 0 -1 770
box -8 -3 16 105
use FILL  FILL_9568
timestamp 1677677812
transform 1 0 2824 0 -1 770
box -8 -3 16 105
use FILL  FILL_9569
timestamp 1677677812
transform 1 0 2832 0 -1 770
box -8 -3 16 105
use FILL  FILL_9570
timestamp 1677677812
transform 1 0 2840 0 -1 770
box -8 -3 16 105
use FILL  FILL_9571
timestamp 1677677812
transform 1 0 2848 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_58
timestamp 1677677812
transform 1 0 2856 0 -1 770
box -8 -3 40 105
use FILL  FILL_9580
timestamp 1677677812
transform 1 0 2888 0 -1 770
box -8 -3 16 105
use FILL  FILL_9581
timestamp 1677677812
transform 1 0 2896 0 -1 770
box -8 -3 16 105
use FILL  FILL_9582
timestamp 1677677812
transform 1 0 2904 0 -1 770
box -8 -3 16 105
use FILL  FILL_9583
timestamp 1677677812
transform 1 0 2912 0 -1 770
box -8 -3 16 105
use FILL  FILL_9584
timestamp 1677677812
transform 1 0 2920 0 -1 770
box -8 -3 16 105
use FILL  FILL_9585
timestamp 1677677812
transform 1 0 2928 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1677677812
transform 1 0 2936 0 -1 770
box -8 -3 32 105
use FILL  FILL_9586
timestamp 1677677812
transform 1 0 2960 0 -1 770
box -8 -3 16 105
use FILL  FILL_9587
timestamp 1677677812
transform 1 0 2968 0 -1 770
box -8 -3 16 105
use FILL  FILL_9588
timestamp 1677677812
transform 1 0 2976 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_613
timestamp 1677677812
transform -1 0 3000 0 -1 770
box -9 -3 26 105
use INVX2  INVX2_614
timestamp 1677677812
transform 1 0 3000 0 -1 770
box -9 -3 26 105
use FILL  FILL_9589
timestamp 1677677812
transform 1 0 3016 0 -1 770
box -8 -3 16 105
use FILL  FILL_9590
timestamp 1677677812
transform 1 0 3024 0 -1 770
box -8 -3 16 105
use FILL  FILL_9591
timestamp 1677677812
transform 1 0 3032 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_174
timestamp 1677677812
transform -1 0 3072 0 -1 770
box -8 -3 34 105
use FILL  FILL_9592
timestamp 1677677812
transform 1 0 3072 0 -1 770
box -8 -3 16 105
use FILL  FILL_9594
timestamp 1677677812
transform 1 0 3080 0 -1 770
box -8 -3 16 105
use FILL  FILL_9597
timestamp 1677677812
transform 1 0 3088 0 -1 770
box -8 -3 16 105
use AOI21X1  AOI21X1_18
timestamp 1677677812
transform 1 0 3096 0 -1 770
box -7 -3 39 105
use FILL  FILL_9598
timestamp 1677677812
transform 1 0 3128 0 -1 770
box -8 -3 16 105
use FILL  FILL_9600
timestamp 1677677812
transform 1 0 3136 0 -1 770
box -8 -3 16 105
use FILL  FILL_9602
timestamp 1677677812
transform 1 0 3144 0 -1 770
box -8 -3 16 105
use NOR2X1  NOR2X1_96
timestamp 1677677812
transform 1 0 3152 0 -1 770
box -8 -3 32 105
use NAND3X1  NAND3X1_74
timestamp 1677677812
transform -1 0 3208 0 -1 770
box -8 -3 40 105
use FILL  FILL_9611
timestamp 1677677812
transform 1 0 3208 0 -1 770
box -8 -3 16 105
use FILL  FILL_9612
timestamp 1677677812
transform 1 0 3216 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_35
timestamp 1677677812
transform -1 0 3248 0 -1 770
box -8 -3 32 105
use FILL  FILL_9613
timestamp 1677677812
transform 1 0 3248 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7713
timestamp 1677677812
transform 1 0 3268 0 1 675
box -3 -3 3 3
use XOR2X1  XOR2X1_5
timestamp 1677677812
transform 1 0 3256 0 -1 770
box -8 -3 64 105
use M3_M2  M3_M2_7714
timestamp 1677677812
transform 1 0 3356 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_524
timestamp 1677677812
transform 1 0 3312 0 -1 770
box -8 -3 104 105
use FILL  FILL_9630
timestamp 1677677812
transform 1 0 3408 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_7715
timestamp 1677677812
transform 1 0 3452 0 1 675
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_525
timestamp 1677677812
transform 1 0 3416 0 -1 770
box -8 -3 104 105
use FILL  FILL_9631
timestamp 1677677812
transform 1 0 3512 0 -1 770
box -8 -3 16 105
use FILL  FILL_9632
timestamp 1677677812
transform 1 0 3520 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_37
timestamp 1677677812
transform 1 0 3528 0 -1 770
box -8 -3 32 105
use FILL  FILL_9633
timestamp 1677677812
transform 1 0 3552 0 -1 770
box -8 -3 16 105
use FILL  FILL_9634
timestamp 1677677812
transform 1 0 3560 0 -1 770
box -8 -3 16 105
use FILL  FILL_9636
timestamp 1677677812
transform 1 0 3568 0 -1 770
box -8 -3 16 105
use FILL  FILL_9638
timestamp 1677677812
transform 1 0 3576 0 -1 770
box -8 -3 16 105
use FILL  FILL_9640
timestamp 1677677812
transform 1 0 3584 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_616
timestamp 1677677812
transform 1 0 3592 0 -1 770
box -9 -3 26 105
use FILL  FILL_9643
timestamp 1677677812
transform 1 0 3608 0 -1 770
box -8 -3 16 105
use FILL  FILL_9644
timestamp 1677677812
transform 1 0 3616 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_363
timestamp 1677677812
transform 1 0 3624 0 -1 770
box -8 -3 46 105
use FILL  FILL_9651
timestamp 1677677812
transform 1 0 3664 0 -1 770
box -8 -3 16 105
use FILL  FILL_9658
timestamp 1677677812
transform 1 0 3672 0 -1 770
box -8 -3 16 105
use FILL  FILL_9659
timestamp 1677677812
transform 1 0 3680 0 -1 770
box -8 -3 16 105
use FILL  FILL_9660
timestamp 1677677812
transform 1 0 3688 0 -1 770
box -8 -3 16 105
use FILL  FILL_9661
timestamp 1677677812
transform 1 0 3696 0 -1 770
box -8 -3 16 105
use FILL  FILL_9662
timestamp 1677677812
transform 1 0 3704 0 -1 770
box -8 -3 16 105
use FILL  FILL_9663
timestamp 1677677812
transform 1 0 3712 0 -1 770
box -8 -3 16 105
use FILL  FILL_9664
timestamp 1677677812
transform 1 0 3720 0 -1 770
box -8 -3 16 105
use FILL  FILL_9665
timestamp 1677677812
transform 1 0 3728 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_365
timestamp 1677677812
transform 1 0 3736 0 -1 770
box -8 -3 46 105
use FILL  FILL_9666
timestamp 1677677812
transform 1 0 3776 0 -1 770
box -8 -3 16 105
use FILL  FILL_9671
timestamp 1677677812
transform 1 0 3784 0 -1 770
box -8 -3 16 105
use FILL  FILL_9672
timestamp 1677677812
transform 1 0 3792 0 -1 770
box -8 -3 16 105
use FILL  FILL_9673
timestamp 1677677812
transform 1 0 3800 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_367
timestamp 1677677812
transform 1 0 3808 0 -1 770
box -8 -3 46 105
use FILL  FILL_9674
timestamp 1677677812
transform 1 0 3848 0 -1 770
box -8 -3 16 105
use FILL  FILL_9676
timestamp 1677677812
transform 1 0 3856 0 -1 770
box -8 -3 16 105
use FILL  FILL_9678
timestamp 1677677812
transform 1 0 3864 0 -1 770
box -8 -3 16 105
use FILL  FILL_9679
timestamp 1677677812
transform 1 0 3872 0 -1 770
box -8 -3 16 105
use FILL  FILL_9680
timestamp 1677677812
transform 1 0 3880 0 -1 770
box -8 -3 16 105
use FILL  FILL_9681
timestamp 1677677812
transform 1 0 3888 0 -1 770
box -8 -3 16 105
use FILL  FILL_9682
timestamp 1677677812
transform 1 0 3896 0 -1 770
box -8 -3 16 105
use FILL  FILL_9683
timestamp 1677677812
transform 1 0 3904 0 -1 770
box -8 -3 16 105
use FILL  FILL_9685
timestamp 1677677812
transform 1 0 3912 0 -1 770
box -8 -3 16 105
use FILL  FILL_9687
timestamp 1677677812
transform 1 0 3920 0 -1 770
box -8 -3 16 105
use FILL  FILL_9689
timestamp 1677677812
transform 1 0 3928 0 -1 770
box -8 -3 16 105
use FILL  FILL_9691
timestamp 1677677812
transform 1 0 3936 0 -1 770
box -8 -3 16 105
use FILL  FILL_9692
timestamp 1677677812
transform 1 0 3944 0 -1 770
box -8 -3 16 105
use FILL  FILL_9693
timestamp 1677677812
transform 1 0 3952 0 -1 770
box -8 -3 16 105
use FILL  FILL_9694
timestamp 1677677812
transform 1 0 3960 0 -1 770
box -8 -3 16 105
use FILL  FILL_9695
timestamp 1677677812
transform 1 0 3968 0 -1 770
box -8 -3 16 105
use FILL  FILL_9696
timestamp 1677677812
transform 1 0 3976 0 -1 770
box -8 -3 16 105
use FILL  FILL_9698
timestamp 1677677812
transform 1 0 3984 0 -1 770
box -8 -3 16 105
use FILL  FILL_9700
timestamp 1677677812
transform 1 0 3992 0 -1 770
box -8 -3 16 105
use FILL  FILL_9702
timestamp 1677677812
transform 1 0 4000 0 -1 770
box -8 -3 16 105
use FILL  FILL_9705
timestamp 1677677812
transform 1 0 4008 0 -1 770
box -8 -3 16 105
use FILL  FILL_9706
timestamp 1677677812
transform 1 0 4016 0 -1 770
box -8 -3 16 105
use FILL  FILL_9707
timestamp 1677677812
transform 1 0 4024 0 -1 770
box -8 -3 16 105
use FILL  FILL_9708
timestamp 1677677812
transform 1 0 4032 0 -1 770
box -8 -3 16 105
use FILL  FILL_9709
timestamp 1677677812
transform 1 0 4040 0 -1 770
box -8 -3 16 105
use FILL  FILL_9710
timestamp 1677677812
transform 1 0 4048 0 -1 770
box -8 -3 16 105
use FILL  FILL_9711
timestamp 1677677812
transform 1 0 4056 0 -1 770
box -8 -3 16 105
use FILL  FILL_9713
timestamp 1677677812
transform 1 0 4064 0 -1 770
box -8 -3 16 105
use FILL  FILL_9715
timestamp 1677677812
transform 1 0 4072 0 -1 770
box -8 -3 16 105
use FILL  FILL_9718
timestamp 1677677812
transform 1 0 4080 0 -1 770
box -8 -3 16 105
use FILL  FILL_9719
timestamp 1677677812
transform 1 0 4088 0 -1 770
box -8 -3 16 105
use FILL  FILL_9720
timestamp 1677677812
transform 1 0 4096 0 -1 770
box -8 -3 16 105
use FILL  FILL_9721
timestamp 1677677812
transform 1 0 4104 0 -1 770
box -8 -3 16 105
use FILL  FILL_9722
timestamp 1677677812
transform 1 0 4112 0 -1 770
box -8 -3 16 105
use FILL  FILL_9723
timestamp 1677677812
transform 1 0 4120 0 -1 770
box -8 -3 16 105
use FILL  FILL_9724
timestamp 1677677812
transform 1 0 4128 0 -1 770
box -8 -3 16 105
use FILL  FILL_9726
timestamp 1677677812
transform 1 0 4136 0 -1 770
box -8 -3 16 105
use FILL  FILL_9728
timestamp 1677677812
transform 1 0 4144 0 -1 770
box -8 -3 16 105
use FILL  FILL_9733
timestamp 1677677812
transform 1 0 4152 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_372
timestamp 1677677812
transform 1 0 4160 0 -1 770
box -8 -3 46 105
use FILL  FILL_9734
timestamp 1677677812
transform 1 0 4200 0 -1 770
box -8 -3 16 105
use FILL  FILL_9736
timestamp 1677677812
transform 1 0 4208 0 -1 770
box -8 -3 16 105
use FILL  FILL_9738
timestamp 1677677812
transform 1 0 4216 0 -1 770
box -8 -3 16 105
use FILL  FILL_9740
timestamp 1677677812
transform 1 0 4224 0 -1 770
box -8 -3 16 105
use FILL  FILL_9745
timestamp 1677677812
transform 1 0 4232 0 -1 770
box -8 -3 16 105
use FILL  FILL_9746
timestamp 1677677812
transform 1 0 4240 0 -1 770
box -8 -3 16 105
use FILL  FILL_9747
timestamp 1677677812
transform 1 0 4248 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_374
timestamp 1677677812
transform 1 0 4256 0 -1 770
box -8 -3 46 105
use FILL  FILL_9748
timestamp 1677677812
transform 1 0 4296 0 -1 770
box -8 -3 16 105
use FILL  FILL_9760
timestamp 1677677812
transform 1 0 4304 0 -1 770
box -8 -3 16 105
use FILL  FILL_9761
timestamp 1677677812
transform 1 0 4312 0 -1 770
box -8 -3 16 105
use FILL  FILL_9762
timestamp 1677677812
transform 1 0 4320 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_379
timestamp 1677677812
transform 1 0 4328 0 -1 770
box -8 -3 46 105
use FILL  FILL_9763
timestamp 1677677812
transform 1 0 4368 0 -1 770
box -8 -3 16 105
use FILL  FILL_9764
timestamp 1677677812
transform 1 0 4376 0 -1 770
box -8 -3 16 105
use FILL  FILL_9765
timestamp 1677677812
transform 1 0 4384 0 -1 770
box -8 -3 16 105
use FILL  FILL_9766
timestamp 1677677812
transform 1 0 4392 0 -1 770
box -8 -3 16 105
use FILL  FILL_9767
timestamp 1677677812
transform 1 0 4400 0 -1 770
box -8 -3 16 105
use FILL  FILL_9768
timestamp 1677677812
transform 1 0 4408 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_380
timestamp 1677677812
transform -1 0 4456 0 -1 770
box -8 -3 46 105
use FILL  FILL_9769
timestamp 1677677812
transform 1 0 4456 0 -1 770
box -8 -3 16 105
use FILL  FILL_9770
timestamp 1677677812
transform 1 0 4464 0 -1 770
box -8 -3 16 105
use FILL  FILL_9771
timestamp 1677677812
transform 1 0 4472 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_381
timestamp 1677677812
transform -1 0 4520 0 -1 770
box -8 -3 46 105
use FILL  FILL_9772
timestamp 1677677812
transform 1 0 4520 0 -1 770
box -8 -3 16 105
use FILL  FILL_9773
timestamp 1677677812
transform 1 0 4528 0 -1 770
box -8 -3 16 105
use FILL  FILL_9774
timestamp 1677677812
transform 1 0 4536 0 -1 770
box -8 -3 16 105
use FILL  FILL_9775
timestamp 1677677812
transform 1 0 4544 0 -1 770
box -8 -3 16 105
use FILL  FILL_9777
timestamp 1677677812
transform 1 0 4552 0 -1 770
box -8 -3 16 105
use FILL  FILL_9779
timestamp 1677677812
transform 1 0 4560 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_382
timestamp 1677677812
transform 1 0 4568 0 -1 770
box -8 -3 46 105
use FILL  FILL_9786
timestamp 1677677812
transform 1 0 4608 0 -1 770
box -8 -3 16 105
use FILL  FILL_9791
timestamp 1677677812
transform 1 0 4616 0 -1 770
box -8 -3 16 105
use FILL  FILL_9792
timestamp 1677677812
transform 1 0 4624 0 -1 770
box -8 -3 16 105
use FILL  FILL_9793
timestamp 1677677812
transform 1 0 4632 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_384
timestamp 1677677812
transform 1 0 4640 0 -1 770
box -8 -3 46 105
use FILL  FILL_9794
timestamp 1677677812
transform 1 0 4680 0 -1 770
box -8 -3 16 105
use FILL  FILL_9796
timestamp 1677677812
transform 1 0 4688 0 -1 770
box -8 -3 16 105
use FILL  FILL_9797
timestamp 1677677812
transform 1 0 4696 0 -1 770
box -8 -3 16 105
use FILL  FILL_9798
timestamp 1677677812
transform 1 0 4704 0 -1 770
box -8 -3 16 105
use OAI22X1  OAI22X1_385
timestamp 1677677812
transform 1 0 4712 0 -1 770
box -8 -3 46 105
use FILL  FILL_9799
timestamp 1677677812
transform 1 0 4752 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_617
timestamp 1677677812
transform -1 0 4776 0 -1 770
box -9 -3 26 105
use FILL  FILL_9800
timestamp 1677677812
transform 1 0 4776 0 -1 770
box -8 -3 16 105
use FILL  FILL_9801
timestamp 1677677812
transform 1 0 4784 0 -1 770
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_81
timestamp 1677677812
transform 1 0 4843 0 1 670
box -10 -3 10 3
use M2_M1  M2_M1_8676
timestamp 1677677812
transform 1 0 108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8677
timestamp 1677677812
transform 1 0 164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8678
timestamp 1677677812
transform 1 0 172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8791
timestamp 1677677812
transform 1 0 84 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7828
timestamp 1677677812
transform 1 0 164 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7753
timestamp 1677677812
transform 1 0 204 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7790
timestamp 1677677812
transform 1 0 196 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7733
timestamp 1677677812
transform 1 0 236 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7754
timestamp 1677677812
transform 1 0 236 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8679
timestamp 1677677812
transform 1 0 204 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8680
timestamp 1677677812
transform 1 0 220 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8681
timestamp 1677677812
transform 1 0 236 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8792
timestamp 1677677812
transform 1 0 188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8793
timestamp 1677677812
transform 1 0 204 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7829
timestamp 1677677812
transform 1 0 204 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7817
timestamp 1677677812
transform 1 0 236 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8794
timestamp 1677677812
transform 1 0 244 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8795
timestamp 1677677812
transform 1 0 268 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7755
timestamp 1677677812
transform 1 0 292 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8682
timestamp 1677677812
transform 1 0 292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8683
timestamp 1677677812
transform 1 0 308 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7791
timestamp 1677677812
transform 1 0 316 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8684
timestamp 1677677812
transform 1 0 324 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8685
timestamp 1677677812
transform 1 0 332 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8796
timestamp 1677677812
transform 1 0 316 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8797
timestamp 1677677812
transform 1 0 340 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7792
timestamp 1677677812
transform 1 0 348 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7830
timestamp 1677677812
transform 1 0 340 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7756
timestamp 1677677812
transform 1 0 364 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8686
timestamp 1677677812
transform 1 0 364 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7734
timestamp 1677677812
transform 1 0 428 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7757
timestamp 1677677812
transform 1 0 420 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7793
timestamp 1677677812
transform 1 0 396 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7758
timestamp 1677677812
transform 1 0 460 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8687
timestamp 1677677812
transform 1 0 404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8688
timestamp 1677677812
transform 1 0 420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8689
timestamp 1677677812
transform 1 0 428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8690
timestamp 1677677812
transform 1 0 444 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8691
timestamp 1677677812
transform 1 0 460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8798
timestamp 1677677812
transform 1 0 388 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8799
timestamp 1677677812
transform 1 0 396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8800
timestamp 1677677812
transform 1 0 412 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7831
timestamp 1677677812
transform 1 0 412 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8801
timestamp 1677677812
transform 1 0 436 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8802
timestamp 1677677812
transform 1 0 452 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7832
timestamp 1677677812
transform 1 0 436 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8692
timestamp 1677677812
transform 1 0 516 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8693
timestamp 1677677812
transform 1 0 572 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8694
timestamp 1677677812
transform 1 0 580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8803
timestamp 1677677812
transform 1 0 492 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7818
timestamp 1677677812
transform 1 0 580 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7833
timestamp 1677677812
transform 1 0 524 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7834
timestamp 1677677812
transform 1 0 572 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7863
timestamp 1677677812
transform 1 0 540 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8695
timestamp 1677677812
transform 1 0 620 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7794
timestamp 1677677812
transform 1 0 628 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8696
timestamp 1677677812
transform 1 0 636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8804
timestamp 1677677812
transform 1 0 604 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8805
timestamp 1677677812
transform 1 0 628 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8806
timestamp 1677677812
transform 1 0 636 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7835
timestamp 1677677812
transform 1 0 604 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7759
timestamp 1677677812
transform 1 0 660 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7836
timestamp 1677677812
transform 1 0 652 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7760
timestamp 1677677812
transform 1 0 676 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8697
timestamp 1677677812
transform 1 0 676 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7761
timestamp 1677677812
transform 1 0 716 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8698
timestamp 1677677812
transform 1 0 716 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7795
timestamp 1677677812
transform 1 0 764 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8699
timestamp 1677677812
transform 1 0 772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8807
timestamp 1677677812
transform 1 0 692 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7864
timestamp 1677677812
transform 1 0 692 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8700
timestamp 1677677812
transform 1 0 788 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7819
timestamp 1677677812
transform 1 0 788 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8808
timestamp 1677677812
transform 1 0 820 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7735
timestamp 1677677812
transform 1 0 852 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8701
timestamp 1677677812
transform 1 0 836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8702
timestamp 1677677812
transform 1 0 852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8703
timestamp 1677677812
transform 1 0 868 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8809
timestamp 1677677812
transform 1 0 844 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8810
timestamp 1677677812
transform 1 0 860 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7736
timestamp 1677677812
transform 1 0 892 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7762
timestamp 1677677812
transform 1 0 884 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7763
timestamp 1677677812
transform 1 0 956 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8704
timestamp 1677677812
transform 1 0 956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8811
timestamp 1677677812
transform 1 0 1004 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8896
timestamp 1677677812
transform 1 0 1020 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7865
timestamp 1677677812
transform 1 0 964 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7866
timestamp 1677677812
transform 1 0 1012 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7716
timestamp 1677677812
transform 1 0 1060 0 1 655
box -3 -3 3 3
use M3_M2  M3_M2_7764
timestamp 1677677812
transform 1 0 1156 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8705
timestamp 1677677812
transform 1 0 1060 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7796
timestamp 1677677812
transform 1 0 1076 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7797
timestamp 1677677812
transform 1 0 1100 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7718
timestamp 1677677812
transform 1 0 1188 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8706
timestamp 1677677812
transform 1 0 1124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8707
timestamp 1677677812
transform 1 0 1156 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8708
timestamp 1677677812
transform 1 0 1164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8709
timestamp 1677677812
transform 1 0 1172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8710
timestamp 1677677812
transform 1 0 1196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8812
timestamp 1677677812
transform 1 0 1052 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7820
timestamp 1677677812
transform 1 0 1060 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8813
timestamp 1677677812
transform 1 0 1076 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7837
timestamp 1677677812
transform 1 0 1116 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7798
timestamp 1677677812
transform 1 0 1204 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8814
timestamp 1677677812
transform 1 0 1180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8815
timestamp 1677677812
transform 1 0 1188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8816
timestamp 1677677812
transform 1 0 1204 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7867
timestamp 1677677812
transform 1 0 1060 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7868
timestamp 1677677812
transform 1 0 1148 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7869
timestamp 1677677812
transform 1 0 1172 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8711
timestamp 1677677812
transform 1 0 1220 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7719
timestamp 1677677812
transform 1 0 1228 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7737
timestamp 1677677812
transform 1 0 1236 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7799
timestamp 1677677812
transform 1 0 1236 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8712
timestamp 1677677812
transform 1 0 1244 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7765
timestamp 1677677812
transform 1 0 1260 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8817
timestamp 1677677812
transform 1 0 1260 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7720
timestamp 1677677812
transform 1 0 1268 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8713
timestamp 1677677812
transform 1 0 1268 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7717
timestamp 1677677812
transform 1 0 1300 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_8714
timestamp 1677677812
transform 1 0 1292 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8715
timestamp 1677677812
transform 1 0 1308 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8818
timestamp 1677677812
transform 1 0 1300 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7721
timestamp 1677677812
transform 1 0 1380 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7766
timestamp 1677677812
transform 1 0 1356 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7800
timestamp 1677677812
transform 1 0 1348 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7722
timestamp 1677677812
transform 1 0 1412 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7767
timestamp 1677677812
transform 1 0 1404 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8716
timestamp 1677677812
transform 1 0 1356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8717
timestamp 1677677812
transform 1 0 1372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8718
timestamp 1677677812
transform 1 0 1388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8819
timestamp 1677677812
transform 1 0 1348 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7838
timestamp 1677677812
transform 1 0 1348 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8820
timestamp 1677677812
transform 1 0 1364 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8821
timestamp 1677677812
transform 1 0 1380 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7839
timestamp 1677677812
transform 1 0 1372 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7801
timestamp 1677677812
transform 1 0 1396 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8719
timestamp 1677677812
transform 1 0 1404 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8822
timestamp 1677677812
transform 1 0 1396 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7738
timestamp 1677677812
transform 1 0 1420 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8720
timestamp 1677677812
transform 1 0 1436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8721
timestamp 1677677812
transform 1 0 1460 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8823
timestamp 1677677812
transform 1 0 1444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8824
timestamp 1677677812
transform 1 0 1452 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7870
timestamp 1677677812
transform 1 0 1420 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7871
timestamp 1677677812
transform 1 0 1452 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8722
timestamp 1677677812
transform 1 0 1476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8825
timestamp 1677677812
transform 1 0 1476 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7872
timestamp 1677677812
transform 1 0 1476 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7873
timestamp 1677677812
transform 1 0 1508 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8723
timestamp 1677677812
transform 1 0 1524 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8724
timestamp 1677677812
transform 1 0 1556 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7874
timestamp 1677677812
transform 1 0 1556 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7802
timestamp 1677677812
transform 1 0 1564 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8826
timestamp 1677677812
transform 1 0 1564 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8827
timestamp 1677677812
transform 1 0 1572 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7840
timestamp 1677677812
transform 1 0 1572 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7768
timestamp 1677677812
transform 1 0 1580 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7769
timestamp 1677677812
transform 1 0 1620 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8725
timestamp 1677677812
transform 1 0 1580 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8726
timestamp 1677677812
transform 1 0 1588 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8727
timestamp 1677677812
transform 1 0 1620 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7803
timestamp 1677677812
transform 1 0 1636 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7723
timestamp 1677677812
transform 1 0 1724 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7770
timestamp 1677677812
transform 1 0 1692 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7771
timestamp 1677677812
transform 1 0 1716 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8728
timestamp 1677677812
transform 1 0 1692 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8729
timestamp 1677677812
transform 1 0 1708 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8828
timestamp 1677677812
transform 1 0 1668 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8829
timestamp 1677677812
transform 1 0 1684 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7875
timestamp 1677677812
transform 1 0 1668 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7821
timestamp 1677677812
transform 1 0 1692 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8830
timestamp 1677677812
transform 1 0 1700 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8730
timestamp 1677677812
transform 1 0 1724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8831
timestamp 1677677812
transform 1 0 1732 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7841
timestamp 1677677812
transform 1 0 1732 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7772
timestamp 1677677812
transform 1 0 1756 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7804
timestamp 1677677812
transform 1 0 1748 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7739
timestamp 1677677812
transform 1 0 1812 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7773
timestamp 1677677812
transform 1 0 1820 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8731
timestamp 1677677812
transform 1 0 1756 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8732
timestamp 1677677812
transform 1 0 1772 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8733
timestamp 1677677812
transform 1 0 1796 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7805
timestamp 1677677812
transform 1 0 1804 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8734
timestamp 1677677812
transform 1 0 1812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8735
timestamp 1677677812
transform 1 0 1828 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8832
timestamp 1677677812
transform 1 0 1748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8833
timestamp 1677677812
transform 1 0 1764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8834
timestamp 1677677812
transform 1 0 1772 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8835
timestamp 1677677812
transform 1 0 1804 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8836
timestamp 1677677812
transform 1 0 1820 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7842
timestamp 1677677812
transform 1 0 1764 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8736
timestamp 1677677812
transform 1 0 1860 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8737
timestamp 1677677812
transform 1 0 1908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8738
timestamp 1677677812
transform 1 0 1964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8739
timestamp 1677677812
transform 1 0 1972 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8740
timestamp 1677677812
transform 1 0 2028 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8837
timestamp 1677677812
transform 1 0 1940 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8838
timestamp 1677677812
transform 1 0 1956 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7806
timestamp 1677677812
transform 1 0 2052 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8839
timestamp 1677677812
transform 1 0 2052 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7843
timestamp 1677677812
transform 1 0 2036 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7844
timestamp 1677677812
transform 1 0 2052 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7845
timestamp 1677677812
transform 1 0 2076 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8741
timestamp 1677677812
transform 1 0 2116 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8742
timestamp 1677677812
transform 1 0 2172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8840
timestamp 1677677812
transform 1 0 2092 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7774
timestamp 1677677812
transform 1 0 2268 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8743
timestamp 1677677812
transform 1 0 2268 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8841
timestamp 1677677812
transform 1 0 2220 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7876
timestamp 1677677812
transform 1 0 2220 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7775
timestamp 1677677812
transform 1 0 2308 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8744
timestamp 1677677812
transform 1 0 2316 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8842
timestamp 1677677812
transform 1 0 2308 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8672
timestamp 1677677812
transform 1 0 2340 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8745
timestamp 1677677812
transform 1 0 2372 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8746
timestamp 1677677812
transform 1 0 2396 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8747
timestamp 1677677812
transform 1 0 2436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8843
timestamp 1677677812
transform 1 0 2412 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8844
timestamp 1677677812
transform 1 0 2420 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7846
timestamp 1677677812
transform 1 0 2420 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7847
timestamp 1677677812
transform 1 0 2468 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7724
timestamp 1677677812
transform 1 0 2532 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7725
timestamp 1677677812
transform 1 0 2556 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7776
timestamp 1677677812
transform 1 0 2524 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7807
timestamp 1677677812
transform 1 0 2516 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8845
timestamp 1677677812
transform 1 0 2516 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7777
timestamp 1677677812
transform 1 0 2548 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8748
timestamp 1677677812
transform 1 0 2540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8749
timestamp 1677677812
transform 1 0 2548 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8846
timestamp 1677677812
transform 1 0 2532 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7778
timestamp 1677677812
transform 1 0 2564 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8847
timestamp 1677677812
transform 1 0 2556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8897
timestamp 1677677812
transform 1 0 2524 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7848
timestamp 1677677812
transform 1 0 2532 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7808
timestamp 1677677812
transform 1 0 2620 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8750
timestamp 1677677812
transform 1 0 2628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8751
timestamp 1677677812
transform 1 0 2644 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7726
timestamp 1677677812
transform 1 0 2660 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8848
timestamp 1677677812
transform 1 0 2660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7740
timestamp 1677677812
transform 1 0 2740 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8752
timestamp 1677677812
transform 1 0 2740 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8849
timestamp 1677677812
transform 1 0 2764 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8850
timestamp 1677677812
transform 1 0 2804 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7741
timestamp 1677677812
transform 1 0 2868 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8753
timestamp 1677677812
transform 1 0 2852 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8851
timestamp 1677677812
transform 1 0 2876 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8754
timestamp 1677677812
transform 1 0 2900 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8852
timestamp 1677677812
transform 1 0 2924 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8673
timestamp 1677677812
transform 1 0 2972 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8674
timestamp 1677677812
transform 1 0 2996 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_8755
timestamp 1677677812
transform 1 0 2988 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8756
timestamp 1677677812
transform 1 0 3004 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8671
timestamp 1677677812
transform 1 0 3012 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_7809
timestamp 1677677812
transform 1 0 3012 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7727
timestamp 1677677812
transform 1 0 3044 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8853
timestamp 1677677812
transform 1 0 3044 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8898
timestamp 1677677812
transform 1 0 3084 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7742
timestamp 1677677812
transform 1 0 3100 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8757
timestamp 1677677812
transform 1 0 3100 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7728
timestamp 1677677812
transform 1 0 3132 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7779
timestamp 1677677812
transform 1 0 3140 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8758
timestamp 1677677812
transform 1 0 3124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8759
timestamp 1677677812
transform 1 0 3140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8854
timestamp 1677677812
transform 1 0 3116 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7877
timestamp 1677677812
transform 1 0 3116 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8855
timestamp 1677677812
transform 1 0 3148 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7849
timestamp 1677677812
transform 1 0 3132 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7878
timestamp 1677677812
transform 1 0 3140 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8760
timestamp 1677677812
transform 1 0 3164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8856
timestamp 1677677812
transform 1 0 3164 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7850
timestamp 1677677812
transform 1 0 3164 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7743
timestamp 1677677812
transform 1 0 3180 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7810
timestamp 1677677812
transform 1 0 3180 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8857
timestamp 1677677812
transform 1 0 3180 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8899
timestamp 1677677812
transform 1 0 3180 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_8900
timestamp 1677677812
transform 1 0 3236 0 1 595
box -2 -2 2 2
use M2_M1  M2_M1_8901
timestamp 1677677812
transform 1 0 3260 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7744
timestamp 1677677812
transform 1 0 3276 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7780
timestamp 1677677812
transform 1 0 3284 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8761
timestamp 1677677812
transform 1 0 3276 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8858
timestamp 1677677812
transform 1 0 3284 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8902
timestamp 1677677812
transform 1 0 3276 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_7745
timestamp 1677677812
transform 1 0 3300 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8762
timestamp 1677677812
transform 1 0 3300 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7729
timestamp 1677677812
transform 1 0 3356 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7746
timestamp 1677677812
transform 1 0 3396 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7747
timestamp 1677677812
transform 1 0 3452 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8763
timestamp 1677677812
transform 1 0 3356 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8764
timestamp 1677677812
transform 1 0 3412 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8765
timestamp 1677677812
transform 1 0 3452 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7811
timestamp 1677677812
transform 1 0 3500 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8859
timestamp 1677677812
transform 1 0 3332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7822
timestamp 1677677812
transform 1 0 3412 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8860
timestamp 1677677812
transform 1 0 3428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8675
timestamp 1677677812
transform 1 0 3548 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_7823
timestamp 1677677812
transform 1 0 3564 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8766
timestamp 1677677812
transform 1 0 3580 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7824
timestamp 1677677812
transform 1 0 3580 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7781
timestamp 1677677812
transform 1 0 3612 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8767
timestamp 1677677812
transform 1 0 3596 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8768
timestamp 1677677812
transform 1 0 3612 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8861
timestamp 1677677812
transform 1 0 3588 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8862
timestamp 1677677812
transform 1 0 3604 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7879
timestamp 1677677812
transform 1 0 3588 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7880
timestamp 1677677812
transform 1 0 3604 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8863
timestamp 1677677812
transform 1 0 3636 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7851
timestamp 1677677812
transform 1 0 3636 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7782
timestamp 1677677812
transform 1 0 3652 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8864
timestamp 1677677812
transform 1 0 3652 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8865
timestamp 1677677812
transform 1 0 3660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7881
timestamp 1677677812
transform 1 0 3660 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8769
timestamp 1677677812
transform 1 0 3684 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8770
timestamp 1677677812
transform 1 0 3700 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8866
timestamp 1677677812
transform 1 0 3692 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8867
timestamp 1677677812
transform 1 0 3708 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7852
timestamp 1677677812
transform 1 0 3708 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8771
timestamp 1677677812
transform 1 0 3780 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7825
timestamp 1677677812
transform 1 0 3828 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8868
timestamp 1677677812
transform 1 0 3836 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7748
timestamp 1677677812
transform 1 0 3908 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7783
timestamp 1677677812
transform 1 0 3892 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8772
timestamp 1677677812
transform 1 0 3892 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8773
timestamp 1677677812
transform 1 0 3908 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8869
timestamp 1677677812
transform 1 0 3884 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8870
timestamp 1677677812
transform 1 0 3900 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8871
timestamp 1677677812
transform 1 0 3916 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8872
timestamp 1677677812
transform 1 0 3924 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7853
timestamp 1677677812
transform 1 0 3884 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7854
timestamp 1677677812
transform 1 0 3924 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7882
timestamp 1677677812
transform 1 0 3916 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7883
timestamp 1677677812
transform 1 0 3940 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7730
timestamp 1677677812
transform 1 0 3964 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_8774
timestamp 1677677812
transform 1 0 3964 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8775
timestamp 1677677812
transform 1 0 3980 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8873
timestamp 1677677812
transform 1 0 3972 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8874
timestamp 1677677812
transform 1 0 3988 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7884
timestamp 1677677812
transform 1 0 3988 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7812
timestamp 1677677812
transform 1 0 4012 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7784
timestamp 1677677812
transform 1 0 4028 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7813
timestamp 1677677812
transform 1 0 4028 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7749
timestamp 1677677812
transform 1 0 4060 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7785
timestamp 1677677812
transform 1 0 4044 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8776
timestamp 1677677812
transform 1 0 4044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8777
timestamp 1677677812
transform 1 0 4060 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8875
timestamp 1677677812
transform 1 0 4036 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8876
timestamp 1677677812
transform 1 0 4052 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7885
timestamp 1677677812
transform 1 0 4036 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7731
timestamp 1677677812
transform 1 0 4124 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7750
timestamp 1677677812
transform 1 0 4116 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7751
timestamp 1677677812
transform 1 0 4148 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_8778
timestamp 1677677812
transform 1 0 4124 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8779
timestamp 1677677812
transform 1 0 4140 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8780
timestamp 1677677812
transform 1 0 4148 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8877
timestamp 1677677812
transform 1 0 4108 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8878
timestamp 1677677812
transform 1 0 4116 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8879
timestamp 1677677812
transform 1 0 4132 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8880
timestamp 1677677812
transform 1 0 4148 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7855
timestamp 1677677812
transform 1 0 4108 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7886
timestamp 1677677812
transform 1 0 4116 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7856
timestamp 1677677812
transform 1 0 4148 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7732
timestamp 1677677812
transform 1 0 4188 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_7752
timestamp 1677677812
transform 1 0 4212 0 1 635
box -3 -3 3 3
use M3_M2  M3_M2_7786
timestamp 1677677812
transform 1 0 4212 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8781
timestamp 1677677812
transform 1 0 4212 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8881
timestamp 1677677812
transform 1 0 4188 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8882
timestamp 1677677812
transform 1 0 4204 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7857
timestamp 1677677812
transform 1 0 4188 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8883
timestamp 1677677812
transform 1 0 4228 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7858
timestamp 1677677812
transform 1 0 4236 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7787
timestamp 1677677812
transform 1 0 4284 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8782
timestamp 1677677812
transform 1 0 4340 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7859
timestamp 1677677812
transform 1 0 4340 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8884
timestamp 1677677812
transform 1 0 4396 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8783
timestamp 1677677812
transform 1 0 4476 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7788
timestamp 1677677812
transform 1 0 4540 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_8784
timestamp 1677677812
transform 1 0 4540 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8785
timestamp 1677677812
transform 1 0 4556 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8786
timestamp 1677677812
transform 1 0 4580 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7814
timestamp 1677677812
transform 1 0 4588 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8885
timestamp 1677677812
transform 1 0 4508 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8886
timestamp 1677677812
transform 1 0 4516 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8887
timestamp 1677677812
transform 1 0 4532 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8888
timestamp 1677677812
transform 1 0 4548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8889
timestamp 1677677812
transform 1 0 4556 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8890
timestamp 1677677812
transform 1 0 4572 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8891
timestamp 1677677812
transform 1 0 4588 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8892
timestamp 1677677812
transform 1 0 4596 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7860
timestamp 1677677812
transform 1 0 4556 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7789
timestamp 1677677812
transform 1 0 4604 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_7861
timestamp 1677677812
transform 1 0 4596 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_8787
timestamp 1677677812
transform 1 0 4636 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8788
timestamp 1677677812
transform 1 0 4652 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7815
timestamp 1677677812
transform 1 0 4660 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_8789
timestamp 1677677812
transform 1 0 4668 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_8893
timestamp 1677677812
transform 1 0 4644 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_8894
timestamp 1677677812
transform 1 0 4660 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_7887
timestamp 1677677812
transform 1 0 4652 0 1 585
box -3 -3 3 3
use M2_M1  M2_M1_8790
timestamp 1677677812
transform 1 0 4684 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_7826
timestamp 1677677812
transform 1 0 4684 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_7888
timestamp 1677677812
transform 1 0 4692 0 1 585
box -3 -3 3 3
use M3_M2  M3_M2_7862
timestamp 1677677812
transform 1 0 4708 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_7816
timestamp 1677677812
transform 1 0 4740 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_7827
timestamp 1677677812
transform 1 0 4748 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_8895
timestamp 1677677812
transform 1 0 4788 0 1 605
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_82
timestamp 1677677812
transform 1 0 48 0 1 570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_527
timestamp 1677677812
transform 1 0 72 0 1 570
box -8 -3 104 105
use INVX2  INVX2_618
timestamp 1677677812
transform -1 0 184 0 1 570
box -9 -3 26 105
use FILL  FILL_9802
timestamp 1677677812
transform 1 0 184 0 1 570
box -8 -3 16 105
use FILL  FILL_9803
timestamp 1677677812
transform 1 0 192 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7889
timestamp 1677677812
transform 1 0 236 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_366
timestamp 1677677812
transform -1 0 240 0 1 570
box -8 -3 46 105
use FILL  FILL_9804
timestamp 1677677812
transform 1 0 240 0 1 570
box -8 -3 16 105
use FILL  FILL_9805
timestamp 1677677812
transform 1 0 248 0 1 570
box -8 -3 16 105
use FILL  FILL_9806
timestamp 1677677812
transform 1 0 256 0 1 570
box -8 -3 16 105
use FILL  FILL_9807
timestamp 1677677812
transform 1 0 264 0 1 570
box -8 -3 16 105
use FILL  FILL_9808
timestamp 1677677812
transform 1 0 272 0 1 570
box -8 -3 16 105
use FILL  FILL_9809
timestamp 1677677812
transform 1 0 280 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_367
timestamp 1677677812
transform -1 0 328 0 1 570
box -8 -3 46 105
use FILL  FILL_9810
timestamp 1677677812
transform 1 0 328 0 1 570
box -8 -3 16 105
use FILL  FILL_9811
timestamp 1677677812
transform 1 0 336 0 1 570
box -8 -3 16 105
use FILL  FILL_9812
timestamp 1677677812
transform 1 0 344 0 1 570
box -8 -3 16 105
use INVX2  INVX2_619
timestamp 1677677812
transform -1 0 368 0 1 570
box -9 -3 26 105
use FILL  FILL_9813
timestamp 1677677812
transform 1 0 368 0 1 570
box -8 -3 16 105
use FILL  FILL_9826
timestamp 1677677812
transform 1 0 376 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_369
timestamp 1677677812
transform -1 0 424 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_370
timestamp 1677677812
transform -1 0 464 0 1 570
box -8 -3 46 105
use FILL  FILL_9828
timestamp 1677677812
transform 1 0 464 0 1 570
box -8 -3 16 105
use FILL  FILL_9829
timestamp 1677677812
transform 1 0 472 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_529
timestamp 1677677812
transform 1 0 480 0 1 570
box -8 -3 104 105
use FILL  FILL_9830
timestamp 1677677812
transform 1 0 576 0 1 570
box -8 -3 16 105
use FILL  FILL_9831
timestamp 1677677812
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_9832
timestamp 1677677812
transform 1 0 592 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_371
timestamp 1677677812
transform 1 0 600 0 1 570
box -8 -3 46 105
use FILL  FILL_9833
timestamp 1677677812
transform 1 0 640 0 1 570
box -8 -3 16 105
use FILL  FILL_9834
timestamp 1677677812
transform 1 0 648 0 1 570
box -8 -3 16 105
use INVX2  INVX2_622
timestamp 1677677812
transform 1 0 656 0 1 570
box -9 -3 26 105
use FILL  FILL_9835
timestamp 1677677812
transform 1 0 672 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_530
timestamp 1677677812
transform 1 0 680 0 1 570
box -8 -3 104 105
use FILL  FILL_9836
timestamp 1677677812
transform 1 0 776 0 1 570
box -8 -3 16 105
use FILL  FILL_9837
timestamp 1677677812
transform 1 0 784 0 1 570
box -8 -3 16 105
use FILL  FILL_9838
timestamp 1677677812
transform 1 0 792 0 1 570
box -8 -3 16 105
use FILL  FILL_9849
timestamp 1677677812
transform 1 0 800 0 1 570
box -8 -3 16 105
use FILL  FILL_9851
timestamp 1677677812
transform 1 0 808 0 1 570
box -8 -3 16 105
use FILL  FILL_9852
timestamp 1677677812
transform 1 0 816 0 1 570
box -8 -3 16 105
use FILL  FILL_9853
timestamp 1677677812
transform 1 0 824 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_374
timestamp 1677677812
transform 1 0 832 0 1 570
box -8 -3 46 105
use FILL  FILL_9854
timestamp 1677677812
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_9857
timestamp 1677677812
transform 1 0 880 0 1 570
box -8 -3 16 105
use FILL  FILL_9859
timestamp 1677677812
transform 1 0 888 0 1 570
box -8 -3 16 105
use FILL  FILL_9861
timestamp 1677677812
transform 1 0 896 0 1 570
box -8 -3 16 105
use FILL  FILL_9862
timestamp 1677677812
transform 1 0 904 0 1 570
box -8 -3 16 105
use FILL  FILL_9863
timestamp 1677677812
transform 1 0 912 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7890
timestamp 1677677812
transform 1 0 1020 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_532
timestamp 1677677812
transform -1 0 1016 0 1 570
box -8 -3 104 105
use FILL  FILL_9864
timestamp 1677677812
transform 1 0 1016 0 1 570
box -8 -3 16 105
use FILL  FILL_9865
timestamp 1677677812
transform 1 0 1024 0 1 570
box -8 -3 16 105
use FILL  FILL_9866
timestamp 1677677812
transform 1 0 1032 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_97
timestamp 1677677812
transform 1 0 1040 0 1 570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_533
timestamp 1677677812
transform 1 0 1064 0 1 570
box -8 -3 104 105
use INVX2  INVX2_625
timestamp 1677677812
transform -1 0 1176 0 1 570
box -9 -3 26 105
use AOI22X1  AOI22X1_376
timestamp 1677677812
transform 1 0 1176 0 1 570
box -8 -3 46 105
use FILL  FILL_9867
timestamp 1677677812
transform 1 0 1216 0 1 570
box -8 -3 16 105
use FILL  FILL_9881
timestamp 1677677812
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_9883
timestamp 1677677812
transform 1 0 1232 0 1 570
box -8 -3 16 105
use INVX2  INVX2_627
timestamp 1677677812
transform -1 0 1256 0 1 570
box -9 -3 26 105
use FILL  FILL_9884
timestamp 1677677812
transform 1 0 1256 0 1 570
box -8 -3 16 105
use FILL  FILL_9885
timestamp 1677677812
transform 1 0 1264 0 1 570
box -8 -3 16 105
use FILL  FILL_9886
timestamp 1677677812
transform 1 0 1272 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_390
timestamp 1677677812
transform -1 0 1320 0 1 570
box -8 -3 46 105
use FILL  FILL_9887
timestamp 1677677812
transform 1 0 1320 0 1 570
box -8 -3 16 105
use FILL  FILL_9888
timestamp 1677677812
transform 1 0 1328 0 1 570
box -8 -3 16 105
use FILL  FILL_9889
timestamp 1677677812
transform 1 0 1336 0 1 570
box -8 -3 16 105
use FILL  FILL_9890
timestamp 1677677812
transform 1 0 1344 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7891
timestamp 1677677812
transform 1 0 1364 0 1 575
box -3 -3 3 3
use AOI22X1  AOI22X1_378
timestamp 1677677812
transform -1 0 1392 0 1 570
box -8 -3 46 105
use FILL  FILL_9891
timestamp 1677677812
transform 1 0 1392 0 1 570
box -8 -3 16 105
use FILL  FILL_9892
timestamp 1677677812
transform 1 0 1400 0 1 570
box -8 -3 16 105
use FILL  FILL_9893
timestamp 1677677812
transform 1 0 1408 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_379
timestamp 1677677812
transform -1 0 1456 0 1 570
box -8 -3 46 105
use INVX2  INVX2_628
timestamp 1677677812
transform 1 0 1456 0 1 570
box -9 -3 26 105
use FILL  FILL_9894
timestamp 1677677812
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_9895
timestamp 1677677812
transform 1 0 1480 0 1 570
box -8 -3 16 105
use FILL  FILL_9896
timestamp 1677677812
transform 1 0 1488 0 1 570
box -8 -3 16 105
use FILL  FILL_9897
timestamp 1677677812
transform 1 0 1496 0 1 570
box -8 -3 16 105
use FILL  FILL_9898
timestamp 1677677812
transform 1 0 1504 0 1 570
box -8 -3 16 105
use INVX2  INVX2_629
timestamp 1677677812
transform 1 0 1512 0 1 570
box -9 -3 26 105
use FILL  FILL_9899
timestamp 1677677812
transform 1 0 1528 0 1 570
box -8 -3 16 105
use FILL  FILL_9900
timestamp 1677677812
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_9901
timestamp 1677677812
transform 1 0 1544 0 1 570
box -8 -3 16 105
use INVX2  INVX2_630
timestamp 1677677812
transform -1 0 1568 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_7892
timestamp 1677677812
transform 1 0 1588 0 1 575
box -3 -3 3 3
use INVX2  INVX2_631
timestamp 1677677812
transform 1 0 1568 0 1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_535
timestamp 1677677812
transform -1 0 1680 0 1 570
box -8 -3 104 105
use OAI22X1  OAI22X1_391
timestamp 1677677812
transform 1 0 1680 0 1 570
box -8 -3 46 105
use FILL  FILL_9902
timestamp 1677677812
transform 1 0 1720 0 1 570
box -8 -3 16 105
use FILL  FILL_9922
timestamp 1677677812
transform 1 0 1728 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_381
timestamp 1677677812
transform 1 0 1736 0 1 570
box -8 -3 46 105
use AOI22X1  AOI22X1_382
timestamp 1677677812
transform -1 0 1816 0 1 570
box -8 -3 46 105
use INVX2  INVX2_633
timestamp 1677677812
transform 1 0 1816 0 1 570
box -9 -3 26 105
use FILL  FILL_9924
timestamp 1677677812
transform 1 0 1832 0 1 570
box -8 -3 16 105
use FILL  FILL_9936
timestamp 1677677812
transform 1 0 1840 0 1 570
box -8 -3 16 105
use FILL  FILL_9937
timestamp 1677677812
transform 1 0 1848 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7893
timestamp 1677677812
transform 1 0 1956 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_537
timestamp 1677677812
transform -1 0 1952 0 1 570
box -8 -3 104 105
use INVX2  INVX2_635
timestamp 1677677812
transform 1 0 1952 0 1 570
box -9 -3 26 105
use M3_M2  M3_M2_7894
timestamp 1677677812
transform 1 0 2004 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_7895
timestamp 1677677812
transform 1 0 2028 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_538
timestamp 1677677812
transform -1 0 2064 0 1 570
box -8 -3 104 105
use FILL  FILL_9938
timestamp 1677677812
transform 1 0 2064 0 1 570
box -8 -3 16 105
use FILL  FILL_9939
timestamp 1677677812
transform 1 0 2072 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_540
timestamp 1677677812
transform 1 0 2080 0 1 570
box -8 -3 104 105
use FILL  FILL_9949
timestamp 1677677812
transform 1 0 2176 0 1 570
box -8 -3 16 105
use FILL  FILL_9950
timestamp 1677677812
transform 1 0 2184 0 1 570
box -8 -3 16 105
use FILL  FILL_9951
timestamp 1677677812
transform 1 0 2192 0 1 570
box -8 -3 16 105
use FILL  FILL_9955
timestamp 1677677812
transform 1 0 2200 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_542
timestamp 1677677812
transform 1 0 2208 0 1 570
box -8 -3 104 105
use FILL  FILL_9957
timestamp 1677677812
transform 1 0 2304 0 1 570
box -8 -3 16 105
use FILL  FILL_9971
timestamp 1677677812
transform 1 0 2312 0 1 570
box -8 -3 16 105
use FILL  FILL_9973
timestamp 1677677812
transform 1 0 2320 0 1 570
box -8 -3 16 105
use FILL  FILL_9975
timestamp 1677677812
transform 1 0 2328 0 1 570
box -8 -3 16 105
use FILL  FILL_9977
timestamp 1677677812
transform 1 0 2336 0 1 570
box -8 -3 16 105
use FILL  FILL_9979
timestamp 1677677812
transform 1 0 2344 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_175
timestamp 1677677812
transform -1 0 2384 0 1 570
box -8 -3 34 105
use FILL  FILL_9980
timestamp 1677677812
transform 1 0 2384 0 1 570
box -8 -3 16 105
use FILL  FILL_9981
timestamp 1677677812
transform 1 0 2392 0 1 570
box -8 -3 16 105
use FILL  FILL_9982
timestamp 1677677812
transform 1 0 2400 0 1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_19
timestamp 1677677812
transform 1 0 2408 0 1 570
box -7 -3 39 105
use FILL  FILL_9983
timestamp 1677677812
transform 1 0 2440 0 1 570
box -8 -3 16 105
use FILL  FILL_9987
timestamp 1677677812
transform 1 0 2448 0 1 570
box -8 -3 16 105
use FILL  FILL_9988
timestamp 1677677812
transform 1 0 2456 0 1 570
box -8 -3 16 105
use INVX2  INVX2_638
timestamp 1677677812
transform -1 0 2480 0 1 570
box -9 -3 26 105
use FILL  FILL_9989
timestamp 1677677812
transform 1 0 2480 0 1 570
box -8 -3 16 105
use FILL  FILL_9990
timestamp 1677677812
transform 1 0 2488 0 1 570
box -8 -3 16 105
use FILL  FILL_9991
timestamp 1677677812
transform 1 0 2496 0 1 570
box -8 -3 16 105
use FILL  FILL_9992
timestamp 1677677812
transform 1 0 2504 0 1 570
box -8 -3 16 105
use FILL  FILL_9993
timestamp 1677677812
transform 1 0 2512 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_102
timestamp 1677677812
transform 1 0 2520 0 1 570
box -8 -3 32 105
use INVX2  INVX2_639
timestamp 1677677812
transform -1 0 2560 0 1 570
box -9 -3 26 105
use FILL  FILL_9994
timestamp 1677677812
transform 1 0 2560 0 1 570
box -8 -3 16 105
use FILL  FILL_9995
timestamp 1677677812
transform 1 0 2568 0 1 570
box -8 -3 16 105
use FILL  FILL_9996
timestamp 1677677812
transform 1 0 2576 0 1 570
box -8 -3 16 105
use FILL  FILL_9998
timestamp 1677677812
transform 1 0 2584 0 1 570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_1
timestamp 1677677812
transform 1 0 2592 0 1 570
box -8 -3 64 105
use FILL  FILL_9999
timestamp 1677677812
transform 1 0 2648 0 1 570
box -8 -3 16 105
use FILL  FILL_10000
timestamp 1677677812
transform 1 0 2656 0 1 570
box -8 -3 16 105
use FILL  FILL_10001
timestamp 1677677812
transform 1 0 2664 0 1 570
box -8 -3 16 105
use FILL  FILL_10002
timestamp 1677677812
transform 1 0 2672 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_544
timestamp 1677677812
transform -1 0 2776 0 1 570
box -8 -3 104 105
use FILL  FILL_10003
timestamp 1677677812
transform 1 0 2776 0 1 570
box -8 -3 16 105
use FILL  FILL_10004
timestamp 1677677812
transform 1 0 2784 0 1 570
box -8 -3 16 105
use FILL  FILL_10007
timestamp 1677677812
transform 1 0 2792 0 1 570
box -8 -3 16 105
use FILL  FILL_10008
timestamp 1677677812
transform 1 0 2800 0 1 570
box -8 -3 16 105
use FILL  FILL_10009
timestamp 1677677812
transform 1 0 2808 0 1 570
box -8 -3 16 105
use FILL  FILL_10010
timestamp 1677677812
transform 1 0 2816 0 1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_7
timestamp 1677677812
transform -1 0 2880 0 1 570
box -8 -3 64 105
use FILL  FILL_10011
timestamp 1677677812
transform 1 0 2880 0 1 570
box -8 -3 16 105
use FILL  FILL_10012
timestamp 1677677812
transform 1 0 2888 0 1 570
box -8 -3 16 105
use FILL  FILL_10013
timestamp 1677677812
transform 1 0 2896 0 1 570
box -8 -3 16 105
use BUFX2  BUFX2_113
timestamp 1677677812
transform 1 0 2904 0 1 570
box -5 -3 28 105
use FILL  FILL_10016
timestamp 1677677812
transform 1 0 2928 0 1 570
box -8 -3 16 105
use FILL  FILL_10018
timestamp 1677677812
transform 1 0 2936 0 1 570
box -8 -3 16 105
use FILL  FILL_10019
timestamp 1677677812
transform 1 0 2944 0 1 570
box -8 -3 16 105
use FILL  FILL_10020
timestamp 1677677812
transform 1 0 2952 0 1 570
box -8 -3 16 105
use FILL  FILL_10021
timestamp 1677677812
transform 1 0 2960 0 1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_75
timestamp 1677677812
transform -1 0 3000 0 1 570
box -8 -3 40 105
use FILL  FILL_10022
timestamp 1677677812
transform 1 0 3000 0 1 570
box -8 -3 16 105
use FILL  FILL_10023
timestamp 1677677812
transform 1 0 3008 0 1 570
box -8 -3 16 105
use INVX2  INVX2_640
timestamp 1677677812
transform -1 0 3032 0 1 570
box -9 -3 26 105
use FILL  FILL_10024
timestamp 1677677812
transform 1 0 3032 0 1 570
box -8 -3 16 105
use FILL  FILL_10032
timestamp 1677677812
transform 1 0 3040 0 1 570
box -8 -3 16 105
use FILL  FILL_10033
timestamp 1677677812
transform 1 0 3048 0 1 570
box -8 -3 16 105
use FILL  FILL_10034
timestamp 1677677812
transform 1 0 3056 0 1 570
box -8 -3 16 105
use FILL  FILL_10035
timestamp 1677677812
transform 1 0 3064 0 1 570
box -8 -3 16 105
use FILL  FILL_10037
timestamp 1677677812
transform 1 0 3072 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_106
timestamp 1677677812
transform 1 0 3080 0 1 570
box -8 -3 32 105
use FILL  FILL_10039
timestamp 1677677812
transform 1 0 3104 0 1 570
box -8 -3 16 105
use FILL  FILL_10040
timestamp 1677677812
transform 1 0 3112 0 1 570
box -8 -3 16 105
use AND2X2  AND2X2_62
timestamp 1677677812
transform -1 0 3152 0 1 570
box -8 -3 40 105
use FILL  FILL_10041
timestamp 1677677812
transform 1 0 3152 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_107
timestamp 1677677812
transform -1 0 3184 0 1 570
box -8 -3 32 105
use FILL  FILL_10042
timestamp 1677677812
transform 1 0 3184 0 1 570
box -8 -3 16 105
use FILL  FILL_10043
timestamp 1677677812
transform 1 0 3192 0 1 570
box -8 -3 16 105
use FILL  FILL_10044
timestamp 1677677812
transform 1 0 3200 0 1 570
box -8 -3 16 105
use FILL  FILL_10045
timestamp 1677677812
transform 1 0 3208 0 1 570
box -8 -3 16 105
use FILL  FILL_10046
timestamp 1677677812
transform 1 0 3216 0 1 570
box -8 -3 16 105
use FILL  FILL_10047
timestamp 1677677812
transform 1 0 3224 0 1 570
box -8 -3 16 105
use FILL  FILL_10048
timestamp 1677677812
transform 1 0 3232 0 1 570
box -8 -3 16 105
use FILL  FILL_10049
timestamp 1677677812
transform 1 0 3240 0 1 570
box -8 -3 16 105
use FILL  FILL_10050
timestamp 1677677812
transform 1 0 3248 0 1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_108
timestamp 1677677812
transform 1 0 3256 0 1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_109
timestamp 1677677812
transform 1 0 3280 0 1 570
box -8 -3 32 105
use FILL  FILL_10051
timestamp 1677677812
transform 1 0 3304 0 1 570
box -8 -3 16 105
use FILL  FILL_10052
timestamp 1677677812
transform 1 0 3312 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_548
timestamp 1677677812
transform 1 0 3320 0 1 570
box -8 -3 104 105
use M3_M2  M3_M2_7896
timestamp 1677677812
transform 1 0 3484 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_549
timestamp 1677677812
transform 1 0 3416 0 1 570
box -8 -3 104 105
use FILL  FILL_10053
timestamp 1677677812
transform 1 0 3512 0 1 570
box -8 -3 16 105
use FILL  FILL_10074
timestamp 1677677812
transform 1 0 3520 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_43
timestamp 1677677812
transform 1 0 3528 0 1 570
box -8 -3 32 105
use FILL  FILL_10075
timestamp 1677677812
transform 1 0 3552 0 1 570
box -8 -3 16 105
use FILL  FILL_10076
timestamp 1677677812
transform 1 0 3560 0 1 570
box -8 -3 16 105
use FILL  FILL_10077
timestamp 1677677812
transform 1 0 3568 0 1 570
box -8 -3 16 105
use FILL  FILL_10078
timestamp 1677677812
transform 1 0 3576 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_395
timestamp 1677677812
transform 1 0 3584 0 1 570
box -8 -3 46 105
use FILL  FILL_10079
timestamp 1677677812
transform 1 0 3624 0 1 570
box -8 -3 16 105
use FILL  FILL_10080
timestamp 1677677812
transform 1 0 3632 0 1 570
box -8 -3 16 105
use INVX2  INVX2_641
timestamp 1677677812
transform -1 0 3656 0 1 570
box -9 -3 26 105
use FILL  FILL_10081
timestamp 1677677812
transform 1 0 3656 0 1 570
box -8 -3 16 105
use FILL  FILL_10082
timestamp 1677677812
transform 1 0 3664 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_396
timestamp 1677677812
transform 1 0 3672 0 1 570
box -8 -3 46 105
use FILL  FILL_10084
timestamp 1677677812
transform 1 0 3712 0 1 570
box -8 -3 16 105
use FILL  FILL_10085
timestamp 1677677812
transform 1 0 3720 0 1 570
box -8 -3 16 105
use FILL  FILL_10086
timestamp 1677677812
transform 1 0 3728 0 1 570
box -8 -3 16 105
use FILL  FILL_10090
timestamp 1677677812
transform 1 0 3736 0 1 570
box -8 -3 16 105
use FILL  FILL_10092
timestamp 1677677812
transform 1 0 3744 0 1 570
box -8 -3 16 105
use FILL  FILL_10093
timestamp 1677677812
transform 1 0 3752 0 1 570
box -8 -3 16 105
use FILL  FILL_10094
timestamp 1677677812
transform 1 0 3760 0 1 570
box -8 -3 16 105
use FILL  FILL_10095
timestamp 1677677812
transform 1 0 3768 0 1 570
box -8 -3 16 105
use FILL  FILL_10096
timestamp 1677677812
transform 1 0 3776 0 1 570
box -8 -3 16 105
use FILL  FILL_10097
timestamp 1677677812
transform 1 0 3784 0 1 570
box -8 -3 16 105
use FILL  FILL_10098
timestamp 1677677812
transform 1 0 3792 0 1 570
box -8 -3 16 105
use INVX2  INVX2_642
timestamp 1677677812
transform -1 0 3816 0 1 570
box -9 -3 26 105
use FILL  FILL_10099
timestamp 1677677812
transform 1 0 3816 0 1 570
box -8 -3 16 105
use FILL  FILL_10105
timestamp 1677677812
transform 1 0 3824 0 1 570
box -8 -3 16 105
use FILL  FILL_10107
timestamp 1677677812
transform 1 0 3832 0 1 570
box -8 -3 16 105
use FILL  FILL_10109
timestamp 1677677812
transform 1 0 3840 0 1 570
box -8 -3 16 105
use FILL  FILL_10110
timestamp 1677677812
transform 1 0 3848 0 1 570
box -8 -3 16 105
use FILL  FILL_10111
timestamp 1677677812
transform 1 0 3856 0 1 570
box -8 -3 16 105
use FILL  FILL_10113
timestamp 1677677812
transform 1 0 3864 0 1 570
box -8 -3 16 105
use FILL  FILL_10115
timestamp 1677677812
transform 1 0 3872 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_399
timestamp 1677677812
transform -1 0 3920 0 1 570
box -8 -3 46 105
use FILL  FILL_10117
timestamp 1677677812
transform 1 0 3920 0 1 570
box -8 -3 16 105
use FILL  FILL_10119
timestamp 1677677812
transform 1 0 3928 0 1 570
box -8 -3 16 105
use FILL  FILL_10121
timestamp 1677677812
transform 1 0 3936 0 1 570
box -8 -3 16 105
use FILL  FILL_10123
timestamp 1677677812
transform 1 0 3944 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_401
timestamp 1677677812
transform -1 0 3992 0 1 570
box -8 -3 46 105
use FILL  FILL_10124
timestamp 1677677812
transform 1 0 3992 0 1 570
box -8 -3 16 105
use FILL  FILL_10130
timestamp 1677677812
transform 1 0 4000 0 1 570
box -8 -3 16 105
use FILL  FILL_10131
timestamp 1677677812
transform 1 0 4008 0 1 570
box -8 -3 16 105
use FILL  FILL_10132
timestamp 1677677812
transform 1 0 4016 0 1 570
box -8 -3 16 105
use FILL  FILL_10133
timestamp 1677677812
transform 1 0 4024 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_402
timestamp 1677677812
transform -1 0 4072 0 1 570
box -8 -3 46 105
use FILL  FILL_10134
timestamp 1677677812
transform 1 0 4072 0 1 570
box -8 -3 16 105
use FILL  FILL_10135
timestamp 1677677812
transform 1 0 4080 0 1 570
box -8 -3 16 105
use FILL  FILL_10136
timestamp 1677677812
transform 1 0 4088 0 1 570
box -8 -3 16 105
use FILL  FILL_10137
timestamp 1677677812
transform 1 0 4096 0 1 570
box -8 -3 16 105
use FILL  FILL_10138
timestamp 1677677812
transform 1 0 4104 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_403
timestamp 1677677812
transform -1 0 4152 0 1 570
box -8 -3 46 105
use FILL  FILL_10139
timestamp 1677677812
transform 1 0 4152 0 1 570
box -8 -3 16 105
use FILL  FILL_10140
timestamp 1677677812
transform 1 0 4160 0 1 570
box -8 -3 16 105
use FILL  FILL_10141
timestamp 1677677812
transform 1 0 4168 0 1 570
box -8 -3 16 105
use FILL  FILL_10142
timestamp 1677677812
transform 1 0 4176 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7897
timestamp 1677677812
transform 1 0 4220 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_404
timestamp 1677677812
transform 1 0 4184 0 1 570
box -8 -3 46 105
use FILL  FILL_10143
timestamp 1677677812
transform 1 0 4224 0 1 570
box -8 -3 16 105
use FILL  FILL_10144
timestamp 1677677812
transform 1 0 4232 0 1 570
box -8 -3 16 105
use FILL  FILL_10145
timestamp 1677677812
transform 1 0 4240 0 1 570
box -8 -3 16 105
use FILL  FILL_10146
timestamp 1677677812
transform 1 0 4248 0 1 570
box -8 -3 16 105
use FILL  FILL_10147
timestamp 1677677812
transform 1 0 4256 0 1 570
box -8 -3 16 105
use FILL  FILL_10148
timestamp 1677677812
transform 1 0 4264 0 1 570
box -8 -3 16 105
use FILL  FILL_10149
timestamp 1677677812
transform 1 0 4272 0 1 570
box -8 -3 16 105
use FILL  FILL_10150
timestamp 1677677812
transform 1 0 4280 0 1 570
box -8 -3 16 105
use FILL  FILL_10159
timestamp 1677677812
transform 1 0 4288 0 1 570
box -8 -3 16 105
use FILL  FILL_10161
timestamp 1677677812
transform 1 0 4296 0 1 570
box -8 -3 16 105
use FILL  FILL_10162
timestamp 1677677812
transform 1 0 4304 0 1 570
box -8 -3 16 105
use FILL  FILL_10163
timestamp 1677677812
transform 1 0 4312 0 1 570
box -8 -3 16 105
use FILL  FILL_10164
timestamp 1677677812
transform 1 0 4320 0 1 570
box -8 -3 16 105
use FILL  FILL_10165
timestamp 1677677812
transform 1 0 4328 0 1 570
box -8 -3 16 105
use FILL  FILL_10166
timestamp 1677677812
transform 1 0 4336 0 1 570
box -8 -3 16 105
use FILL  FILL_10167
timestamp 1677677812
transform 1 0 4344 0 1 570
box -8 -3 16 105
use FILL  FILL_10168
timestamp 1677677812
transform 1 0 4352 0 1 570
box -8 -3 16 105
use FILL  FILL_10170
timestamp 1677677812
transform 1 0 4360 0 1 570
box -8 -3 16 105
use FILL  FILL_10172
timestamp 1677677812
transform 1 0 4368 0 1 570
box -8 -3 16 105
use FILL  FILL_10173
timestamp 1677677812
transform 1 0 4376 0 1 570
box -8 -3 16 105
use INVX2  INVX2_649
timestamp 1677677812
transform -1 0 4400 0 1 570
box -9 -3 26 105
use FILL  FILL_10174
timestamp 1677677812
transform 1 0 4400 0 1 570
box -8 -3 16 105
use FILL  FILL_10175
timestamp 1677677812
transform 1 0 4408 0 1 570
box -8 -3 16 105
use FILL  FILL_10176
timestamp 1677677812
transform 1 0 4416 0 1 570
box -8 -3 16 105
use FILL  FILL_10177
timestamp 1677677812
transform 1 0 4424 0 1 570
box -8 -3 16 105
use FILL  FILL_10178
timestamp 1677677812
transform 1 0 4432 0 1 570
box -8 -3 16 105
use FILL  FILL_10179
timestamp 1677677812
transform 1 0 4440 0 1 570
box -8 -3 16 105
use FILL  FILL_10180
timestamp 1677677812
transform 1 0 4448 0 1 570
box -8 -3 16 105
use FILL  FILL_10181
timestamp 1677677812
transform 1 0 4456 0 1 570
box -8 -3 16 105
use FILL  FILL_10182
timestamp 1677677812
transform 1 0 4464 0 1 570
box -8 -3 16 105
use FILL  FILL_10183
timestamp 1677677812
transform 1 0 4472 0 1 570
box -8 -3 16 105
use FILL  FILL_10186
timestamp 1677677812
transform 1 0 4480 0 1 570
box -8 -3 16 105
use INVX2  INVX2_650
timestamp 1677677812
transform -1 0 4504 0 1 570
box -9 -3 26 105
use FILL  FILL_10187
timestamp 1677677812
transform 1 0 4504 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_7898
timestamp 1677677812
transform 1 0 4540 0 1 575
box -3 -3 3 3
use M3_M2  M3_M2_7899
timestamp 1677677812
transform 1 0 4556 0 1 575
box -3 -3 3 3
use OAI22X1  OAI22X1_408
timestamp 1677677812
transform 1 0 4512 0 1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_409
timestamp 1677677812
transform 1 0 4552 0 1 570
box -8 -3 46 105
use FILL  FILL_10188
timestamp 1677677812
transform 1 0 4592 0 1 570
box -8 -3 16 105
use FILL  FILL_10189
timestamp 1677677812
transform 1 0 4600 0 1 570
box -8 -3 16 105
use FILL  FILL_10194
timestamp 1677677812
transform 1 0 4608 0 1 570
box -8 -3 16 105
use FILL  FILL_10195
timestamp 1677677812
transform 1 0 4616 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_410
timestamp 1677677812
transform 1 0 4624 0 1 570
box -8 -3 46 105
use FILL  FILL_10196
timestamp 1677677812
transform 1 0 4664 0 1 570
box -8 -3 16 105
use FILL  FILL_10197
timestamp 1677677812
transform 1 0 4672 0 1 570
box -8 -3 16 105
use FILL  FILL_10198
timestamp 1677677812
transform 1 0 4680 0 1 570
box -8 -3 16 105
use FILL  FILL_10199
timestamp 1677677812
transform 1 0 4688 0 1 570
box -8 -3 16 105
use FILL  FILL_10200
timestamp 1677677812
transform 1 0 4696 0 1 570
box -8 -3 16 105
use FILL  FILL_10201
timestamp 1677677812
transform 1 0 4704 0 1 570
box -8 -3 16 105
use INVX2  INVX2_651
timestamp 1677677812
transform -1 0 4728 0 1 570
box -9 -3 26 105
use FILL  FILL_10202
timestamp 1677677812
transform 1 0 4728 0 1 570
box -8 -3 16 105
use FILL  FILL_10203
timestamp 1677677812
transform 1 0 4736 0 1 570
box -8 -3 16 105
use FILL  FILL_10204
timestamp 1677677812
transform 1 0 4744 0 1 570
box -8 -3 16 105
use FILL  FILL_10205
timestamp 1677677812
transform 1 0 4752 0 1 570
box -8 -3 16 105
use FILL  FILL_10206
timestamp 1677677812
transform 1 0 4760 0 1 570
box -8 -3 16 105
use FILL  FILL_10207
timestamp 1677677812
transform 1 0 4768 0 1 570
box -8 -3 16 105
use FILL  FILL_10208
timestamp 1677677812
transform 1 0 4776 0 1 570
box -8 -3 16 105
use FILL  FILL_10209
timestamp 1677677812
transform 1 0 4784 0 1 570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_83
timestamp 1677677812
transform 1 0 4819 0 1 570
box -10 -3 10 3
use M3_M2  M3_M2_8065
timestamp 1677677812
transform 1 0 84 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7935
timestamp 1677677812
transform 1 0 100 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8910
timestamp 1677677812
transform 1 0 100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9022
timestamp 1677677812
transform 1 0 108 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7983
timestamp 1677677812
transform 1 0 132 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8911
timestamp 1677677812
transform 1 0 164 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7984
timestamp 1677677812
transform 1 0 172 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7936
timestamp 1677677812
transform 1 0 220 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8912
timestamp 1677677812
transform 1 0 196 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8913
timestamp 1677677812
transform 1 0 204 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8005
timestamp 1677677812
transform 1 0 164 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7985
timestamp 1677677812
transform 1 0 212 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9023
timestamp 1677677812
transform 1 0 172 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9024
timestamp 1677677812
transform 1 0 188 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9025
timestamp 1677677812
transform 1 0 204 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9026
timestamp 1677677812
transform 1 0 212 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8026
timestamp 1677677812
transform 1 0 196 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8027
timestamp 1677677812
transform 1 0 212 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8085
timestamp 1677677812
transform 1 0 204 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7937
timestamp 1677677812
transform 1 0 348 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8914
timestamp 1677677812
transform 1 0 236 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8915
timestamp 1677677812
transform 1 0 252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8916
timestamp 1677677812
transform 1 0 268 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9027
timestamp 1677677812
transform 1 0 244 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8006
timestamp 1677677812
transform 1 0 252 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7914
timestamp 1677677812
transform 1 0 372 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9028
timestamp 1677677812
transform 1 0 316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9029
timestamp 1677677812
transform 1 0 348 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9030
timestamp 1677677812
transform 1 0 356 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9031
timestamp 1677677812
transform 1 0 364 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8028
timestamp 1677677812
transform 1 0 244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8066
timestamp 1677677812
transform 1 0 252 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8086
timestamp 1677677812
transform 1 0 228 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_8917
timestamp 1677677812
transform 1 0 388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8918
timestamp 1677677812
transform 1 0 396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8919
timestamp 1677677812
transform 1 0 412 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8007
timestamp 1677677812
transform 1 0 396 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9032
timestamp 1677677812
transform 1 0 404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8920
timestamp 1677677812
transform 1 0 444 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9033
timestamp 1677677812
transform 1 0 436 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8008
timestamp 1677677812
transform 1 0 444 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8067
timestamp 1677677812
transform 1 0 436 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7900
timestamp 1677677812
transform 1 0 468 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7915
timestamp 1677677812
transform 1 0 492 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7938
timestamp 1677677812
transform 1 0 492 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8921
timestamp 1677677812
transform 1 0 468 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7986
timestamp 1677677812
transform 1 0 476 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8922
timestamp 1677677812
transform 1 0 484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8923
timestamp 1677677812
transform 1 0 492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8924
timestamp 1677677812
transform 1 0 508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9034
timestamp 1677677812
transform 1 0 460 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9035
timestamp 1677677812
transform 1 0 476 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8029
timestamp 1677677812
transform 1 0 460 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8068
timestamp 1677677812
transform 1 0 460 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7987
timestamp 1677677812
transform 1 0 516 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7916
timestamp 1677677812
transform 1 0 660 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7939
timestamp 1677677812
transform 1 0 620 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7940
timestamp 1677677812
transform 1 0 636 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8925
timestamp 1677677812
transform 1 0 524 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8926
timestamp 1677677812
transform 1 0 540 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9036
timestamp 1677677812
transform 1 0 500 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8009
timestamp 1677677812
transform 1 0 508 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9037
timestamp 1677677812
transform 1 0 516 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8030
timestamp 1677677812
transform 1 0 500 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8069
timestamp 1677677812
transform 1 0 516 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8087
timestamp 1677677812
transform 1 0 500 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7988
timestamp 1677677812
transform 1 0 588 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8927
timestamp 1677677812
transform 1 0 628 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8928
timestamp 1677677812
transform 1 0 636 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8929
timestamp 1677677812
transform 1 0 652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8930
timestamp 1677677812
transform 1 0 660 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9038
timestamp 1677677812
transform 1 0 588 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9039
timestamp 1677677812
transform 1 0 620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9040
timestamp 1677677812
transform 1 0 644 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8031
timestamp 1677677812
transform 1 0 644 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7989
timestamp 1677677812
transform 1 0 668 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9041
timestamp 1677677812
transform 1 0 668 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8931
timestamp 1677677812
transform 1 0 684 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8032
timestamp 1677677812
transform 1 0 684 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9042
timestamp 1677677812
transform 1 0 708 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7941
timestamp 1677677812
transform 1 0 732 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8932
timestamp 1677677812
transform 1 0 724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8933
timestamp 1677677812
transform 1 0 732 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9043
timestamp 1677677812
transform 1 0 732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9044
timestamp 1677677812
transform 1 0 740 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8033
timestamp 1677677812
transform 1 0 732 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8034
timestamp 1677677812
transform 1 0 748 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7917
timestamp 1677677812
transform 1 0 772 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8934
timestamp 1677677812
transform 1 0 772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9045
timestamp 1677677812
transform 1 0 780 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8070
timestamp 1677677812
transform 1 0 756 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8088
timestamp 1677677812
transform 1 0 756 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8089
timestamp 1677677812
transform 1 0 780 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9136
timestamp 1677677812
transform 1 0 796 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_7942
timestamp 1677677812
transform 1 0 812 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8935
timestamp 1677677812
transform 1 0 812 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8936
timestamp 1677677812
transform 1 0 820 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8937
timestamp 1677677812
transform 1 0 836 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8938
timestamp 1677677812
transform 1 0 844 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9046
timestamp 1677677812
transform 1 0 828 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9047
timestamp 1677677812
transform 1 0 844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9048
timestamp 1677677812
transform 1 0 852 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8071
timestamp 1677677812
transform 1 0 828 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8072
timestamp 1677677812
transform 1 0 844 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8098
timestamp 1677677812
transform 1 0 812 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_7943
timestamp 1677677812
transform 1 0 868 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8939
timestamp 1677677812
transform 1 0 868 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9049
timestamp 1677677812
transform 1 0 868 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8073
timestamp 1677677812
transform 1 0 868 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8090
timestamp 1677677812
transform 1 0 860 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9050
timestamp 1677677812
transform 1 0 876 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8940
timestamp 1677677812
transform 1 0 892 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8099
timestamp 1677677812
transform 1 0 900 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_8941
timestamp 1677677812
transform 1 0 932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8942
timestamp 1677677812
transform 1 0 940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9051
timestamp 1677677812
transform 1 0 924 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8074
timestamp 1677677812
transform 1 0 916 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7990
timestamp 1677677812
transform 1 0 956 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9052
timestamp 1677677812
transform 1 0 956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9053
timestamp 1677677812
transform 1 0 964 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8903
timestamp 1677677812
transform 1 0 980 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_8010
timestamp 1677677812
transform 1 0 980 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7918
timestamp 1677677812
transform 1 0 1028 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7944
timestamp 1677677812
transform 1 0 1020 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8904
timestamp 1677677812
transform 1 0 1028 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8943
timestamp 1677677812
transform 1 0 1020 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7945
timestamp 1677677812
transform 1 0 1044 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9054
timestamp 1677677812
transform 1 0 1036 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8011
timestamp 1677677812
transform 1 0 1044 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7919
timestamp 1677677812
transform 1 0 1068 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8944
timestamp 1677677812
transform 1 0 1060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9055
timestamp 1677677812
transform 1 0 1068 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7946
timestamp 1677677812
transform 1 0 1172 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8905
timestamp 1677677812
transform 1 0 1180 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8945
timestamp 1677677812
transform 1 0 1084 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7991
timestamp 1677677812
transform 1 0 1132 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7992
timestamp 1677677812
transform 1 0 1164 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9056
timestamp 1677677812
transform 1 0 1132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9057
timestamp 1677677812
transform 1 0 1188 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8035
timestamp 1677677812
transform 1 0 1180 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7901
timestamp 1677677812
transform 1 0 1212 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7947
timestamp 1677677812
transform 1 0 1204 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8906
timestamp 1677677812
transform 1 0 1212 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8946
timestamp 1677677812
transform 1 0 1236 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7948
timestamp 1677677812
transform 1 0 1260 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8947
timestamp 1677677812
transform 1 0 1252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8948
timestamp 1677677812
transform 1 0 1260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9058
timestamp 1677677812
transform 1 0 1244 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8036
timestamp 1677677812
transform 1 0 1244 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8091
timestamp 1677677812
transform 1 0 1236 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9059
timestamp 1677677812
transform 1 0 1268 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7920
timestamp 1677677812
transform 1 0 1292 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8949
timestamp 1677677812
transform 1 0 1292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9060
timestamp 1677677812
transform 1 0 1284 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9061
timestamp 1677677812
transform 1 0 1308 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8037
timestamp 1677677812
transform 1 0 1292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8038
timestamp 1677677812
transform 1 0 1308 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8075
timestamp 1677677812
transform 1 0 1284 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7949
timestamp 1677677812
transform 1 0 1324 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8950
timestamp 1677677812
transform 1 0 1324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8951
timestamp 1677677812
transform 1 0 1332 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7993
timestamp 1677677812
transform 1 0 1340 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8952
timestamp 1677677812
transform 1 0 1348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8953
timestamp 1677677812
transform 1 0 1364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9062
timestamp 1677677812
transform 1 0 1340 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9063
timestamp 1677677812
transform 1 0 1356 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8039
timestamp 1677677812
transform 1 0 1356 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8076
timestamp 1677677812
transform 1 0 1340 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8092
timestamp 1677677812
transform 1 0 1380 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7902
timestamp 1677677812
transform 1 0 1388 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_8954
timestamp 1677677812
transform 1 0 1388 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7903
timestamp 1677677812
transform 1 0 1412 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7921
timestamp 1677677812
transform 1 0 1404 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_9064
timestamp 1677677812
transform 1 0 1404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9065
timestamp 1677677812
transform 1 0 1412 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8955
timestamp 1677677812
transform 1 0 1420 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7904
timestamp 1677677812
transform 1 0 1460 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7922
timestamp 1677677812
transform 1 0 1468 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7950
timestamp 1677677812
transform 1 0 1460 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7951
timestamp 1677677812
transform 1 0 1476 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8956
timestamp 1677677812
transform 1 0 1460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8957
timestamp 1677677812
transform 1 0 1556 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9066
timestamp 1677677812
transform 1 0 1436 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9067
timestamp 1677677812
transform 1 0 1452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9068
timestamp 1677677812
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9069
timestamp 1677677812
transform 1 0 1476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9070
timestamp 1677677812
transform 1 0 1524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8958
timestamp 1677677812
transform 1 0 1588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9071
timestamp 1677677812
transform 1 0 1612 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_8959
timestamp 1677677812
transform 1 0 1636 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8040
timestamp 1677677812
transform 1 0 1636 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7952
timestamp 1677677812
transform 1 0 1684 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8960
timestamp 1677677812
transform 1 0 1676 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8961
timestamp 1677677812
transform 1 0 1692 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7994
timestamp 1677677812
transform 1 0 1700 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9072
timestamp 1677677812
transform 1 0 1684 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8012
timestamp 1677677812
transform 1 0 1692 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9073
timestamp 1677677812
transform 1 0 1700 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8041
timestamp 1677677812
transform 1 0 1676 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8077
timestamp 1677677812
transform 1 0 1684 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7905
timestamp 1677677812
transform 1 0 1724 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_8078
timestamp 1677677812
transform 1 0 1716 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_8962
timestamp 1677677812
transform 1 0 1772 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8100
timestamp 1677677812
transform 1 0 1772 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_8963
timestamp 1677677812
transform 1 0 1788 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8013
timestamp 1677677812
transform 1 0 1812 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8101
timestamp 1677677812
transform 1 0 1812 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_8964
timestamp 1677677812
transform 1 0 1932 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9074
timestamp 1677677812
transform 1 0 1844 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9075
timestamp 1677677812
transform 1 0 1852 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9076
timestamp 1677677812
transform 1 0 1908 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8042
timestamp 1677677812
transform 1 0 1852 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8043
timestamp 1677677812
transform 1 0 1908 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8079
timestamp 1677677812
transform 1 0 1908 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7923
timestamp 1677677812
transform 1 0 1948 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8965
timestamp 1677677812
transform 1 0 1956 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9077
timestamp 1677677812
transform 1 0 1948 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8044
timestamp 1677677812
transform 1 0 1948 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7953
timestamp 1677677812
transform 1 0 1972 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8966
timestamp 1677677812
transform 1 0 1972 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9078
timestamp 1677677812
transform 1 0 1972 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8014
timestamp 1677677812
transform 1 0 1980 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7906
timestamp 1677677812
transform 1 0 2036 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7954
timestamp 1677677812
transform 1 0 2012 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8967
timestamp 1677677812
transform 1 0 2012 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8968
timestamp 1677677812
transform 1 0 2028 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8969
timestamp 1677677812
transform 1 0 2036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8970
timestamp 1677677812
transform 1 0 2044 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9079
timestamp 1677677812
transform 1 0 2020 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8015
timestamp 1677677812
transform 1 0 2028 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8016
timestamp 1677677812
transform 1 0 2044 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7924
timestamp 1677677812
transform 1 0 2060 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7907
timestamp 1677677812
transform 1 0 2076 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7995
timestamp 1677677812
transform 1 0 2084 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7908
timestamp 1677677812
transform 1 0 2124 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7925
timestamp 1677677812
transform 1 0 2180 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7955
timestamp 1677677812
transform 1 0 2100 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7996
timestamp 1677677812
transform 1 0 2132 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8971
timestamp 1677677812
transform 1 0 2180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9080
timestamp 1677677812
transform 1 0 2092 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9081
timestamp 1677677812
transform 1 0 2100 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9082
timestamp 1677677812
transform 1 0 2132 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8045
timestamp 1677677812
transform 1 0 2092 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8046
timestamp 1677677812
transform 1 0 2132 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8972
timestamp 1677677812
transform 1 0 2316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8973
timestamp 1677677812
transform 1 0 2348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9083
timestamp 1677677812
transform 1 0 2340 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7956
timestamp 1677677812
transform 1 0 2364 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8974
timestamp 1677677812
transform 1 0 2364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9084
timestamp 1677677812
transform 1 0 2388 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9137
timestamp 1677677812
transform 1 0 2380 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_8975
timestamp 1677677812
transform 1 0 2444 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8047
timestamp 1677677812
transform 1 0 2444 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_8976
timestamp 1677677812
transform 1 0 2460 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7957
timestamp 1677677812
transform 1 0 2572 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8977
timestamp 1677677812
transform 1 0 2572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9085
timestamp 1677677812
transform 1 0 2500 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9086
timestamp 1677677812
transform 1 0 2540 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9087
timestamp 1677677812
transform 1 0 2548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9088
timestamp 1677677812
transform 1 0 2564 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8048
timestamp 1677677812
transform 1 0 2564 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7958
timestamp 1677677812
transform 1 0 2588 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7959
timestamp 1677677812
transform 1 0 2676 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8978
timestamp 1677677812
transform 1 0 2676 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7909
timestamp 1677677812
transform 1 0 2748 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7960
timestamp 1677677812
transform 1 0 2732 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7961
timestamp 1677677812
transform 1 0 2772 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8979
timestamp 1677677812
transform 1 0 2772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9089
timestamp 1677677812
transform 1 0 2596 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9090
timestamp 1677677812
transform 1 0 2652 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9091
timestamp 1677677812
transform 1 0 2692 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9092
timestamp 1677677812
transform 1 0 2748 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8049
timestamp 1677677812
transform 1 0 2692 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7962
timestamp 1677677812
transform 1 0 2788 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7910
timestamp 1677677812
transform 1 0 2876 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7963
timestamp 1677677812
transform 1 0 2884 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8980
timestamp 1677677812
transform 1 0 2884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9093
timestamp 1677677812
transform 1 0 2804 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9094
timestamp 1677677812
transform 1 0 2860 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8050
timestamp 1677677812
transform 1 0 2860 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7926
timestamp 1677677812
transform 1 0 2908 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8907
timestamp 1677677812
transform 1 0 2908 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8981
timestamp 1677677812
transform 1 0 2900 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8051
timestamp 1677677812
transform 1 0 2900 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9138
timestamp 1677677812
transform 1 0 2948 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_7927
timestamp 1677677812
transform 1 0 2980 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8908
timestamp 1677677812
transform 1 0 2972 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8982
timestamp 1677677812
transform 1 0 2972 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8983
timestamp 1677677812
transform 1 0 2980 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8017
timestamp 1677677812
transform 1 0 2972 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8018
timestamp 1677677812
transform 1 0 3012 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9095
timestamp 1677677812
transform 1 0 3020 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7928
timestamp 1677677812
transform 1 0 3044 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8909
timestamp 1677677812
transform 1 0 3044 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_8984
timestamp 1677677812
transform 1 0 3052 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8019
timestamp 1677677812
transform 1 0 3068 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9139
timestamp 1677677812
transform 1 0 3068 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_9096
timestamp 1677677812
transform 1 0 3108 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8052
timestamp 1677677812
transform 1 0 3108 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9097
timestamp 1677677812
transform 1 0 3132 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9140
timestamp 1677677812
transform 1 0 3140 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_9144
timestamp 1677677812
transform 1 0 3124 0 1 505
box -2 -2 2 2
use M3_M2  M3_M2_8053
timestamp 1677677812
transform 1 0 3164 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7929
timestamp 1677677812
transform 1 0 3180 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7964
timestamp 1677677812
transform 1 0 3180 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8985
timestamp 1677677812
transform 1 0 3180 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9098
timestamp 1677677812
transform 1 0 3204 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8054
timestamp 1677677812
transform 1 0 3204 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7997
timestamp 1677677812
transform 1 0 3292 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9099
timestamp 1677677812
transform 1 0 3292 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7911
timestamp 1677677812
transform 1 0 3308 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7912
timestamp 1677677812
transform 1 0 3332 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7930
timestamp 1677677812
transform 1 0 3332 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7965
timestamp 1677677812
transform 1 0 3308 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8986
timestamp 1677677812
transform 1 0 3308 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7998
timestamp 1677677812
transform 1 0 3388 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8987
timestamp 1677677812
transform 1 0 3396 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9100
timestamp 1677677812
transform 1 0 3332 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7913
timestamp 1677677812
transform 1 0 3428 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_7966
timestamp 1677677812
transform 1 0 3428 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9101
timestamp 1677677812
transform 1 0 3428 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7999
timestamp 1677677812
transform 1 0 3452 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8988
timestamp 1677677812
transform 1 0 3460 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7967
timestamp 1677677812
transform 1 0 3492 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8989
timestamp 1677677812
transform 1 0 3484 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9102
timestamp 1677677812
transform 1 0 3452 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9103
timestamp 1677677812
transform 1 0 3468 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9141
timestamp 1677677812
transform 1 0 3452 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8080
timestamp 1677677812
transform 1 0 3452 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9142
timestamp 1677677812
transform 1 0 3484 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_8990
timestamp 1677677812
transform 1 0 3492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9104
timestamp 1677677812
transform 1 0 3548 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9143
timestamp 1677677812
transform 1 0 3540 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_8081
timestamp 1677677812
transform 1 0 3540 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_8093
timestamp 1677677812
transform 1 0 3548 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7968
timestamp 1677677812
transform 1 0 3628 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8991
timestamp 1677677812
transform 1 0 3564 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8992
timestamp 1677677812
transform 1 0 3580 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9105
timestamp 1677677812
transform 1 0 3564 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9106
timestamp 1677677812
transform 1 0 3628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9107
timestamp 1677677812
transform 1 0 3660 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8000
timestamp 1677677812
transform 1 0 3676 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8055
timestamp 1677677812
transform 1 0 3668 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7931
timestamp 1677677812
transform 1 0 3692 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7969
timestamp 1677677812
transform 1 0 3708 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_8993
timestamp 1677677812
transform 1 0 3692 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8994
timestamp 1677677812
transform 1 0 3708 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8001
timestamp 1677677812
transform 1 0 3716 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_8995
timestamp 1677677812
transform 1 0 3724 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9108
timestamp 1677677812
transform 1 0 3700 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9109
timestamp 1677677812
transform 1 0 3716 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8056
timestamp 1677677812
transform 1 0 3700 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8057
timestamp 1677677812
transform 1 0 3724 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8094
timestamp 1677677812
transform 1 0 3716 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8095
timestamp 1677677812
transform 1 0 3732 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_7932
timestamp 1677677812
transform 1 0 3788 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8996
timestamp 1677677812
transform 1 0 3772 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8997
timestamp 1677677812
transform 1 0 3788 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8002
timestamp 1677677812
transform 1 0 3796 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_9110
timestamp 1677677812
transform 1 0 3764 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9111
timestamp 1677677812
transform 1 0 3780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9112
timestamp 1677677812
transform 1 0 3788 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8058
timestamp 1677677812
transform 1 0 3788 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7970
timestamp 1677677812
transform 1 0 3884 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7933
timestamp 1677677812
transform 1 0 3916 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_8998
timestamp 1677677812
transform 1 0 3884 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_8999
timestamp 1677677812
transform 1 0 3900 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9000
timestamp 1677677812
transform 1 0 3916 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9113
timestamp 1677677812
transform 1 0 3892 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8082
timestamp 1677677812
transform 1 0 3892 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_9114
timestamp 1677677812
transform 1 0 3924 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9001
timestamp 1677677812
transform 1 0 3948 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_7934
timestamp 1677677812
transform 1 0 3972 0 1 555
box -3 -3 3 3
use M3_M2  M3_M2_7971
timestamp 1677677812
transform 1 0 3964 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9002
timestamp 1677677812
transform 1 0 3972 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8083
timestamp 1677677812
transform 1 0 3996 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7972
timestamp 1677677812
transform 1 0 4036 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9003
timestamp 1677677812
transform 1 0 4020 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9004
timestamp 1677677812
transform 1 0 4036 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9115
timestamp 1677677812
transform 1 0 4012 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9116
timestamp 1677677812
transform 1 0 4028 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8059
timestamp 1677677812
transform 1 0 4012 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9005
timestamp 1677677812
transform 1 0 4060 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9117
timestamp 1677677812
transform 1 0 4052 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8060
timestamp 1677677812
transform 1 0 4052 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8096
timestamp 1677677812
transform 1 0 4076 0 1 495
box -3 -3 3 3
use M2_M1  M2_M1_9006
timestamp 1677677812
transform 1 0 4092 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9118
timestamp 1677677812
transform 1 0 4084 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7973
timestamp 1677677812
transform 1 0 4164 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9007
timestamp 1677677812
transform 1 0 4116 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9119
timestamp 1677677812
transform 1 0 4100 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8020
timestamp 1677677812
transform 1 0 4116 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8021
timestamp 1677677812
transform 1 0 4156 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9120
timestamp 1677677812
transform 1 0 4164 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8097
timestamp 1677677812
transform 1 0 4132 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_8102
timestamp 1677677812
transform 1 0 4124 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8103
timestamp 1677677812
transform 1 0 4148 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_7974
timestamp 1677677812
transform 1 0 4260 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9008
timestamp 1677677812
transform 1 0 4244 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9009
timestamp 1677677812
transform 1 0 4260 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9121
timestamp 1677677812
transform 1 0 4252 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9122
timestamp 1677677812
transform 1 0 4268 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8084
timestamp 1677677812
transform 1 0 4268 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_7975
timestamp 1677677812
transform 1 0 4292 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9010
timestamp 1677677812
transform 1 0 4292 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9011
timestamp 1677677812
transform 1 0 4300 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8061
timestamp 1677677812
transform 1 0 4292 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_7976
timestamp 1677677812
transform 1 0 4316 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7977
timestamp 1677677812
transform 1 0 4332 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9012
timestamp 1677677812
transform 1 0 4316 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9013
timestamp 1677677812
transform 1 0 4332 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9014
timestamp 1677677812
transform 1 0 4348 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9123
timestamp 1677677812
transform 1 0 4308 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9124
timestamp 1677677812
transform 1 0 4324 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9125
timestamp 1677677812
transform 1 0 4340 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7978
timestamp 1677677812
transform 1 0 4412 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9015
timestamp 1677677812
transform 1 0 4460 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9126
timestamp 1677677812
transform 1 0 4380 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9127
timestamp 1677677812
transform 1 0 4412 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8022
timestamp 1677677812
transform 1 0 4460 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8062
timestamp 1677677812
transform 1 0 4380 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8023
timestamp 1677677812
transform 1 0 4476 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_7979
timestamp 1677677812
transform 1 0 4516 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9016
timestamp 1677677812
transform 1 0 4588 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9128
timestamp 1677677812
transform 1 0 4508 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9129
timestamp 1677677812
transform 1 0 4540 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8024
timestamp 1677677812
transform 1 0 4588 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_8063
timestamp 1677677812
transform 1 0 4548 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_9130
timestamp 1677677812
transform 1 0 4620 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9131
timestamp 1677677812
transform 1 0 4636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_7980
timestamp 1677677812
transform 1 0 4652 0 1 545
box -3 -3 3 3
use M3_M2  M3_M2_7981
timestamp 1677677812
transform 1 0 4668 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9017
timestamp 1677677812
transform 1 0 4644 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9018
timestamp 1677677812
transform 1 0 4652 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9019
timestamp 1677677812
transform 1 0 4668 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_8104
timestamp 1677677812
transform 1 0 4644 0 1 485
box -3 -3 3 3
use M3_M2  M3_M2_8003
timestamp 1677677812
transform 1 0 4676 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_7982
timestamp 1677677812
transform 1 0 4724 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_9020
timestamp 1677677812
transform 1 0 4684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9021
timestamp 1677677812
transform 1 0 4700 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_9132
timestamp 1677677812
transform 1 0 4660 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9133
timestamp 1677677812
transform 1 0 4676 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8004
timestamp 1677677812
transform 1 0 4764 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_8025
timestamp 1677677812
transform 1 0 4700 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_9134
timestamp 1677677812
transform 1 0 4724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_9135
timestamp 1677677812
transform 1 0 4788 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_8064
timestamp 1677677812
transform 1 0 4684 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_8105
timestamp 1677677812
transform 1 0 4788 0 1 485
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_84
timestamp 1677677812
transform 1 0 24 0 1 470
box -10 -3 10 3
use FILL  FILL_9814
timestamp 1677677812
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_9815
timestamp 1677677812
transform 1 0 80 0 -1 570
box -8 -3 16 105
use FILL  FILL_9816
timestamp 1677677812
transform 1 0 88 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_620
timestamp 1677677812
transform 1 0 96 0 -1 570
box -9 -3 26 105
use FILL  FILL_9817
timestamp 1677677812
transform 1 0 112 0 -1 570
box -8 -3 16 105
use FILL  FILL_9818
timestamp 1677677812
transform 1 0 120 0 -1 570
box -8 -3 16 105
use FILL  FILL_9819
timestamp 1677677812
transform 1 0 128 0 -1 570
box -8 -3 16 105
use FILL  FILL_9820
timestamp 1677677812
transform 1 0 136 0 -1 570
box -8 -3 16 105
use FILL  FILL_9821
timestamp 1677677812
transform 1 0 144 0 -1 570
box -8 -3 16 105
use FILL  FILL_9822
timestamp 1677677812
transform 1 0 152 0 -1 570
box -8 -3 16 105
use FILL  FILL_9823
timestamp 1677677812
transform 1 0 160 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_368
timestamp 1677677812
transform -1 0 208 0 -1 570
box -8 -3 46 105
use FILL  FILL_9824
timestamp 1677677812
transform 1 0 208 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_386
timestamp 1677677812
transform 1 0 216 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_528
timestamp 1677677812
transform 1 0 256 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_621
timestamp 1677677812
transform -1 0 368 0 -1 570
box -9 -3 26 105
use FILL  FILL_9825
timestamp 1677677812
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_9827
timestamp 1677677812
transform 1 0 376 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_372
timestamp 1677677812
transform -1 0 424 0 -1 570
box -8 -3 46 105
use FILL  FILL_9839
timestamp 1677677812
transform 1 0 424 0 -1 570
box -8 -3 16 105
use FILL  FILL_9840
timestamp 1677677812
transform 1 0 432 0 -1 570
box -8 -3 16 105
use FILL  FILL_9841
timestamp 1677677812
transform 1 0 440 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_387
timestamp 1677677812
transform -1 0 488 0 -1 570
box -8 -3 46 105
use OAI22X1  OAI22X1_388
timestamp 1677677812
transform -1 0 528 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_531
timestamp 1677677812
transform 1 0 528 0 -1 570
box -8 -3 104 105
use AOI22X1  AOI22X1_373
timestamp 1677677812
transform -1 0 664 0 -1 570
box -8 -3 46 105
use FILL  FILL_9842
timestamp 1677677812
transform 1 0 664 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_623
timestamp 1677677812
transform -1 0 688 0 -1 570
box -9 -3 26 105
use FILL  FILL_9843
timestamp 1677677812
transform 1 0 688 0 -1 570
box -8 -3 16 105
use FILL  FILL_9844
timestamp 1677677812
transform 1 0 696 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_110
timestamp 1677677812
transform 1 0 704 0 -1 570
box -5 -3 28 105
use FILL  FILL_9845
timestamp 1677677812
transform 1 0 728 0 -1 570
box -8 -3 16 105
use FILL  FILL_9846
timestamp 1677677812
transform 1 0 736 0 -1 570
box -8 -3 16 105
use FILL  FILL_9847
timestamp 1677677812
transform 1 0 744 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_389
timestamp 1677677812
transform 1 0 752 0 -1 570
box -8 -3 46 105
use FILL  FILL_9848
timestamp 1677677812
transform 1 0 792 0 -1 570
box -8 -3 16 105
use FILL  FILL_9850
timestamp 1677677812
transform 1 0 800 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_375
timestamp 1677677812
transform 1 0 808 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_624
timestamp 1677677812
transform 1 0 848 0 -1 570
box -9 -3 26 105
use FILL  FILL_9855
timestamp 1677677812
transform 1 0 864 0 -1 570
box -8 -3 16 105
use FILL  FILL_9856
timestamp 1677677812
transform 1 0 872 0 -1 570
box -8 -3 16 105
use FILL  FILL_9858
timestamp 1677677812
transform 1 0 880 0 -1 570
box -8 -3 16 105
use FILL  FILL_9860
timestamp 1677677812
transform 1 0 888 0 -1 570
box -8 -3 16 105
use FILL  FILL_9868
timestamp 1677677812
transform 1 0 896 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_377
timestamp 1677677812
transform -1 0 944 0 -1 570
box -8 -3 46 105
use FILL  FILL_9869
timestamp 1677677812
transform 1 0 944 0 -1 570
box -8 -3 16 105
use FILL  FILL_9870
timestamp 1677677812
transform 1 0 952 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_626
timestamp 1677677812
transform 1 0 960 0 -1 570
box -9 -3 26 105
use FILL  FILL_9871
timestamp 1677677812
transform 1 0 976 0 -1 570
box -8 -3 16 105
use FILL  FILL_9872
timestamp 1677677812
transform 1 0 984 0 -1 570
box -8 -3 16 105
use FILL  FILL_9873
timestamp 1677677812
transform 1 0 992 0 -1 570
box -8 -3 16 105
use FILL  FILL_9874
timestamp 1677677812
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_98
timestamp 1677677812
transform 1 0 1008 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_99
timestamp 1677677812
transform 1 0 1032 0 -1 570
box -8 -3 32 105
use FILL  FILL_9875
timestamp 1677677812
transform 1 0 1056 0 -1 570
box -8 -3 16 105
use FILL  FILL_9876
timestamp 1677677812
transform 1 0 1064 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_534
timestamp 1677677812
transform 1 0 1072 0 -1 570
box -8 -3 104 105
use FILL  FILL_9877
timestamp 1677677812
transform 1 0 1168 0 -1 570
box -8 -3 16 105
use FILL  FILL_9878
timestamp 1677677812
transform 1 0 1176 0 -1 570
box -8 -3 16 105
use FILL  FILL_9879
timestamp 1677677812
transform 1 0 1184 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_100
timestamp 1677677812
transform 1 0 1192 0 -1 570
box -8 -3 32 105
use FILL  FILL_9880
timestamp 1677677812
transform 1 0 1216 0 -1 570
box -8 -3 16 105
use FILL  FILL_9882
timestamp 1677677812
transform 1 0 1224 0 -1 570
box -8 -3 16 105
use FILL  FILL_9903
timestamp 1677677812
transform 1 0 1232 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8106
timestamp 1677677812
transform 1 0 1268 0 1 475
box -3 -3 3 3
use NOR2X1  NOR2X1_101
timestamp 1677677812
transform 1 0 1240 0 -1 570
box -8 -3 32 105
use FILL  FILL_9904
timestamp 1677677812
transform 1 0 1264 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_392
timestamp 1677677812
transform -1 0 1312 0 -1 570
box -8 -3 46 105
use FILL  FILL_9905
timestamp 1677677812
transform 1 0 1312 0 -1 570
box -8 -3 16 105
use FILL  FILL_9906
timestamp 1677677812
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_393
timestamp 1677677812
transform -1 0 1368 0 -1 570
box -8 -3 46 105
use FILL  FILL_9907
timestamp 1677677812
transform 1 0 1368 0 -1 570
box -8 -3 16 105
use FILL  FILL_9908
timestamp 1677677812
transform 1 0 1376 0 -1 570
box -8 -3 16 105
use FILL  FILL_9909
timestamp 1677677812
transform 1 0 1384 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_632
timestamp 1677677812
transform 1 0 1392 0 -1 570
box -9 -3 26 105
use FILL  FILL_9910
timestamp 1677677812
transform 1 0 1408 0 -1 570
box -8 -3 16 105
use FILL  FILL_9911
timestamp 1677677812
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use FILL  FILL_9912
timestamp 1677677812
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_380
timestamp 1677677812
transform 1 0 1432 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_536
timestamp 1677677812
transform -1 0 1568 0 -1 570
box -8 -3 104 105
use FILL  FILL_9913
timestamp 1677677812
transform 1 0 1568 0 -1 570
box -8 -3 16 105
use FILL  FILL_9914
timestamp 1677677812
transform 1 0 1576 0 -1 570
box -8 -3 16 105
use FILL  FILL_9915
timestamp 1677677812
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_111
timestamp 1677677812
transform -1 0 1616 0 -1 570
box -5 -3 28 105
use BUFX2  BUFX2_112
timestamp 1677677812
transform 1 0 1616 0 -1 570
box -5 -3 28 105
use FILL  FILL_9916
timestamp 1677677812
transform 1 0 1640 0 -1 570
box -8 -3 16 105
use FILL  FILL_9917
timestamp 1677677812
transform 1 0 1648 0 -1 570
box -8 -3 16 105
use FILL  FILL_9918
timestamp 1677677812
transform 1 0 1656 0 -1 570
box -8 -3 16 105
use FILL  FILL_9919
timestamp 1677677812
transform 1 0 1664 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8107
timestamp 1677677812
transform 1 0 1708 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_394
timestamp 1677677812
transform 1 0 1672 0 -1 570
box -8 -3 46 105
use FILL  FILL_9920
timestamp 1677677812
transform 1 0 1712 0 -1 570
box -8 -3 16 105
use FILL  FILL_9921
timestamp 1677677812
transform 1 0 1720 0 -1 570
box -8 -3 16 105
use FILL  FILL_9923
timestamp 1677677812
transform 1 0 1728 0 -1 570
box -8 -3 16 105
use FILL  FILL_9925
timestamp 1677677812
transform 1 0 1736 0 -1 570
box -8 -3 16 105
use FILL  FILL_9926
timestamp 1677677812
transform 1 0 1744 0 -1 570
box -8 -3 16 105
use FILL  FILL_9927
timestamp 1677677812
transform 1 0 1752 0 -1 570
box -8 -3 16 105
use FILL  FILL_9928
timestamp 1677677812
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use FILL  FILL_9929
timestamp 1677677812
transform 1 0 1768 0 -1 570
box -8 -3 16 105
use FILL  FILL_9930
timestamp 1677677812
transform 1 0 1776 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_634
timestamp 1677677812
transform 1 0 1784 0 -1 570
box -9 -3 26 105
use FILL  FILL_9931
timestamp 1677677812
transform 1 0 1800 0 -1 570
box -8 -3 16 105
use FILL  FILL_9932
timestamp 1677677812
transform 1 0 1808 0 -1 570
box -8 -3 16 105
use FILL  FILL_9933
timestamp 1677677812
transform 1 0 1816 0 -1 570
box -8 -3 16 105
use FILL  FILL_9934
timestamp 1677677812
transform 1 0 1824 0 -1 570
box -8 -3 16 105
use FILL  FILL_9935
timestamp 1677677812
transform 1 0 1832 0 -1 570
box -8 -3 16 105
use FILL  FILL_9940
timestamp 1677677812
transform 1 0 1840 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_539
timestamp 1677677812
transform -1 0 1944 0 -1 570
box -8 -3 104 105
use FILL  FILL_9941
timestamp 1677677812
transform 1 0 1944 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_636
timestamp 1677677812
transform 1 0 1952 0 -1 570
box -9 -3 26 105
use FILL  FILL_9942
timestamp 1677677812
transform 1 0 1968 0 -1 570
box -8 -3 16 105
use FILL  FILL_9943
timestamp 1677677812
transform 1 0 1976 0 -1 570
box -8 -3 16 105
use FILL  FILL_9944
timestamp 1677677812
transform 1 0 1984 0 -1 570
box -8 -3 16 105
use FILL  FILL_9945
timestamp 1677677812
transform 1 0 1992 0 -1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_383
timestamp 1677677812
transform -1 0 2040 0 -1 570
box -8 -3 46 105
use FILL  FILL_9946
timestamp 1677677812
transform 1 0 2040 0 -1 570
box -8 -3 16 105
use FILL  FILL_9947
timestamp 1677677812
transform 1 0 2048 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_637
timestamp 1677677812
transform 1 0 2056 0 -1 570
box -9 -3 26 105
use FILL  FILL_9948
timestamp 1677677812
transform 1 0 2072 0 -1 570
box -8 -3 16 105
use FILL  FILL_9952
timestamp 1677677812
transform 1 0 2080 0 -1 570
box -8 -3 16 105
use FILL  FILL_9953
timestamp 1677677812
transform 1 0 2088 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_541
timestamp 1677677812
transform -1 0 2192 0 -1 570
box -8 -3 104 105
use FILL  FILL_9954
timestamp 1677677812
transform 1 0 2192 0 -1 570
box -8 -3 16 105
use FILL  FILL_9956
timestamp 1677677812
transform 1 0 2200 0 -1 570
box -8 -3 16 105
use FILL  FILL_9958
timestamp 1677677812
transform 1 0 2208 0 -1 570
box -8 -3 16 105
use FILL  FILL_9959
timestamp 1677677812
transform 1 0 2216 0 -1 570
box -8 -3 16 105
use FILL  FILL_9960
timestamp 1677677812
transform 1 0 2224 0 -1 570
box -8 -3 16 105
use FILL  FILL_9961
timestamp 1677677812
transform 1 0 2232 0 -1 570
box -8 -3 16 105
use FILL  FILL_9962
timestamp 1677677812
transform 1 0 2240 0 -1 570
box -8 -3 16 105
use FILL  FILL_9963
timestamp 1677677812
transform 1 0 2248 0 -1 570
box -8 -3 16 105
use FILL  FILL_9964
timestamp 1677677812
transform 1 0 2256 0 -1 570
box -8 -3 16 105
use FILL  FILL_9965
timestamp 1677677812
transform 1 0 2264 0 -1 570
box -8 -3 16 105
use FILL  FILL_9966
timestamp 1677677812
transform 1 0 2272 0 -1 570
box -8 -3 16 105
use FILL  FILL_9967
timestamp 1677677812
transform 1 0 2280 0 -1 570
box -8 -3 16 105
use FILL  FILL_9968
timestamp 1677677812
transform 1 0 2288 0 -1 570
box -8 -3 16 105
use FILL  FILL_9969
timestamp 1677677812
transform 1 0 2296 0 -1 570
box -8 -3 16 105
use FILL  FILL_9970
timestamp 1677677812
transform 1 0 2304 0 -1 570
box -8 -3 16 105
use FILL  FILL_9972
timestamp 1677677812
transform 1 0 2312 0 -1 570
box -8 -3 16 105
use FILL  FILL_9974
timestamp 1677677812
transform 1 0 2320 0 -1 570
box -8 -3 16 105
use FILL  FILL_9976
timestamp 1677677812
transform 1 0 2328 0 -1 570
box -8 -3 16 105
use FILL  FILL_9978
timestamp 1677677812
transform 1 0 2336 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_40
timestamp 1677677812
transform 1 0 2344 0 -1 570
box -8 -3 32 105
use FILL  FILL_9984
timestamp 1677677812
transform 1 0 2368 0 -1 570
box -8 -3 16 105
use FILL  FILL_9985
timestamp 1677677812
transform 1 0 2376 0 -1 570
box -8 -3 16 105
use XOR2X1  XOR2X1_6
timestamp 1677677812
transform -1 0 2440 0 -1 570
box -8 -3 64 105
use FILL  FILL_9986
timestamp 1677677812
transform 1 0 2440 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_543
timestamp 1677677812
transform 1 0 2448 0 -1 570
box -8 -3 104 105
use AND2X2  AND2X2_61
timestamp 1677677812
transform -1 0 2576 0 -1 570
box -8 -3 40 105
use FILL  FILL_9997
timestamp 1677677812
transform 1 0 2576 0 -1 570
box -8 -3 16 105
use FILL  FILL_10005
timestamp 1677677812
transform 1 0 2584 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_545
timestamp 1677677812
transform -1 0 2688 0 -1 570
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_546
timestamp 1677677812
transform -1 0 2784 0 -1 570
box -8 -3 104 105
use FILL  FILL_10006
timestamp 1677677812
transform 1 0 2784 0 -1 570
box -8 -3 16 105
use FILL  FILL_10014
timestamp 1677677812
transform 1 0 2792 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_547
timestamp 1677677812
transform -1 0 2896 0 -1 570
box -8 -3 104 105
use FILL  FILL_10015
timestamp 1677677812
transform 1 0 2896 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_103
timestamp 1677677812
transform 1 0 2904 0 -1 570
box -8 -3 32 105
use FILL  FILL_10017
timestamp 1677677812
transform 1 0 2928 0 -1 570
box -8 -3 16 105
use FILL  FILL_10025
timestamp 1677677812
transform 1 0 2936 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_41
timestamp 1677677812
transform -1 0 2968 0 -1 570
box -8 -3 32 105
use FILL  FILL_10026
timestamp 1677677812
transform 1 0 2968 0 -1 570
box -8 -3 16 105
use FILL  FILL_10027
timestamp 1677677812
transform 1 0 2976 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_104
timestamp 1677677812
transform 1 0 2984 0 -1 570
box -8 -3 32 105
use FILL  FILL_10028
timestamp 1677677812
transform 1 0 3008 0 -1 570
box -8 -3 16 105
use FILL  FILL_10029
timestamp 1677677812
transform 1 0 3016 0 -1 570
box -8 -3 16 105
use FILL  FILL_10030
timestamp 1677677812
transform 1 0 3024 0 -1 570
box -8 -3 16 105
use FILL  FILL_10031
timestamp 1677677812
transform 1 0 3032 0 -1 570
box -8 -3 16 105
use NOR2X1  NOR2X1_105
timestamp 1677677812
transform 1 0 3040 0 -1 570
box -8 -3 32 105
use FILL  FILL_10036
timestamp 1677677812
transform 1 0 3064 0 -1 570
box -8 -3 16 105
use FILL  FILL_10038
timestamp 1677677812
transform 1 0 3072 0 -1 570
box -8 -3 16 105
use FILL  FILL_10054
timestamp 1677677812
transform 1 0 3080 0 -1 570
box -8 -3 16 105
use FILL  FILL_10055
timestamp 1677677812
transform 1 0 3088 0 -1 570
box -8 -3 16 105
use FILL  FILL_10056
timestamp 1677677812
transform 1 0 3096 0 -1 570
box -8 -3 16 105
use FILL  FILL_10057
timestamp 1677677812
transform 1 0 3104 0 -1 570
box -8 -3 16 105
use NAND3X1  NAND3X1_76
timestamp 1677677812
transform -1 0 3144 0 -1 570
box -8 -3 40 105
use FILL  FILL_10058
timestamp 1677677812
transform 1 0 3144 0 -1 570
box -8 -3 16 105
use FILL  FILL_10059
timestamp 1677677812
transform 1 0 3152 0 -1 570
box -8 -3 16 105
use FILL  FILL_10060
timestamp 1677677812
transform 1 0 3160 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_550
timestamp 1677677812
transform 1 0 3168 0 -1 570
box -8 -3 104 105
use FILL  FILL_10061
timestamp 1677677812
transform 1 0 3264 0 -1 570
box -8 -3 16 105
use FILL  FILL_10062
timestamp 1677677812
transform 1 0 3272 0 -1 570
box -8 -3 16 105
use FILL  FILL_10063
timestamp 1677677812
transform 1 0 3280 0 -1 570
box -8 -3 16 105
use FILL  FILL_10064
timestamp 1677677812
transform 1 0 3288 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_551
timestamp 1677677812
transform 1 0 3296 0 -1 570
box -8 -3 104 105
use FILL  FILL_10065
timestamp 1677677812
transform 1 0 3392 0 -1 570
box -8 -3 16 105
use FILL  FILL_10066
timestamp 1677677812
transform 1 0 3400 0 -1 570
box -8 -3 16 105
use FILL  FILL_10067
timestamp 1677677812
transform 1 0 3408 0 -1 570
box -8 -3 16 105
use FILL  FILL_10068
timestamp 1677677812
transform 1 0 3416 0 -1 570
box -8 -3 16 105
use FILL  FILL_10069
timestamp 1677677812
transform 1 0 3424 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_42
timestamp 1677677812
transform 1 0 3432 0 -1 570
box -8 -3 32 105
use OAI21X1  OAI21X1_176
timestamp 1677677812
transform 1 0 3456 0 -1 570
box -8 -3 34 105
use FILL  FILL_10070
timestamp 1677677812
transform 1 0 3488 0 -1 570
box -8 -3 16 105
use FILL  FILL_10071
timestamp 1677677812
transform 1 0 3496 0 -1 570
box -8 -3 16 105
use FILL  FILL_10072
timestamp 1677677812
transform 1 0 3504 0 -1 570
box -8 -3 16 105
use FILL  FILL_10073
timestamp 1677677812
transform 1 0 3512 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_44
timestamp 1677677812
transform 1 0 3520 0 -1 570
box -8 -3 32 105
use M3_M2  M3_M2_8108
timestamp 1677677812
transform 1 0 3564 0 1 475
box -3 -3 3 3
use NAND2X1  NAND2X1_45
timestamp 1677677812
transform -1 0 3568 0 -1 570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_552
timestamp 1677677812
transform 1 0 3568 0 -1 570
box -8 -3 104 105
use FILL  FILL_10083
timestamp 1677677812
transform 1 0 3664 0 -1 570
box -8 -3 16 105
use FILL  FILL_10087
timestamp 1677677812
transform 1 0 3672 0 -1 570
box -8 -3 16 105
use FILL  FILL_10088
timestamp 1677677812
transform 1 0 3680 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_8109
timestamp 1677677812
transform 1 0 3732 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_397
timestamp 1677677812
transform 1 0 3688 0 -1 570
box -8 -3 46 105
use FILL  FILL_10089
timestamp 1677677812
transform 1 0 3728 0 -1 570
box -8 -3 16 105
use FILL  FILL_10091
timestamp 1677677812
transform 1 0 3736 0 -1 570
box -8 -3 16 105
use FILL  FILL_10100
timestamp 1677677812
transform 1 0 3744 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_398
timestamp 1677677812
transform -1 0 3792 0 -1 570
box -8 -3 46 105
use FILL  FILL_10101
timestamp 1677677812
transform 1 0 3792 0 -1 570
box -8 -3 16 105
use FILL  FILL_10102
timestamp 1677677812
transform 1 0 3800 0 -1 570
box -8 -3 16 105
use FILL  FILL_10103
timestamp 1677677812
transform 1 0 3808 0 -1 570
box -8 -3 16 105
use FILL  FILL_10104
timestamp 1677677812
transform 1 0 3816 0 -1 570
box -8 -3 16 105
use FILL  FILL_10106
timestamp 1677677812
transform 1 0 3824 0 -1 570
box -8 -3 16 105
use FILL  FILL_10108
timestamp 1677677812
transform 1 0 3832 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_643
timestamp 1677677812
transform 1 0 3840 0 -1 570
box -9 -3 26 105
use FILL  FILL_10112
timestamp 1677677812
transform 1 0 3856 0 -1 570
box -8 -3 16 105
use FILL  FILL_10114
timestamp 1677677812
transform 1 0 3864 0 -1 570
box -8 -3 16 105
use FILL  FILL_10116
timestamp 1677677812
transform 1 0 3872 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_400
timestamp 1677677812
transform -1 0 3920 0 -1 570
box -8 -3 46 105
use FILL  FILL_10118
timestamp 1677677812
transform 1 0 3920 0 -1 570
box -8 -3 16 105
use FILL  FILL_10120
timestamp 1677677812
transform 1 0 3928 0 -1 570
box -8 -3 16 105
use FILL  FILL_10122
timestamp 1677677812
transform 1 0 3936 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_644
timestamp 1677677812
transform 1 0 3944 0 -1 570
box -9 -3 26 105
use FILL  FILL_10125
timestamp 1677677812
transform 1 0 3960 0 -1 570
box -8 -3 16 105
use FILL  FILL_10126
timestamp 1677677812
transform 1 0 3968 0 -1 570
box -8 -3 16 105
use FILL  FILL_10127
timestamp 1677677812
transform 1 0 3976 0 -1 570
box -8 -3 16 105
use FILL  FILL_10128
timestamp 1677677812
transform 1 0 3984 0 -1 570
box -8 -3 16 105
use FILL  FILL_10129
timestamp 1677677812
transform 1 0 3992 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_405
timestamp 1677677812
transform 1 0 4000 0 -1 570
box -8 -3 46 105
use FILL  FILL_10151
timestamp 1677677812
transform 1 0 4040 0 -1 570
box -8 -3 16 105
use FILL  FILL_10152
timestamp 1677677812
transform 1 0 4048 0 -1 570
box -8 -3 16 105
use FILL  FILL_10153
timestamp 1677677812
transform 1 0 4056 0 -1 570
box -8 -3 16 105
use FILL  FILL_10154
timestamp 1677677812
transform 1 0 4064 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_645
timestamp 1677677812
transform 1 0 4072 0 -1 570
box -9 -3 26 105
use INVX2  INVX2_646
timestamp 1677677812
transform 1 0 4088 0 -1 570
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_553
timestamp 1677677812
transform 1 0 4104 0 -1 570
box -8 -3 104 105
use FILL  FILL_10155
timestamp 1677677812
transform 1 0 4200 0 -1 570
box -8 -3 16 105
use FILL  FILL_10156
timestamp 1677677812
transform 1 0 4208 0 -1 570
box -8 -3 16 105
use FILL  FILL_10157
timestamp 1677677812
transform 1 0 4216 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_647
timestamp 1677677812
transform 1 0 4224 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_406
timestamp 1677677812
transform 1 0 4240 0 -1 570
box -8 -3 46 105
use FILL  FILL_10158
timestamp 1677677812
transform 1 0 4280 0 -1 570
box -8 -3 16 105
use FILL  FILL_10160
timestamp 1677677812
transform 1 0 4288 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_648
timestamp 1677677812
transform 1 0 4296 0 -1 570
box -9 -3 26 105
use OAI22X1  OAI22X1_407
timestamp 1677677812
transform -1 0 4352 0 -1 570
box -8 -3 46 105
use FILL  FILL_10169
timestamp 1677677812
transform 1 0 4352 0 -1 570
box -8 -3 16 105
use FILL  FILL_10171
timestamp 1677677812
transform 1 0 4360 0 -1 570
box -8 -3 16 105
use FILL  FILL_10184
timestamp 1677677812
transform 1 0 4368 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_554
timestamp 1677677812
transform -1 0 4472 0 -1 570
box -8 -3 104 105
use FILL  FILL_10185
timestamp 1677677812
transform 1 0 4472 0 -1 570
box -8 -3 16 105
use FILL  FILL_10190
timestamp 1677677812
transform 1 0 4480 0 -1 570
box -8 -3 16 105
use FILL  FILL_10191
timestamp 1677677812
transform 1 0 4488 0 -1 570
box -8 -3 16 105
use FILL  FILL_10192
timestamp 1677677812
transform 1 0 4496 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_555
timestamp 1677677812
transform -1 0 4600 0 -1 570
box -8 -3 104 105
use FILL  FILL_10193
timestamp 1677677812
transform 1 0 4600 0 -1 570
box -8 -3 16 105
use FILL  FILL_10210
timestamp 1677677812
transform 1 0 4608 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_652
timestamp 1677677812
transform -1 0 4632 0 -1 570
box -9 -3 26 105
use FILL  FILL_10211
timestamp 1677677812
transform 1 0 4632 0 -1 570
box -8 -3 16 105
use FILL  FILL_10212
timestamp 1677677812
transform 1 0 4640 0 -1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_411
timestamp 1677677812
transform 1 0 4648 0 -1 570
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_556
timestamp 1677677812
transform 1 0 4688 0 -1 570
box -8 -3 104 105
use FILL  FILL_10213
timestamp 1677677812
transform 1 0 4784 0 -1 570
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_85
timestamp 1677677812
transform 1 0 4843 0 1 470
box -10 -3 10 3
use M3_M2  M3_M2_8156
timestamp 1677677812
transform 1 0 188 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9154
timestamp 1677677812
transform 1 0 132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9155
timestamp 1677677812
transform 1 0 164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9156
timestamp 1677677812
transform 1 0 172 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9272
timestamp 1677677812
transform 1 0 84 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8236
timestamp 1677677812
transform 1 0 84 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8237
timestamp 1677677812
transform 1 0 116 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8195
timestamp 1677677812
transform 1 0 180 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9157
timestamp 1677677812
transform 1 0 188 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8196
timestamp 1677677812
transform 1 0 196 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9158
timestamp 1677677812
transform 1 0 204 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9273
timestamp 1677677812
transform 1 0 188 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9274
timestamp 1677677812
transform 1 0 196 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9275
timestamp 1677677812
transform 1 0 212 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8157
timestamp 1677677812
transform 1 0 228 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8273
timestamp 1677677812
transform 1 0 252 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8238
timestamp 1677677812
transform 1 0 268 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9159
timestamp 1677677812
transform 1 0 284 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8158
timestamp 1677677812
transform 1 0 364 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8197
timestamp 1677677812
transform 1 0 300 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8198
timestamp 1677677812
transform 1 0 324 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9160
timestamp 1677677812
transform 1 0 348 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8199
timestamp 1677677812
transform 1 0 364 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9276
timestamp 1677677812
transform 1 0 300 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8239
timestamp 1677677812
transform 1 0 300 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8274
timestamp 1677677812
transform 1 0 372 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9161
timestamp 1677677812
transform 1 0 396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9277
timestamp 1677677812
transform 1 0 388 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8136
timestamp 1677677812
transform 1 0 460 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8159
timestamp 1677677812
transform 1 0 452 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9162
timestamp 1677677812
transform 1 0 428 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8200
timestamp 1677677812
transform 1 0 436 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9163
timestamp 1677677812
transform 1 0 444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9164
timestamp 1677677812
transform 1 0 460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9278
timestamp 1677677812
transform 1 0 436 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9279
timestamp 1677677812
transform 1 0 452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9280
timestamp 1677677812
transform 1 0 460 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8160
timestamp 1677677812
transform 1 0 492 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8161
timestamp 1677677812
transform 1 0 532 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8201
timestamp 1677677812
transform 1 0 484 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9165
timestamp 1677677812
transform 1 0 492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9166
timestamp 1677677812
transform 1 0 532 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8202
timestamp 1677677812
transform 1 0 580 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9167
timestamp 1677677812
transform 1 0 588 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9281
timestamp 1677677812
transform 1 0 508 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8223
timestamp 1677677812
transform 1 0 532 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8224
timestamp 1677677812
transform 1 0 556 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8275
timestamp 1677677812
transform 1 0 508 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8137
timestamp 1677677812
transform 1 0 604 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9168
timestamp 1677677812
transform 1 0 604 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9282
timestamp 1677677812
transform 1 0 596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9169
timestamp 1677677812
transform 1 0 628 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8203
timestamp 1677677812
transform 1 0 636 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9170
timestamp 1677677812
transform 1 0 644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9283
timestamp 1677677812
transform 1 0 636 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9284
timestamp 1677677812
transform 1 0 644 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9171
timestamp 1677677812
transform 1 0 684 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8162
timestamp 1677677812
transform 1 0 732 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8204
timestamp 1677677812
transform 1 0 724 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8163
timestamp 1677677812
transform 1 0 764 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9172
timestamp 1677677812
transform 1 0 732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9173
timestamp 1677677812
transform 1 0 756 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9285
timestamp 1677677812
transform 1 0 724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9286
timestamp 1677677812
transform 1 0 732 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9287
timestamp 1677677812
transform 1 0 748 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8114
timestamp 1677677812
transform 1 0 820 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8115
timestamp 1677677812
transform 1 0 844 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8138
timestamp 1677677812
transform 1 0 796 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8164
timestamp 1677677812
transform 1 0 796 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8165
timestamp 1677677812
transform 1 0 836 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9174
timestamp 1677677812
transform 1 0 796 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8205
timestamp 1677677812
transform 1 0 804 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8206
timestamp 1677677812
transform 1 0 836 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9175
timestamp 1677677812
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9288
timestamp 1677677812
transform 1 0 876 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8240
timestamp 1677677812
transform 1 0 876 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9176
timestamp 1677677812
transform 1 0 892 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8116
timestamp 1677677812
transform 1 0 932 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9177
timestamp 1677677812
transform 1 0 964 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9289
timestamp 1677677812
transform 1 0 988 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8241
timestamp 1677677812
transform 1 0 988 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9369
timestamp 1677677812
transform 1 0 1004 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_9290
timestamp 1677677812
transform 1 0 1028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9178
timestamp 1677677812
transform 1 0 1044 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8225
timestamp 1677677812
transform 1 0 1044 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8117
timestamp 1677677812
transform 1 0 1084 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8207
timestamp 1677677812
transform 1 0 1060 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8208
timestamp 1677677812
transform 1 0 1084 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9179
timestamp 1677677812
transform 1 0 1108 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9291
timestamp 1677677812
transform 1 0 1060 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8110
timestamp 1677677812
transform 1 0 1164 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_8166
timestamp 1677677812
transform 1 0 1164 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9180
timestamp 1677677812
transform 1 0 1156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9181
timestamp 1677677812
transform 1 0 1164 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9182
timestamp 1677677812
transform 1 0 1180 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9183
timestamp 1677677812
transform 1 0 1196 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9292
timestamp 1677677812
transform 1 0 1164 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9293
timestamp 1677677812
transform 1 0 1188 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8242
timestamp 1677677812
transform 1 0 1156 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8243
timestamp 1677677812
transform 1 0 1188 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8276
timestamp 1677677812
transform 1 0 1164 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9294
timestamp 1677677812
transform 1 0 1204 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8277
timestamp 1677677812
transform 1 0 1204 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8125
timestamp 1677677812
transform 1 0 1220 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9184
timestamp 1677677812
transform 1 0 1220 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8226
timestamp 1677677812
transform 1 0 1220 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8126
timestamp 1677677812
transform 1 0 1268 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8139
timestamp 1677677812
transform 1 0 1260 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8167
timestamp 1677677812
transform 1 0 1252 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8168
timestamp 1677677812
transform 1 0 1316 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9185
timestamp 1677677812
transform 1 0 1236 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9186
timestamp 1677677812
transform 1 0 1252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9187
timestamp 1677677812
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9188
timestamp 1677677812
transform 1 0 1284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9189
timestamp 1677677812
transform 1 0 1300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9295
timestamp 1677677812
transform 1 0 1228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8209
timestamp 1677677812
transform 1 0 1308 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9296
timestamp 1677677812
transform 1 0 1260 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9297
timestamp 1677677812
transform 1 0 1268 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9298
timestamp 1677677812
transform 1 0 1292 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9299
timestamp 1677677812
transform 1 0 1308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9300
timestamp 1677677812
transform 1 0 1316 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8244
timestamp 1677677812
transform 1 0 1268 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8118
timestamp 1677677812
transform 1 0 1356 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8140
timestamp 1677677812
transform 1 0 1332 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8111
timestamp 1677677812
transform 1 0 1444 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_8141
timestamp 1677677812
transform 1 0 1436 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8169
timestamp 1677677812
transform 1 0 1340 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8170
timestamp 1677677812
transform 1 0 1380 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8171
timestamp 1677677812
transform 1 0 1404 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9190
timestamp 1677677812
transform 1 0 1340 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9191
timestamp 1677677812
transform 1 0 1380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9192
timestamp 1677677812
transform 1 0 1436 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9301
timestamp 1677677812
transform 1 0 1356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9193
timestamp 1677677812
transform 1 0 1452 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9302
timestamp 1677677812
transform 1 0 1444 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8172
timestamp 1677677812
transform 1 0 1492 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9194
timestamp 1677677812
transform 1 0 1476 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8210
timestamp 1677677812
transform 1 0 1484 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9195
timestamp 1677677812
transform 1 0 1492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9303
timestamp 1677677812
transform 1 0 1484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9304
timestamp 1677677812
transform 1 0 1492 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8112
timestamp 1677677812
transform 1 0 1596 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_8173
timestamp 1677677812
transform 1 0 1532 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8174
timestamp 1677677812
transform 1 0 1572 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9196
timestamp 1677677812
transform 1 0 1532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9197
timestamp 1677677812
transform 1 0 1540 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8211
timestamp 1677677812
transform 1 0 1548 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9198
timestamp 1677677812
transform 1 0 1572 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9305
timestamp 1677677812
transform 1 0 1620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9199
timestamp 1677677812
transform 1 0 1644 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8175
timestamp 1677677812
transform 1 0 1684 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9200
timestamp 1677677812
transform 1 0 1700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9201
timestamp 1677677812
transform 1 0 1716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9306
timestamp 1677677812
transform 1 0 1684 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9307
timestamp 1677677812
transform 1 0 1692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9308
timestamp 1677677812
transform 1 0 1708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9309
timestamp 1677677812
transform 1 0 1724 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9310
timestamp 1677677812
transform 1 0 1732 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8245
timestamp 1677677812
transform 1 0 1692 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8246
timestamp 1677677812
transform 1 0 1732 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8278
timestamp 1677677812
transform 1 0 1724 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8113
timestamp 1677677812
transform 1 0 1804 0 1 465
box -3 -3 3 3
use M3_M2  M3_M2_8176
timestamp 1677677812
transform 1 0 1788 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8177
timestamp 1677677812
transform 1 0 1804 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9202
timestamp 1677677812
transform 1 0 1764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9203
timestamp 1677677812
transform 1 0 1772 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9204
timestamp 1677677812
transform 1 0 1788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9205
timestamp 1677677812
transform 1 0 1804 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9206
timestamp 1677677812
transform 1 0 1812 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9207
timestamp 1677677812
transform 1 0 1844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9311
timestamp 1677677812
transform 1 0 1796 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9312
timestamp 1677677812
transform 1 0 1804 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9313
timestamp 1677677812
transform 1 0 1892 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9314
timestamp 1677677812
transform 1 0 1908 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8142
timestamp 1677677812
transform 1 0 1940 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8143
timestamp 1677677812
transform 1 0 1972 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9208
timestamp 1677677812
transform 1 0 1940 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9209
timestamp 1677677812
transform 1 0 1956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9210
timestamp 1677677812
transform 1 0 1980 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8127
timestamp 1677677812
transform 1 0 1996 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8128
timestamp 1677677812
transform 1 0 2020 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8129
timestamp 1677677812
transform 1 0 2036 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8144
timestamp 1677677812
transform 1 0 2028 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8178
timestamp 1677677812
transform 1 0 1996 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8179
timestamp 1677677812
transform 1 0 2012 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8180
timestamp 1677677812
transform 1 0 2036 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9211
timestamp 1677677812
transform 1 0 1996 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9212
timestamp 1677677812
transform 1 0 2012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9213
timestamp 1677677812
transform 1 0 2028 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9315
timestamp 1677677812
transform 1 0 1996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9316
timestamp 1677677812
transform 1 0 2004 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9317
timestamp 1677677812
transform 1 0 2028 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9318
timestamp 1677677812
transform 1 0 2036 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8279
timestamp 1677677812
transform 1 0 2028 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8181
timestamp 1677677812
transform 1 0 2092 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8182
timestamp 1677677812
transform 1 0 2132 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9214
timestamp 1677677812
transform 1 0 2092 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9215
timestamp 1677677812
transform 1 0 2100 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9216
timestamp 1677677812
transform 1 0 2132 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9319
timestamp 1677677812
transform 1 0 2180 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8247
timestamp 1677677812
transform 1 0 2140 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8248
timestamp 1677677812
transform 1 0 2180 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8280
timestamp 1677677812
transform 1 0 2100 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9217
timestamp 1677677812
transform 1 0 2244 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9218
timestamp 1677677812
transform 1 0 2300 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9320
timestamp 1677677812
transform 1 0 2220 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8130
timestamp 1677677812
transform 1 0 2332 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9321
timestamp 1677677812
transform 1 0 2316 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9370
timestamp 1677677812
transform 1 0 2308 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_8249
timestamp 1677677812
transform 1 0 2316 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8281
timestamp 1677677812
transform 1 0 2308 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9322
timestamp 1677677812
transform 1 0 2340 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8282
timestamp 1677677812
transform 1 0 2340 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9219
timestamp 1677677812
transform 1 0 2356 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9371
timestamp 1677677812
transform 1 0 2356 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_9220
timestamp 1677677812
transform 1 0 2372 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9323
timestamp 1677677812
transform 1 0 2380 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8250
timestamp 1677677812
transform 1 0 2372 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8212
timestamp 1677677812
transform 1 0 2460 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9221
timestamp 1677677812
transform 1 0 2476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9222
timestamp 1677677812
transform 1 0 2500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9223
timestamp 1677677812
transform 1 0 2540 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9324
timestamp 1677677812
transform 1 0 2484 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9325
timestamp 1677677812
transform 1 0 2580 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8251
timestamp 1677677812
transform 1 0 2580 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8283
timestamp 1677677812
transform 1 0 2580 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8213
timestamp 1677677812
transform 1 0 2620 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8131
timestamp 1677677812
transform 1 0 2804 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9224
timestamp 1677677812
transform 1 0 2644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9225
timestamp 1677677812
transform 1 0 2700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9226
timestamp 1677677812
transform 1 0 2708 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9227
timestamp 1677677812
transform 1 0 2764 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9326
timestamp 1677677812
transform 1 0 2620 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8284
timestamp 1677677812
transform 1 0 2644 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8214
timestamp 1677677812
transform 1 0 2788 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8227
timestamp 1677677812
transform 1 0 2764 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9327
timestamp 1677677812
transform 1 0 2788 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9328
timestamp 1677677812
transform 1 0 2804 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8252
timestamp 1677677812
transform 1 0 2748 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8253
timestamp 1677677812
transform 1 0 2804 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8145
timestamp 1677677812
transform 1 0 2836 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8132
timestamp 1677677812
transform 1 0 2852 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8146
timestamp 1677677812
transform 1 0 2924 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8183
timestamp 1677677812
transform 1 0 2900 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9228
timestamp 1677677812
transform 1 0 2836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9229
timestamp 1677677812
transform 1 0 2844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9230
timestamp 1677677812
transform 1 0 2900 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8215
timestamp 1677677812
transform 1 0 2924 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9329
timestamp 1677677812
transform 1 0 2924 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9146
timestamp 1677677812
transform 1 0 2940 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8228
timestamp 1677677812
transform 1 0 2940 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8229
timestamp 1677677812
transform 1 0 2964 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8184
timestamp 1677677812
transform 1 0 2996 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9330
timestamp 1677677812
transform 1 0 2988 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9331
timestamp 1677677812
transform 1 0 2996 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9147
timestamp 1677677812
transform 1 0 3020 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9372
timestamp 1677677812
transform 1 0 3012 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_8147
timestamp 1677677812
transform 1 0 3044 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9145
timestamp 1677677812
transform 1 0 3052 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_9148
timestamp 1677677812
transform 1 0 3052 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9231
timestamp 1677677812
transform 1 0 3068 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8185
timestamp 1677677812
transform 1 0 3084 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9332
timestamp 1677677812
transform 1 0 3084 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8148
timestamp 1677677812
transform 1 0 3100 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8186
timestamp 1677677812
transform 1 0 3140 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9232
timestamp 1677677812
transform 1 0 3140 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9333
timestamp 1677677812
transform 1 0 3100 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9334
timestamp 1677677812
transform 1 0 3116 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8187
timestamp 1677677812
transform 1 0 3212 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9233
timestamp 1677677812
transform 1 0 3212 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8149
timestamp 1677677812
transform 1 0 3260 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9234
timestamp 1677677812
transform 1 0 3260 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9335
timestamp 1677677812
transform 1 0 3228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8188
timestamp 1677677812
transform 1 0 3316 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9336
timestamp 1677677812
transform 1 0 3316 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8216
timestamp 1677677812
transform 1 0 3332 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9235
timestamp 1677677812
transform 1 0 3340 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8254
timestamp 1677677812
transform 1 0 3340 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9149
timestamp 1677677812
transform 1 0 3364 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8217
timestamp 1677677812
transform 1 0 3364 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9337
timestamp 1677677812
transform 1 0 3364 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8255
timestamp 1677677812
transform 1 0 3364 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9236
timestamp 1677677812
transform 1 0 3380 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8230
timestamp 1677677812
transform 1 0 3380 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8133
timestamp 1677677812
transform 1 0 3396 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9150
timestamp 1677677812
transform 1 0 3412 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9237
timestamp 1677677812
transform 1 0 3396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9238
timestamp 1677677812
transform 1 0 3404 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8218
timestamp 1677677812
transform 1 0 3412 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9338
timestamp 1677677812
transform 1 0 3420 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8219
timestamp 1677677812
transform 1 0 3452 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8231
timestamp 1677677812
transform 1 0 3444 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8119
timestamp 1677677812
transform 1 0 3484 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8150
timestamp 1677677812
transform 1 0 3476 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9151
timestamp 1677677812
transform 1 0 3476 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_8151
timestamp 1677677812
transform 1 0 3508 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9152
timestamp 1677677812
transform 1 0 3508 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9239
timestamp 1677677812
transform 1 0 3484 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9240
timestamp 1677677812
transform 1 0 3492 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9339
timestamp 1677677812
transform 1 0 3484 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8256
timestamp 1677677812
transform 1 0 3460 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8257
timestamp 1677677812
transform 1 0 3484 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8152
timestamp 1677677812
transform 1 0 3548 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9153
timestamp 1677677812
transform 1 0 3548 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_9241
timestamp 1677677812
transform 1 0 3524 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9242
timestamp 1677677812
transform 1 0 3532 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9340
timestamp 1677677812
transform 1 0 3516 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8258
timestamp 1677677812
transform 1 0 3516 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9243
timestamp 1677677812
transform 1 0 3612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9341
timestamp 1677677812
transform 1 0 3548 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9342
timestamp 1677677812
transform 1 0 3564 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8259
timestamp 1677677812
transform 1 0 3612 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8285
timestamp 1677677812
transform 1 0 3548 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8286
timestamp 1677677812
transform 1 0 3628 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_9343
timestamp 1677677812
transform 1 0 3652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9244
timestamp 1677677812
transform 1 0 3684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9245
timestamp 1677677812
transform 1 0 3700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9246
timestamp 1677677812
transform 1 0 3716 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9344
timestamp 1677677812
transform 1 0 3692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9345
timestamp 1677677812
transform 1 0 3708 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9346
timestamp 1677677812
transform 1 0 3724 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8287
timestamp 1677677812
transform 1 0 3684 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8260
timestamp 1677677812
transform 1 0 3708 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8261
timestamp 1677677812
transform 1 0 3732 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8288
timestamp 1677677812
transform 1 0 3724 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8134
timestamp 1677677812
transform 1 0 3892 0 1 445
box -3 -3 3 3
use M3_M2  M3_M2_8135
timestamp 1677677812
transform 1 0 3908 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_9247
timestamp 1677677812
transform 1 0 3788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9248
timestamp 1677677812
transform 1 0 3844 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9249
timestamp 1677677812
transform 1 0 3860 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9250
timestamp 1677677812
transform 1 0 3900 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9251
timestamp 1677677812
transform 1 0 3956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9347
timestamp 1677677812
transform 1 0 3764 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9348
timestamp 1677677812
transform 1 0 3852 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9349
timestamp 1677677812
transform 1 0 3876 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9252
timestamp 1677677812
transform 1 0 4020 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9253
timestamp 1677677812
transform 1 0 4060 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9350
timestamp 1677677812
transform 1 0 3980 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8232
timestamp 1677677812
transform 1 0 4028 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8262
timestamp 1677677812
transform 1 0 4028 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_9254
timestamp 1677677812
transform 1 0 4076 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9255
timestamp 1677677812
transform 1 0 4108 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8289
timestamp 1677677812
transform 1 0 4068 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8233
timestamp 1677677812
transform 1 0 4084 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_9351
timestamp 1677677812
transform 1 0 4156 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8263
timestamp 1677677812
transform 1 0 4156 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8189
timestamp 1677677812
transform 1 0 4172 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8190
timestamp 1677677812
transform 1 0 4196 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8120
timestamp 1677677812
transform 1 0 4244 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8220
timestamp 1677677812
transform 1 0 4228 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_8221
timestamp 1677677812
transform 1 0 4252 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9256
timestamp 1677677812
transform 1 0 4276 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9257
timestamp 1677677812
transform 1 0 4308 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9258
timestamp 1677677812
transform 1 0 4316 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9352
timestamp 1677677812
transform 1 0 4228 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8264
timestamp 1677677812
transform 1 0 4228 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8265
timestamp 1677677812
transform 1 0 4276 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8121
timestamp 1677677812
transform 1 0 4332 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9353
timestamp 1677677812
transform 1 0 4332 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8290
timestamp 1677677812
transform 1 0 4332 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8122
timestamp 1677677812
transform 1 0 4348 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9259
timestamp 1677677812
transform 1 0 4364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9260
timestamp 1677677812
transform 1 0 4380 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9354
timestamp 1677677812
transform 1 0 4356 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9355
timestamp 1677677812
transform 1 0 4372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9356
timestamp 1677677812
transform 1 0 4380 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8266
timestamp 1677677812
transform 1 0 4356 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8291
timestamp 1677677812
transform 1 0 4380 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8292
timestamp 1677677812
transform 1 0 4396 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8123
timestamp 1677677812
transform 1 0 4452 0 1 455
box -3 -3 3 3
use M2_M1  M2_M1_9261
timestamp 1677677812
transform 1 0 4428 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8234
timestamp 1677677812
transform 1 0 4428 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8153
timestamp 1677677812
transform 1 0 4460 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9262
timestamp 1677677812
transform 1 0 4460 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9357
timestamp 1677677812
transform 1 0 4436 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9358
timestamp 1677677812
transform 1 0 4452 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8267
timestamp 1677677812
transform 1 0 4436 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8293
timestamp 1677677812
transform 1 0 4452 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8124
timestamp 1677677812
transform 1 0 4516 0 1 455
box -3 -3 3 3
use M3_M2  M3_M2_8154
timestamp 1677677812
transform 1 0 4524 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_8155
timestamp 1677677812
transform 1 0 4564 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_9263
timestamp 1677677812
transform 1 0 4500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9264
timestamp 1677677812
transform 1 0 4556 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9265
timestamp 1677677812
transform 1 0 4564 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9359
timestamp 1677677812
transform 1 0 4476 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8268
timestamp 1677677812
transform 1 0 4500 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8269
timestamp 1677677812
transform 1 0 4564 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8294
timestamp 1677677812
transform 1 0 4476 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8191
timestamp 1677677812
transform 1 0 4588 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9266
timestamp 1677677812
transform 1 0 4588 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_8222
timestamp 1677677812
transform 1 0 4612 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_9267
timestamp 1677677812
transform 1 0 4628 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9268
timestamp 1677677812
transform 1 0 4636 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9360
timestamp 1677677812
transform 1 0 4572 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9361
timestamp 1677677812
transform 1 0 4580 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9362
timestamp 1677677812
transform 1 0 4596 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9363
timestamp 1677677812
transform 1 0 4612 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8270
timestamp 1677677812
transform 1 0 4604 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8295
timestamp 1677677812
transform 1 0 4580 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_8192
timestamp 1677677812
transform 1 0 4684 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9269
timestamp 1677677812
transform 1 0 4684 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9364
timestamp 1677677812
transform 1 0 4652 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9365
timestamp 1677677812
transform 1 0 4660 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9366
timestamp 1677677812
transform 1 0 4676 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8235
timestamp 1677677812
transform 1 0 4684 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_8193
timestamp 1677677812
transform 1 0 4732 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_8194
timestamp 1677677812
transform 1 0 4748 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_9270
timestamp 1677677812
transform 1 0 4732 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9271
timestamp 1677677812
transform 1 0 4788 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_9367
timestamp 1677677812
transform 1 0 4692 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_9368
timestamp 1677677812
transform 1 0 4708 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_8271
timestamp 1677677812
transform 1 0 4676 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8272
timestamp 1677677812
transform 1 0 4732 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_8296
timestamp 1677677812
transform 1 0 4724 0 1 385
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_86
timestamp 1677677812
transform 1 0 48 0 1 370
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_557
timestamp 1677677812
transform 1 0 72 0 1 370
box -8 -3 104 105
use INVX2  INVX2_653
timestamp 1677677812
transform -1 0 184 0 1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_384
timestamp 1677677812
transform -1 0 224 0 1 370
box -8 -3 46 105
use FILL  FILL_10214
timestamp 1677677812
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_10223
timestamp 1677677812
transform 1 0 232 0 1 370
box -8 -3 16 105
use FILL  FILL_10225
timestamp 1677677812
transform 1 0 240 0 1 370
box -8 -3 16 105
use FILL  FILL_10226
timestamp 1677677812
transform 1 0 248 0 1 370
box -8 -3 16 105
use FILL  FILL_10227
timestamp 1677677812
transform 1 0 256 0 1 370
box -8 -3 16 105
use FILL  FILL_10228
timestamp 1677677812
transform 1 0 264 0 1 370
box -8 -3 16 105
use FILL  FILL_10229
timestamp 1677677812
transform 1 0 272 0 1 370
box -8 -3 16 105
use FILL  FILL_10230
timestamp 1677677812
transform 1 0 280 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_559
timestamp 1677677812
transform 1 0 288 0 1 370
box -8 -3 104 105
use FILL  FILL_10231
timestamp 1677677812
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_10232
timestamp 1677677812
transform 1 0 392 0 1 370
box -8 -3 16 105
use FILL  FILL_10233
timestamp 1677677812
transform 1 0 400 0 1 370
box -8 -3 16 105
use FILL  FILL_10234
timestamp 1677677812
transform 1 0 408 0 1 370
box -8 -3 16 105
use FILL  FILL_10235
timestamp 1677677812
transform 1 0 416 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_385
timestamp 1677677812
transform -1 0 464 0 1 370
box -8 -3 46 105
use FILL  FILL_10236
timestamp 1677677812
transform 1 0 464 0 1 370
box -8 -3 16 105
use FILL  FILL_10237
timestamp 1677677812
transform 1 0 472 0 1 370
box -8 -3 16 105
use INVX2  INVX2_654
timestamp 1677677812
transform 1 0 480 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_560
timestamp 1677677812
transform 1 0 496 0 1 370
box -8 -3 104 105
use FILL  FILL_10238
timestamp 1677677812
transform 1 0 592 0 1 370
box -8 -3 16 105
use FILL  FILL_10251
timestamp 1677677812
transform 1 0 600 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_386
timestamp 1677677812
transform 1 0 608 0 1 370
box -8 -3 46 105
use FILL  FILL_10252
timestamp 1677677812
transform 1 0 648 0 1 370
box -8 -3 16 105
use FILL  FILL_10253
timestamp 1677677812
transform 1 0 656 0 1 370
box -8 -3 16 105
use INVX2  INVX2_657
timestamp 1677677812
transform 1 0 664 0 1 370
box -9 -3 26 105
use FILL  FILL_10254
timestamp 1677677812
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_10255
timestamp 1677677812
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_10256
timestamp 1677677812
transform 1 0 696 0 1 370
box -8 -3 16 105
use FILL  FILL_10257
timestamp 1677677812
transform 1 0 704 0 1 370
box -8 -3 16 105
use FILL  FILL_10258
timestamp 1677677812
transform 1 0 712 0 1 370
box -8 -3 16 105
use FILL  FILL_10259
timestamp 1677677812
transform 1 0 720 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_413
timestamp 1677677812
transform 1 0 728 0 1 370
box -8 -3 46 105
use FILL  FILL_10260
timestamp 1677677812
transform 1 0 768 0 1 370
box -8 -3 16 105
use FILL  FILL_10261
timestamp 1677677812
transform 1 0 776 0 1 370
box -8 -3 16 105
use FILL  FILL_10262
timestamp 1677677812
transform 1 0 784 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_563
timestamp 1677677812
transform -1 0 888 0 1 370
box -8 -3 104 105
use FILL  FILL_10263
timestamp 1677677812
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_10264
timestamp 1677677812
transform 1 0 896 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_564
timestamp 1677677812
transform -1 0 1000 0 1 370
box -8 -3 104 105
use FILL  FILL_10265
timestamp 1677677812
transform 1 0 1000 0 1 370
box -8 -3 16 105
use FILL  FILL_10282
timestamp 1677677812
transform 1 0 1008 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_112
timestamp 1677677812
transform 1 0 1016 0 1 370
box -8 -3 32 105
use FILL  FILL_10284
timestamp 1677677812
transform 1 0 1040 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_566
timestamp 1677677812
transform 1 0 1048 0 1 370
box -8 -3 104 105
use FILL  FILL_10286
timestamp 1677677812
transform 1 0 1144 0 1 370
box -8 -3 16 105
use FILL  FILL_10296
timestamp 1677677812
transform 1 0 1152 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_389
timestamp 1677677812
transform 1 0 1160 0 1 370
box -8 -3 46 105
use FILL  FILL_10298
timestamp 1677677812
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_10299
timestamp 1677677812
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_10300
timestamp 1677677812
transform 1 0 1216 0 1 370
box -8 -3 16 105
use FILL  FILL_10301
timestamp 1677677812
transform 1 0 1224 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_390
timestamp 1677677812
transform 1 0 1232 0 1 370
box -8 -3 46 105
use OAI22X1  OAI22X1_415
timestamp 1677677812
transform -1 0 1312 0 1 370
box -8 -3 46 105
use FILL  FILL_10302
timestamp 1677677812
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_10313
timestamp 1677677812
transform 1 0 1320 0 1 370
box -8 -3 16 105
use INVX2  INVX2_661
timestamp 1677677812
transform 1 0 1328 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_567
timestamp 1677677812
transform 1 0 1344 0 1 370
box -8 -3 104 105
use FILL  FILL_10315
timestamp 1677677812
transform 1 0 1440 0 1 370
box -8 -3 16 105
use FILL  FILL_10316
timestamp 1677677812
transform 1 0 1448 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_391
timestamp 1677677812
transform 1 0 1456 0 1 370
box -8 -3 46 105
use FILL  FILL_10317
timestamp 1677677812
transform 1 0 1496 0 1 370
box -8 -3 16 105
use FILL  FILL_10318
timestamp 1677677812
transform 1 0 1504 0 1 370
box -8 -3 16 105
use FILL  FILL_10319
timestamp 1677677812
transform 1 0 1512 0 1 370
box -8 -3 16 105
use INVX2  INVX2_662
timestamp 1677677812
transform 1 0 1520 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_568
timestamp 1677677812
transform -1 0 1632 0 1 370
box -8 -3 104 105
use FILL  FILL_10320
timestamp 1677677812
transform 1 0 1632 0 1 370
box -8 -3 16 105
use INVX2  INVX2_663
timestamp 1677677812
transform -1 0 1656 0 1 370
box -9 -3 26 105
use FILL  FILL_10321
timestamp 1677677812
transform 1 0 1656 0 1 370
box -8 -3 16 105
use FILL  FILL_10322
timestamp 1677677812
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_10323
timestamp 1677677812
transform 1 0 1672 0 1 370
box -8 -3 16 105
use FILL  FILL_10324
timestamp 1677677812
transform 1 0 1680 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_418
timestamp 1677677812
transform -1 0 1728 0 1 370
box -8 -3 46 105
use FILL  FILL_10325
timestamp 1677677812
transform 1 0 1728 0 1 370
box -8 -3 16 105
use FILL  FILL_10326
timestamp 1677677812
transform 1 0 1736 0 1 370
box -8 -3 16 105
use FILL  FILL_10327
timestamp 1677677812
transform 1 0 1744 0 1 370
box -8 -3 16 105
use FILL  FILL_10328
timestamp 1677677812
transform 1 0 1752 0 1 370
box -8 -3 16 105
use FILL  FILL_10329
timestamp 1677677812
transform 1 0 1760 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_392
timestamp 1677677812
transform -1 0 1808 0 1 370
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_569
timestamp 1677677812
transform -1 0 1904 0 1 370
box -8 -3 104 105
use FILL  FILL_10330
timestamp 1677677812
transform 1 0 1904 0 1 370
box -8 -3 16 105
use FILL  FILL_10331
timestamp 1677677812
transform 1 0 1912 0 1 370
box -8 -3 16 105
use FILL  FILL_10332
timestamp 1677677812
transform 1 0 1920 0 1 370
box -8 -3 16 105
use FILL  FILL_10333
timestamp 1677677812
transform 1 0 1928 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_393
timestamp 1677677812
transform -1 0 1976 0 1 370
box -8 -3 46 105
use FILL  FILL_10334
timestamp 1677677812
transform 1 0 1976 0 1 370
box -8 -3 16 105
use FILL  FILL_10360
timestamp 1677677812
transform 1 0 1984 0 1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_395
timestamp 1677677812
transform 1 0 1992 0 1 370
box -8 -3 46 105
use FILL  FILL_10362
timestamp 1677677812
transform 1 0 2032 0 1 370
box -8 -3 16 105
use FILL  FILL_10363
timestamp 1677677812
transform 1 0 2040 0 1 370
box -8 -3 16 105
use FILL  FILL_10364
timestamp 1677677812
transform 1 0 2048 0 1 370
box -8 -3 16 105
use INVX2  INVX2_667
timestamp 1677677812
transform 1 0 2056 0 1 370
box -9 -3 26 105
use FILL  FILL_10368
timestamp 1677677812
transform 1 0 2072 0 1 370
box -8 -3 16 105
use FILL  FILL_10372
timestamp 1677677812
transform 1 0 2080 0 1 370
box -8 -3 16 105
use FILL  FILL_10374
timestamp 1677677812
transform 1 0 2088 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_573
timestamp 1677677812
transform -1 0 2192 0 1 370
box -8 -3 104 105
use FILL  FILL_10375
timestamp 1677677812
transform 1 0 2192 0 1 370
box -8 -3 16 105
use FILL  FILL_10376
timestamp 1677677812
transform 1 0 2200 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8297
timestamp 1677677812
transform 1 0 2252 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_574
timestamp 1677677812
transform 1 0 2208 0 1 370
box -8 -3 104 105
use M3_M2  M3_M2_8298
timestamp 1677677812
transform 1 0 2316 0 1 375
box -3 -3 3 3
use OR2X1  OR2X1_1
timestamp 1677677812
transform 1 0 2304 0 1 370
box -8 -3 40 105
use FILL  FILL_10377
timestamp 1677677812
transform 1 0 2336 0 1 370
box -8 -3 16 105
use FILL  FILL_10384
timestamp 1677677812
transform 1 0 2344 0 1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_114
timestamp 1677677812
transform 1 0 2352 0 1 370
box -8 -3 32 105
use FILL  FILL_10385
timestamp 1677677812
transform 1 0 2376 0 1 370
box -8 -3 16 105
use FILL  FILL_10386
timestamp 1677677812
transform 1 0 2384 0 1 370
box -8 -3 16 105
use FILL  FILL_10387
timestamp 1677677812
transform 1 0 2392 0 1 370
box -8 -3 16 105
use FILL  FILL_10388
timestamp 1677677812
transform 1 0 2400 0 1 370
box -8 -3 16 105
use FILL  FILL_10389
timestamp 1677677812
transform 1 0 2408 0 1 370
box -8 -3 16 105
use FILL  FILL_10390
timestamp 1677677812
transform 1 0 2416 0 1 370
box -8 -3 16 105
use FILL  FILL_10391
timestamp 1677677812
transform 1 0 2424 0 1 370
box -8 -3 16 105
use FILL  FILL_10392
timestamp 1677677812
transform 1 0 2432 0 1 370
box -8 -3 16 105
use FILL  FILL_10393
timestamp 1677677812
transform 1 0 2440 0 1 370
box -8 -3 16 105
use FILL  FILL_10394
timestamp 1677677812
transform 1 0 2448 0 1 370
box -8 -3 16 105
use FILL  FILL_10397
timestamp 1677677812
transform 1 0 2456 0 1 370
box -8 -3 16 105
use FILL  FILL_10399
timestamp 1677677812
transform 1 0 2464 0 1 370
box -8 -3 16 105
use FILL  FILL_10401
timestamp 1677677812
transform 1 0 2472 0 1 370
box -8 -3 16 105
use INVX2  INVX2_669
timestamp 1677677812
transform 1 0 2480 0 1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_578
timestamp 1677677812
transform -1 0 2592 0 1 370
box -8 -3 104 105
use FILL  FILL_10403
timestamp 1677677812
transform 1 0 2592 0 1 370
box -8 -3 16 105
use FILL  FILL_10411
timestamp 1677677812
transform 1 0 2600 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_579
timestamp 1677677812
transform 1 0 2608 0 1 370
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_580
timestamp 1677677812
transform -1 0 2800 0 1 370
box -8 -3 104 105
use BUFX2  BUFX2_114
timestamp 1677677812
transform -1 0 2824 0 1 370
box -5 -3 28 105
use FILL  FILL_10412
timestamp 1677677812
transform 1 0 2824 0 1 370
box -8 -3 16 105
use FILL  FILL_10413
timestamp 1677677812
transform 1 0 2832 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8299
timestamp 1677677812
transform 1 0 2940 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_581
timestamp 1677677812
transform -1 0 2936 0 1 370
box -8 -3 104 105
use FILL  FILL_10414
timestamp 1677677812
transform 1 0 2936 0 1 370
box -8 -3 16 105
use FILL  FILL_10415
timestamp 1677677812
transform 1 0 2944 0 1 370
box -8 -3 16 105
use FILL  FILL_10416
timestamp 1677677812
transform 1 0 2952 0 1 370
box -8 -3 16 105
use FILL  FILL_10417
timestamp 1677677812
transform 1 0 2960 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_46
timestamp 1677677812
transform -1 0 2992 0 1 370
box -8 -3 32 105
use NOR2X1  NOR2X1_115
timestamp 1677677812
transform -1 0 3016 0 1 370
box -8 -3 32 105
use FILL  FILL_10418
timestamp 1677677812
transform 1 0 3016 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_78
timestamp 1677677812
transform -1 0 3056 0 1 370
box -8 -3 40 105
use INVX2  INVX2_670
timestamp 1677677812
transform -1 0 3072 0 1 370
box -9 -3 26 105
use FILL  FILL_10419
timestamp 1677677812
transform 1 0 3072 0 1 370
box -8 -3 16 105
use FILL  FILL_10435
timestamp 1677677812
transform 1 0 3080 0 1 370
box -8 -3 16 105
use INVX2  INVX2_673
timestamp 1677677812
transform -1 0 3104 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_8300
timestamp 1677677812
transform 1 0 3116 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8301
timestamp 1677677812
transform 1 0 3172 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_584
timestamp 1677677812
transform 1 0 3104 0 1 370
box -8 -3 104 105
use FILL  FILL_10436
timestamp 1677677812
transform 1 0 3200 0 1 370
box -8 -3 16 105
use FILL  FILL_10437
timestamp 1677677812
transform 1 0 3208 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8302
timestamp 1677677812
transform 1 0 3228 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_585
timestamp 1677677812
transform 1 0 3216 0 1 370
box -8 -3 104 105
use FILL  FILL_10438
timestamp 1677677812
transform 1 0 3312 0 1 370
box -8 -3 16 105
use FILL  FILL_10447
timestamp 1677677812
transform 1 0 3320 0 1 370
box -8 -3 16 105
use FILL  FILL_10449
timestamp 1677677812
transform 1 0 3328 0 1 370
box -8 -3 16 105
use FILL  FILL_10451
timestamp 1677677812
transform 1 0 3336 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_48
timestamp 1677677812
transform 1 0 3344 0 1 370
box -8 -3 32 105
use FILL  FILL_10452
timestamp 1677677812
transform 1 0 3368 0 1 370
box -8 -3 16 105
use FILL  FILL_10453
timestamp 1677677812
transform 1 0 3376 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_49
timestamp 1677677812
transform 1 0 3384 0 1 370
box -8 -3 32 105
use FILL  FILL_10454
timestamp 1677677812
transform 1 0 3408 0 1 370
box -8 -3 16 105
use FILL  FILL_10455
timestamp 1677677812
transform 1 0 3416 0 1 370
box -8 -3 16 105
use FILL  FILL_10456
timestamp 1677677812
transform 1 0 3424 0 1 370
box -8 -3 16 105
use FILL  FILL_10459
timestamp 1677677812
transform 1 0 3432 0 1 370
box -8 -3 16 105
use FILL  FILL_10461
timestamp 1677677812
transform 1 0 3440 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_178
timestamp 1677677812
transform 1 0 3448 0 1 370
box -8 -3 34 105
use M3_M2  M3_M2_8303
timestamp 1677677812
transform 1 0 3516 0 1 375
box -3 -3 3 3
use OAI21X1  OAI21X1_179
timestamp 1677677812
transform 1 0 3480 0 1 370
box -8 -3 34 105
use FILL  FILL_10463
timestamp 1677677812
transform 1 0 3512 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_180
timestamp 1677677812
transform 1 0 3520 0 1 370
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_587
timestamp 1677677812
transform 1 0 3552 0 1 370
box -8 -3 104 105
use FILL  FILL_10464
timestamp 1677677812
transform 1 0 3648 0 1 370
box -8 -3 16 105
use FILL  FILL_10465
timestamp 1677677812
transform 1 0 3656 0 1 370
box -8 -3 16 105
use FILL  FILL_10466
timestamp 1677677812
transform 1 0 3664 0 1 370
box -8 -3 16 105
use FILL  FILL_10467
timestamp 1677677812
transform 1 0 3672 0 1 370
box -8 -3 16 105
use FILL  FILL_10479
timestamp 1677677812
transform 1 0 3680 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_422
timestamp 1677677812
transform 1 0 3688 0 1 370
box -8 -3 46 105
use FILL  FILL_10481
timestamp 1677677812
transform 1 0 3728 0 1 370
box -8 -3 16 105
use FILL  FILL_10486
timestamp 1677677812
transform 1 0 3736 0 1 370
box -8 -3 16 105
use FILL  FILL_10488
timestamp 1677677812
transform 1 0 3744 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_588
timestamp 1677677812
transform 1 0 3752 0 1 370
box -8 -3 104 105
use INVX2  INVX2_680
timestamp 1677677812
transform 1 0 3848 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_8304
timestamp 1677677812
transform 1 0 3924 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_589
timestamp 1677677812
transform 1 0 3864 0 1 370
box -8 -3 104 105
use FILL  FILL_10490
timestamp 1677677812
transform 1 0 3960 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_590
timestamp 1677677812
transform 1 0 3968 0 1 370
box -8 -3 104 105
use FILL  FILL_10491
timestamp 1677677812
transform 1 0 4064 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_591
timestamp 1677677812
transform -1 0 4168 0 1 370
box -8 -3 104 105
use FILL  FILL_10492
timestamp 1677677812
transform 1 0 4168 0 1 370
box -8 -3 16 105
use FILL  FILL_10493
timestamp 1677677812
transform 1 0 4176 0 1 370
box -8 -3 16 105
use FILL  FILL_10494
timestamp 1677677812
transform 1 0 4184 0 1 370
box -8 -3 16 105
use FILL  FILL_10513
timestamp 1677677812
transform 1 0 4192 0 1 370
box -8 -3 16 105
use FILL  FILL_10514
timestamp 1677677812
transform 1 0 4200 0 1 370
box -8 -3 16 105
use FILL  FILL_10515
timestamp 1677677812
transform 1 0 4208 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_593
timestamp 1677677812
transform 1 0 4216 0 1 370
box -8 -3 104 105
use FILL  FILL_10516
timestamp 1677677812
transform 1 0 4312 0 1 370
box -8 -3 16 105
use FILL  FILL_10517
timestamp 1677677812
transform 1 0 4320 0 1 370
box -8 -3 16 105
use FILL  FILL_10518
timestamp 1677677812
transform 1 0 4328 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8305
timestamp 1677677812
transform 1 0 4364 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_428
timestamp 1677677812
transform 1 0 4336 0 1 370
box -8 -3 46 105
use INVX2  INVX2_681
timestamp 1677677812
transform 1 0 4376 0 1 370
box -9 -3 26 105
use FILL  FILL_10519
timestamp 1677677812
transform 1 0 4392 0 1 370
box -8 -3 16 105
use FILL  FILL_10520
timestamp 1677677812
transform 1 0 4400 0 1 370
box -8 -3 16 105
use FILL  FILL_10521
timestamp 1677677812
transform 1 0 4408 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8306
timestamp 1677677812
transform 1 0 4436 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_429
timestamp 1677677812
transform -1 0 4456 0 1 370
box -8 -3 46 105
use FILL  FILL_10522
timestamp 1677677812
transform 1 0 4456 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_594
timestamp 1677677812
transform 1 0 4464 0 1 370
box -8 -3 104 105
use INVX2  INVX2_682
timestamp 1677677812
transform -1 0 4576 0 1 370
box -9 -3 26 105
use M3_M2  M3_M2_8307
timestamp 1677677812
transform 1 0 4612 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_430
timestamp 1677677812
transform -1 0 4616 0 1 370
box -8 -3 46 105
use INVX2  INVX2_683
timestamp 1677677812
transform -1 0 4632 0 1 370
box -9 -3 26 105
use FILL  FILL_10523
timestamp 1677677812
transform 1 0 4632 0 1 370
box -8 -3 16 105
use FILL  FILL_10524
timestamp 1677677812
transform 1 0 4640 0 1 370
box -8 -3 16 105
use FILL  FILL_10525
timestamp 1677677812
transform 1 0 4648 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_8308
timestamp 1677677812
transform 1 0 4668 0 1 375
box -3 -3 3 3
use OAI22X1  OAI22X1_431
timestamp 1677677812
transform 1 0 4656 0 1 370
box -8 -3 46 105
use M3_M2  M3_M2_8309
timestamp 1677677812
transform 1 0 4716 0 1 375
box -3 -3 3 3
use M3_M2  M3_M2_8310
timestamp 1677677812
transform 1 0 4748 0 1 375
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_595
timestamp 1677677812
transform 1 0 4696 0 1 370
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_87
timestamp 1677677812
transform 1 0 4819 0 1 370
box -10 -3 10 3
use M2_M1  M2_M1_9379
timestamp 1677677812
transform 1 0 84 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8369
timestamp 1677677812
transform 1 0 132 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9483
timestamp 1677677812
transform 1 0 132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8488
timestamp 1677677812
transform 1 0 4 0 1 275
box -3 -3 3 3
use M3_M2  M3_M2_8335
timestamp 1677677812
transform 1 0 180 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8370
timestamp 1677677812
transform 1 0 172 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9484
timestamp 1677677812
transform 1 0 180 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9380
timestamp 1677677812
transform 1 0 252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9381
timestamp 1677677812
transform 1 0 340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9485
timestamp 1677677812
transform 1 0 300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9486
timestamp 1677677812
transform 1 0 332 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9487
timestamp 1677677812
transform 1 0 340 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8414
timestamp 1677677812
transform 1 0 300 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8415
timestamp 1677677812
transform 1 0 340 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8452
timestamp 1677677812
transform 1 0 332 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8476
timestamp 1677677812
transform 1 0 308 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9382
timestamp 1677677812
transform 1 0 356 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8453
timestamp 1677677812
transform 1 0 356 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8322
timestamp 1677677812
transform 1 0 396 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8336
timestamp 1677677812
transform 1 0 412 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9383
timestamp 1677677812
transform 1 0 396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9384
timestamp 1677677812
transform 1 0 412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9488
timestamp 1677677812
transform 1 0 388 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9489
timestamp 1677677812
transform 1 0 404 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8371
timestamp 1677677812
transform 1 0 444 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8337
timestamp 1677677812
transform 1 0 548 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9385
timestamp 1677677812
transform 1 0 468 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8394
timestamp 1677677812
transform 1 0 468 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9490
timestamp 1677677812
transform 1 0 516 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8395
timestamp 1677677812
transform 1 0 540 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9491
timestamp 1677677812
transform 1 0 548 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9492
timestamp 1677677812
transform 1 0 556 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8416
timestamp 1677677812
transform 1 0 516 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8477
timestamp 1677677812
transform 1 0 532 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8417
timestamp 1677677812
transform 1 0 556 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8396
timestamp 1677677812
transform 1 0 572 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9493
timestamp 1677677812
transform 1 0 580 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8418
timestamp 1677677812
transform 1 0 580 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8338
timestamp 1677677812
transform 1 0 628 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9386
timestamp 1677677812
transform 1 0 604 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9387
timestamp 1677677812
transform 1 0 612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9388
timestamp 1677677812
transform 1 0 628 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9494
timestamp 1677677812
transform 1 0 620 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9495
timestamp 1677677812
transform 1 0 636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9389
timestamp 1677677812
transform 1 0 660 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8397
timestamp 1677677812
transform 1 0 660 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8339
timestamp 1677677812
transform 1 0 748 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9390
timestamp 1677677812
transform 1 0 748 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9496
timestamp 1677677812
transform 1 0 684 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9497
timestamp 1677677812
transform 1 0 740 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8311
timestamp 1677677812
transform 1 0 772 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9391
timestamp 1677677812
transform 1 0 772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9498
timestamp 1677677812
transform 1 0 764 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9499
timestamp 1677677812
transform 1 0 780 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8323
timestamp 1677677812
transform 1 0 796 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9373
timestamp 1677677812
transform 1 0 796 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8340
timestamp 1677677812
transform 1 0 820 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9392
timestamp 1677677812
transform 1 0 820 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9393
timestamp 1677677812
transform 1 0 836 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9394
timestamp 1677677812
transform 1 0 844 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8341
timestamp 1677677812
transform 1 0 892 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9395
timestamp 1677677812
transform 1 0 892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9396
timestamp 1677677812
transform 1 0 908 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9500
timestamp 1677677812
transform 1 0 860 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9501
timestamp 1677677812
transform 1 0 868 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9502
timestamp 1677677812
transform 1 0 884 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9503
timestamp 1677677812
transform 1 0 900 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8419
timestamp 1677677812
transform 1 0 868 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8420
timestamp 1677677812
transform 1 0 884 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8478
timestamp 1677677812
transform 1 0 860 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9504
timestamp 1677677812
transform 1 0 916 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8421
timestamp 1677677812
transform 1 0 908 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9374
timestamp 1677677812
transform 1 0 956 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9397
timestamp 1677677812
transform 1 0 948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9505
timestamp 1677677812
transform 1 0 948 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9375
timestamp 1677677812
transform 1 0 972 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8372
timestamp 1677677812
transform 1 0 972 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8312
timestamp 1677677812
transform 1 0 1004 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8324
timestamp 1677677812
transform 1 0 1020 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9398
timestamp 1677677812
transform 1 0 1012 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9506
timestamp 1677677812
transform 1 0 1020 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9507
timestamp 1677677812
transform 1 0 1084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9508
timestamp 1677677812
transform 1 0 1092 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8454
timestamp 1677677812
transform 1 0 1084 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9509
timestamp 1677677812
transform 1 0 1108 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9399
timestamp 1677677812
transform 1 0 1124 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8398
timestamp 1677677812
transform 1 0 1124 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9400
timestamp 1677677812
transform 1 0 1180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9401
timestamp 1677677812
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8399
timestamp 1677677812
transform 1 0 1180 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9402
timestamp 1677677812
transform 1 0 1220 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9510
timestamp 1677677812
transform 1 0 1212 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9511
timestamp 1677677812
transform 1 0 1228 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8422
timestamp 1677677812
transform 1 0 1228 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8467
timestamp 1677677812
transform 1 0 1212 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8342
timestamp 1677677812
transform 1 0 1244 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9403
timestamp 1677677812
transform 1 0 1244 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9404
timestamp 1677677812
transform 1 0 1268 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9405
timestamp 1677677812
transform 1 0 1284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9512
timestamp 1677677812
transform 1 0 1276 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9513
timestamp 1677677812
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8423
timestamp 1677677812
transform 1 0 1292 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8468
timestamp 1677677812
transform 1 0 1276 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9406
timestamp 1677677812
transform 1 0 1324 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9407
timestamp 1677677812
transform 1 0 1332 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8400
timestamp 1677677812
transform 1 0 1324 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8424
timestamp 1677677812
transform 1 0 1332 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8343
timestamp 1677677812
transform 1 0 1348 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9408
timestamp 1677677812
transform 1 0 1348 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9409
timestamp 1677677812
transform 1 0 1372 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9514
timestamp 1677677812
transform 1 0 1340 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9515
timestamp 1677677812
transform 1 0 1348 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9516
timestamp 1677677812
transform 1 0 1364 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9517
timestamp 1677677812
transform 1 0 1380 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8401
timestamp 1677677812
transform 1 0 1388 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9518
timestamp 1677677812
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8425
timestamp 1677677812
transform 1 0 1364 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8426
timestamp 1677677812
transform 1 0 1380 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8469
timestamp 1677677812
transform 1 0 1348 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8470
timestamp 1677677812
transform 1 0 1404 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8313
timestamp 1677677812
transform 1 0 1500 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9410
timestamp 1677677812
transform 1 0 1500 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9411
timestamp 1677677812
transform 1 0 1516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9519
timestamp 1677677812
transform 1 0 1476 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9520
timestamp 1677677812
transform 1 0 1516 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8427
timestamp 1677677812
transform 1 0 1436 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8428
timestamp 1677677812
transform 1 0 1452 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8429
timestamp 1677677812
transform 1 0 1476 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8430
timestamp 1677677812
transform 1 0 1516 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8431
timestamp 1677677812
transform 1 0 1572 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8373
timestamp 1677677812
transform 1 0 1588 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8479
timestamp 1677677812
transform 1 0 1580 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8314
timestamp 1677677812
transform 1 0 1620 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9412
timestamp 1677677812
transform 1 0 1612 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9521
timestamp 1677677812
transform 1 0 1644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9522
timestamp 1677677812
transform 1 0 1692 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8325
timestamp 1677677812
transform 1 0 1748 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9413
timestamp 1677677812
transform 1 0 1732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9414
timestamp 1677677812
transform 1 0 1748 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8374
timestamp 1677677812
transform 1 0 1756 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9523
timestamp 1677677812
transform 1 0 1740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9524
timestamp 1677677812
transform 1 0 1756 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8432
timestamp 1677677812
transform 1 0 1740 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9415
timestamp 1677677812
transform 1 0 1772 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9416
timestamp 1677677812
transform 1 0 1780 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9417
timestamp 1677677812
transform 1 0 1796 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8375
timestamp 1677677812
transform 1 0 1804 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9525
timestamp 1677677812
transform 1 0 1788 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9526
timestamp 1677677812
transform 1 0 1804 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8433
timestamp 1677677812
transform 1 0 1788 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8455
timestamp 1677677812
transform 1 0 1796 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9527
timestamp 1677677812
transform 1 0 1828 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8344
timestamp 1677677812
transform 1 0 1844 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9418
timestamp 1677677812
transform 1 0 1844 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9419
timestamp 1677677812
transform 1 0 1932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9528
timestamp 1677677812
transform 1 0 1908 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8434
timestamp 1677677812
transform 1 0 1908 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9420
timestamp 1677677812
transform 1 0 1956 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9529
timestamp 1677677812
transform 1 0 1948 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8435
timestamp 1677677812
transform 1 0 1948 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8345
timestamp 1677677812
transform 1 0 1972 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9421
timestamp 1677677812
transform 1 0 1972 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8376
timestamp 1677677812
transform 1 0 1980 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9530
timestamp 1677677812
transform 1 0 1972 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8402
timestamp 1677677812
transform 1 0 1996 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9422
timestamp 1677677812
transform 1 0 2004 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9423
timestamp 1677677812
transform 1 0 2036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9424
timestamp 1677677812
transform 1 0 2044 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9531
timestamp 1677677812
transform 1 0 2028 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8403
timestamp 1677677812
transform 1 0 2036 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9532
timestamp 1677677812
transform 1 0 2060 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8346
timestamp 1677677812
transform 1 0 2108 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9533
timestamp 1677677812
transform 1 0 2100 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8347
timestamp 1677677812
transform 1 0 2140 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8348
timestamp 1677677812
transform 1 0 2220 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9425
timestamp 1677677812
transform 1 0 2140 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8377
timestamp 1677677812
transform 1 0 2220 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9534
timestamp 1677677812
transform 1 0 2172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9535
timestamp 1677677812
transform 1 0 2220 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8349
timestamp 1677677812
transform 1 0 2252 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9426
timestamp 1677677812
transform 1 0 2252 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9536
timestamp 1677677812
transform 1 0 2300 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9537
timestamp 1677677812
transform 1 0 2332 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8480
timestamp 1677677812
transform 1 0 2284 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8481
timestamp 1677677812
transform 1 0 2308 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8350
timestamp 1677677812
transform 1 0 2436 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9427
timestamp 1677677812
transform 1 0 2436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9538
timestamp 1677677812
transform 1 0 2356 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9539
timestamp 1677677812
transform 1 0 2412 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8436
timestamp 1677677812
transform 1 0 2412 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8351
timestamp 1677677812
transform 1 0 2460 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8378
timestamp 1677677812
transform 1 0 2468 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9540
timestamp 1677677812
transform 1 0 2476 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8437
timestamp 1677677812
transform 1 0 2476 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9428
timestamp 1677677812
transform 1 0 2492 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8438
timestamp 1677677812
transform 1 0 2492 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9429
timestamp 1677677812
transform 1 0 2540 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9541
timestamp 1677677812
transform 1 0 2572 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8439
timestamp 1677677812
transform 1 0 2572 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9376
timestamp 1677677812
transform 1 0 2604 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9430
timestamp 1677677812
transform 1 0 2596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9593
timestamp 1677677812
transform 1 0 2588 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_9600
timestamp 1677677812
transform 1 0 2596 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_8440
timestamp 1677677812
transform 1 0 2628 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9542
timestamp 1677677812
transform 1 0 2644 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8326
timestamp 1677677812
transform 1 0 2668 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9431
timestamp 1677677812
transform 1 0 2668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9543
timestamp 1677677812
transform 1 0 2660 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8441
timestamp 1677677812
transform 1 0 2660 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9377
timestamp 1677677812
transform 1 0 2676 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_8379
timestamp 1677677812
transform 1 0 2676 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8327
timestamp 1677677812
transform 1 0 2708 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9544
timestamp 1677677812
transform 1 0 2708 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8482
timestamp 1677677812
transform 1 0 2716 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8352
timestamp 1677677812
transform 1 0 2732 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9432
timestamp 1677677812
transform 1 0 2732 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9433
timestamp 1677677812
transform 1 0 2748 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8380
timestamp 1677677812
transform 1 0 2844 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9434
timestamp 1677677812
transform 1 0 2852 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9545
timestamp 1677677812
transform 1 0 2796 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9546
timestamp 1677677812
transform 1 0 2828 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9547
timestamp 1677677812
transform 1 0 2836 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9435
timestamp 1677677812
transform 1 0 2868 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8381
timestamp 1677677812
transform 1 0 2892 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9548
timestamp 1677677812
transform 1 0 2876 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9549
timestamp 1677677812
transform 1 0 2892 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8483
timestamp 1677677812
transform 1 0 2876 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9436
timestamp 1677677812
transform 1 0 2924 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8353
timestamp 1677677812
transform 1 0 3028 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8354
timestamp 1677677812
transform 1 0 3044 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9437
timestamp 1677677812
transform 1 0 2940 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9438
timestamp 1677677812
transform 1 0 3028 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9550
timestamp 1677677812
transform 1 0 2964 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9551
timestamp 1677677812
transform 1 0 3028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9552
timestamp 1677677812
transform 1 0 3044 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9553
timestamp 1677677812
transform 1 0 3052 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9594
timestamp 1677677812
transform 1 0 3044 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8456
timestamp 1677677812
transform 1 0 3044 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8315
timestamp 1677677812
transform 1 0 3084 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9439
timestamp 1677677812
transform 1 0 3084 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9554
timestamp 1677677812
transform 1 0 3076 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9440
timestamp 1677677812
transform 1 0 3108 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9441
timestamp 1677677812
transform 1 0 3116 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8404
timestamp 1677677812
transform 1 0 3116 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8484
timestamp 1677677812
transform 1 0 3108 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8457
timestamp 1677677812
transform 1 0 3148 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9555
timestamp 1677677812
transform 1 0 3156 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8471
timestamp 1677677812
transform 1 0 3156 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8355
timestamp 1677677812
transform 1 0 3260 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9378
timestamp 1677677812
transform 1 0 3276 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_9442
timestamp 1677677812
transform 1 0 3172 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9443
timestamp 1677677812
transform 1 0 3260 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9444
timestamp 1677677812
transform 1 0 3284 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9556
timestamp 1677677812
transform 1 0 3196 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9557
timestamp 1677677812
transform 1 0 3260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9558
timestamp 1677677812
transform 1 0 3276 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8405
timestamp 1677677812
transform 1 0 3284 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9559
timestamp 1677677812
transform 1 0 3292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8442
timestamp 1677677812
transform 1 0 3260 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8458
timestamp 1677677812
transform 1 0 3196 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8459
timestamp 1677677812
transform 1 0 3276 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8443
timestamp 1677677812
transform 1 0 3292 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8460
timestamp 1677677812
transform 1 0 3332 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8328
timestamp 1677677812
transform 1 0 3348 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8382
timestamp 1677677812
transform 1 0 3356 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9445
timestamp 1677677812
transform 1 0 3364 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9560
timestamp 1677677812
transform 1 0 3356 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8406
timestamp 1677677812
transform 1 0 3372 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9595
timestamp 1677677812
transform 1 0 3356 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8444
timestamp 1677677812
transform 1 0 3364 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8461
timestamp 1677677812
transform 1 0 3356 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9446
timestamp 1677677812
transform 1 0 3396 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9561
timestamp 1677677812
transform 1 0 3388 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8407
timestamp 1677677812
transform 1 0 3396 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9596
timestamp 1677677812
transform 1 0 3388 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8462
timestamp 1677677812
transform 1 0 3388 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8356
timestamp 1677677812
transform 1 0 3404 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9447
timestamp 1677677812
transform 1 0 3412 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9562
timestamp 1677677812
transform 1 0 3404 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9448
timestamp 1677677812
transform 1 0 3428 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9563
timestamp 1677677812
transform 1 0 3420 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8445
timestamp 1677677812
transform 1 0 3428 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8446
timestamp 1677677812
transform 1 0 3444 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8472
timestamp 1677677812
transform 1 0 3436 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8329
timestamp 1677677812
transform 1 0 3468 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8383
timestamp 1677677812
transform 1 0 3460 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9449
timestamp 1677677812
transform 1 0 3468 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9597
timestamp 1677677812
transform 1 0 3468 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8463
timestamp 1677677812
transform 1 0 3484 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8485
timestamp 1677677812
transform 1 0 3492 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8357
timestamp 1677677812
transform 1 0 3524 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9450
timestamp 1677677812
transform 1 0 3516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9598
timestamp 1677677812
transform 1 0 3516 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8473
timestamp 1677677812
transform 1 0 3516 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_9451
timestamp 1677677812
transform 1 0 3524 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9564
timestamp 1677677812
transform 1 0 3524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9565
timestamp 1677677812
transform 1 0 3532 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8316
timestamp 1677677812
transform 1 0 3564 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_9599
timestamp 1677677812
transform 1 0 3556 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_8474
timestamp 1677677812
transform 1 0 3540 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8475
timestamp 1677677812
transform 1 0 3556 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_8358
timestamp 1677677812
transform 1 0 3572 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9452
timestamp 1677677812
transform 1 0 3572 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9453
timestamp 1677677812
transform 1 0 3580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9454
timestamp 1677677812
transform 1 0 3612 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8359
timestamp 1677677812
transform 1 0 3652 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9455
timestamp 1677677812
transform 1 0 3652 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8384
timestamp 1677677812
transform 1 0 3660 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9456
timestamp 1677677812
transform 1 0 3668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9566
timestamp 1677677812
transform 1 0 3644 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9567
timestamp 1677677812
transform 1 0 3660 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8464
timestamp 1677677812
transform 1 0 3660 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8385
timestamp 1677677812
transform 1 0 3692 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9568
timestamp 1677677812
transform 1 0 3700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9457
timestamp 1677677812
transform 1 0 3724 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8465
timestamp 1677677812
transform 1 0 3716 0 1 305
box -3 -3 3 3
use M3_M2  M3_M2_8317
timestamp 1677677812
transform 1 0 3764 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8360
timestamp 1677677812
transform 1 0 3820 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9458
timestamp 1677677812
transform 1 0 3772 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8386
timestamp 1677677812
transform 1 0 3836 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9569
timestamp 1677677812
transform 1 0 3820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9570
timestamp 1677677812
transform 1 0 3852 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9571
timestamp 1677677812
transform 1 0 3860 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8318
timestamp 1677677812
transform 1 0 3876 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8330
timestamp 1677677812
transform 1 0 3892 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8331
timestamp 1677677812
transform 1 0 3916 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8361
timestamp 1677677812
transform 1 0 3908 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9459
timestamp 1677677812
transform 1 0 3892 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9460
timestamp 1677677812
transform 1 0 3908 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8387
timestamp 1677677812
transform 1 0 3916 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9572
timestamp 1677677812
transform 1 0 3916 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8388
timestamp 1677677812
transform 1 0 3932 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_8319
timestamp 1677677812
transform 1 0 3980 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8332
timestamp 1677677812
transform 1 0 3980 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8362
timestamp 1677677812
transform 1 0 3948 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_8363
timestamp 1677677812
transform 1 0 3964 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9461
timestamp 1677677812
transform 1 0 3948 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8389
timestamp 1677677812
transform 1 0 3956 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9462
timestamp 1677677812
transform 1 0 3964 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9463
timestamp 1677677812
transform 1 0 3980 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9573
timestamp 1677677812
transform 1 0 3956 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8447
timestamp 1677677812
transform 1 0 3956 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8364
timestamp 1677677812
transform 1 0 4036 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9464
timestamp 1677677812
transform 1 0 4020 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8390
timestamp 1677677812
transform 1 0 4028 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9465
timestamp 1677677812
transform 1 0 4036 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9574
timestamp 1677677812
transform 1 0 4004 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9575
timestamp 1677677812
transform 1 0 4012 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9576
timestamp 1677677812
transform 1 0 4028 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8448
timestamp 1677677812
transform 1 0 4004 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8449
timestamp 1677677812
transform 1 0 4036 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_9466
timestamp 1677677812
transform 1 0 4076 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9467
timestamp 1677677812
transform 1 0 4092 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9468
timestamp 1677677812
transform 1 0 4108 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8408
timestamp 1677677812
transform 1 0 4076 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9577
timestamp 1677677812
transform 1 0 4084 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8466
timestamp 1677677812
transform 1 0 4084 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_9578
timestamp 1677677812
transform 1 0 4116 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9579
timestamp 1677677812
transform 1 0 4132 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8365
timestamp 1677677812
transform 1 0 4164 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9469
timestamp 1677677812
transform 1 0 4164 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8391
timestamp 1677677812
transform 1 0 4172 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9470
timestamp 1677677812
transform 1 0 4180 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9580
timestamp 1677677812
transform 1 0 4156 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9581
timestamp 1677677812
transform 1 0 4172 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8409
timestamp 1677677812
transform 1 0 4180 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8450
timestamp 1677677812
transform 1 0 4156 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8320
timestamp 1677677812
transform 1 0 4276 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8366
timestamp 1677677812
transform 1 0 4228 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9471
timestamp 1677677812
transform 1 0 4204 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8410
timestamp 1677677812
transform 1 0 4204 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_8321
timestamp 1677677812
transform 1 0 4324 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_8367
timestamp 1677677812
transform 1 0 4364 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9472
timestamp 1677677812
transform 1 0 4300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9473
timestamp 1677677812
transform 1 0 4316 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9582
timestamp 1677677812
transform 1 0 4228 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9583
timestamp 1677677812
transform 1 0 4284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9584
timestamp 1677677812
transform 1 0 4292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8451
timestamp 1677677812
transform 1 0 4292 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_8486
timestamp 1677677812
transform 1 0 4268 0 1 285
box -3 -3 3 3
use M3_M2  M3_M2_8411
timestamp 1677677812
transform 1 0 4316 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9585
timestamp 1677677812
transform 1 0 4364 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8487
timestamp 1677677812
transform 1 0 4324 0 1 285
box -3 -3 3 3
use M2_M1  M2_M1_9586
timestamp 1677677812
transform 1 0 4412 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8333
timestamp 1677677812
transform 1 0 4428 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_9474
timestamp 1677677812
transform 1 0 4428 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8334
timestamp 1677677812
transform 1 0 4468 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_8368
timestamp 1677677812
transform 1 0 4460 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_9475
timestamp 1677677812
transform 1 0 4460 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9476
timestamp 1677677812
transform 1 0 4476 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9587
timestamp 1677677812
transform 1 0 4468 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8412
timestamp 1677677812
transform 1 0 4532 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9477
timestamp 1677677812
transform 1 0 4580 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8413
timestamp 1677677812
transform 1 0 4580 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_9478
timestamp 1677677812
transform 1 0 4668 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9588
timestamp 1677677812
transform 1 0 4604 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9589
timestamp 1677677812
transform 1 0 4660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9479
timestamp 1677677812
transform 1 0 4692 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_8392
timestamp 1677677812
transform 1 0 4700 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9480
timestamp 1677677812
transform 1 0 4708 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9481
timestamp 1677677812
transform 1 0 4724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_9590
timestamp 1677677812
transform 1 0 4700 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9591
timestamp 1677677812
transform 1 0 4716 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_8393
timestamp 1677677812
transform 1 0 4740 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_9592
timestamp 1677677812
transform 1 0 4740 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_9482
timestamp 1677677812
transform 1 0 4788 0 1 335
box -2 -2 2 2
use top_level_VIA0  top_level_VIA0_88
timestamp 1677677812
transform 1 0 24 0 1 270
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_558
timestamp 1677677812
transform 1 0 72 0 -1 370
box -8 -3 104 105
use FILL  FILL_10215
timestamp 1677677812
transform 1 0 168 0 -1 370
box -8 -3 16 105
use FILL  FILL_10216
timestamp 1677677812
transform 1 0 176 0 -1 370
box -8 -3 16 105
use FILL  FILL_10217
timestamp 1677677812
transform 1 0 184 0 -1 370
box -8 -3 16 105
use FILL  FILL_10218
timestamp 1677677812
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_10219
timestamp 1677677812
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_10220
timestamp 1677677812
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_10221
timestamp 1677677812
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_10222
timestamp 1677677812
transform 1 0 224 0 -1 370
box -8 -3 16 105
use FILL  FILL_10224
timestamp 1677677812
transform 1 0 232 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8489
timestamp 1677677812
transform 1 0 268 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_561
timestamp 1677677812
transform 1 0 240 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_655
timestamp 1677677812
transform 1 0 336 0 -1 370
box -9 -3 26 105
use FILL  FILL_10239
timestamp 1677677812
transform 1 0 352 0 -1 370
box -8 -3 16 105
use FILL  FILL_10240
timestamp 1677677812
transform 1 0 360 0 -1 370
box -8 -3 16 105
use FILL  FILL_10241
timestamp 1677677812
transform 1 0 368 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_412
timestamp 1677677812
transform 1 0 376 0 -1 370
box -8 -3 46 105
use FILL  FILL_10242
timestamp 1677677812
transform 1 0 416 0 -1 370
box -8 -3 16 105
use FILL  FILL_10243
timestamp 1677677812
transform 1 0 424 0 -1 370
box -8 -3 16 105
use FILL  FILL_10244
timestamp 1677677812
transform 1 0 432 0 -1 370
box -8 -3 16 105
use FILL  FILL_10245
timestamp 1677677812
transform 1 0 440 0 -1 370
box -8 -3 16 105
use FILL  FILL_10246
timestamp 1677677812
transform 1 0 448 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_562
timestamp 1677677812
transform 1 0 456 0 -1 370
box -8 -3 104 105
use FILL  FILL_10247
timestamp 1677677812
transform 1 0 552 0 -1 370
box -8 -3 16 105
use FILL  FILL_10248
timestamp 1677677812
transform 1 0 560 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_656
timestamp 1677677812
transform -1 0 584 0 -1 370
box -9 -3 26 105
use FILL  FILL_10249
timestamp 1677677812
transform 1 0 584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10250
timestamp 1677677812
transform 1 0 592 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_387
timestamp 1677677812
transform 1 0 600 0 -1 370
box -8 -3 46 105
use FILL  FILL_10266
timestamp 1677677812
transform 1 0 640 0 -1 370
box -8 -3 16 105
use M3_M2  M3_M2_8490
timestamp 1677677812
transform 1 0 692 0 1 275
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_565
timestamp 1677677812
transform 1 0 648 0 -1 370
box -8 -3 104 105
use FILL  FILL_10267
timestamp 1677677812
transform 1 0 744 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_414
timestamp 1677677812
transform 1 0 752 0 -1 370
box -8 -3 46 105
use FILL  FILL_10268
timestamp 1677677812
transform 1 0 792 0 -1 370
box -8 -3 16 105
use FILL  FILL_10269
timestamp 1677677812
transform 1 0 800 0 -1 370
box -8 -3 16 105
use FILL  FILL_10270
timestamp 1677677812
transform 1 0 808 0 -1 370
box -8 -3 16 105
use FILL  FILL_10271
timestamp 1677677812
transform 1 0 816 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_110
timestamp 1677677812
transform 1 0 824 0 -1 370
box -8 -3 32 105
use FILL  FILL_10272
timestamp 1677677812
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_10273
timestamp 1677677812
transform 1 0 856 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_388
timestamp 1677677812
transform 1 0 864 0 -1 370
box -8 -3 46 105
use FILL  FILL_10274
timestamp 1677677812
transform 1 0 904 0 -1 370
box -8 -3 16 105
use FILL  FILL_10275
timestamp 1677677812
transform 1 0 912 0 -1 370
box -8 -3 16 105
use FILL  FILL_10276
timestamp 1677677812
transform 1 0 920 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_658
timestamp 1677677812
transform 1 0 928 0 -1 370
box -9 -3 26 105
use FILL  FILL_10277
timestamp 1677677812
transform 1 0 944 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_111
timestamp 1677677812
transform 1 0 952 0 -1 370
box -8 -3 32 105
use FILL  FILL_10278
timestamp 1677677812
transform 1 0 976 0 -1 370
box -8 -3 16 105
use FILL  FILL_10279
timestamp 1677677812
transform 1 0 984 0 -1 370
box -8 -3 16 105
use FILL  FILL_10280
timestamp 1677677812
transform 1 0 992 0 -1 370
box -8 -3 16 105
use FILL  FILL_10281
timestamp 1677677812
transform 1 0 1000 0 -1 370
box -8 -3 16 105
use FILL  FILL_10283
timestamp 1677677812
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_113
timestamp 1677677812
transform 1 0 1016 0 -1 370
box -8 -3 32 105
use FILL  FILL_10285
timestamp 1677677812
transform 1 0 1040 0 -1 370
box -8 -3 16 105
use FILL  FILL_10287
timestamp 1677677812
transform 1 0 1048 0 -1 370
box -8 -3 16 105
use FILL  FILL_10288
timestamp 1677677812
transform 1 0 1056 0 -1 370
box -8 -3 16 105
use FILL  FILL_10289
timestamp 1677677812
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use FILL  FILL_10290
timestamp 1677677812
transform 1 0 1072 0 -1 370
box -8 -3 16 105
use FILL  FILL_10291
timestamp 1677677812
transform 1 0 1080 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_659
timestamp 1677677812
transform -1 0 1104 0 -1 370
box -9 -3 26 105
use FILL  FILL_10292
timestamp 1677677812
transform 1 0 1104 0 -1 370
box -8 -3 16 105
use FILL  FILL_10293
timestamp 1677677812
transform 1 0 1112 0 -1 370
box -8 -3 16 105
use FILL  FILL_10294
timestamp 1677677812
transform 1 0 1120 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_660
timestamp 1677677812
transform -1 0 1144 0 -1 370
box -9 -3 26 105
use FILL  FILL_10295
timestamp 1677677812
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_10297
timestamp 1677677812
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use FILL  FILL_10303
timestamp 1677677812
transform 1 0 1160 0 -1 370
box -8 -3 16 105
use FILL  FILL_10304
timestamp 1677677812
transform 1 0 1168 0 -1 370
box -8 -3 16 105
use FILL  FILL_10305
timestamp 1677677812
transform 1 0 1176 0 -1 370
box -8 -3 16 105
use FILL  FILL_10306
timestamp 1677677812
transform 1 0 1184 0 -1 370
box -8 -3 16 105
use FILL  FILL_10307
timestamp 1677677812
transform 1 0 1192 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_416
timestamp 1677677812
transform -1 0 1240 0 -1 370
box -8 -3 46 105
use FILL  FILL_10308
timestamp 1677677812
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use FILL  FILL_10309
timestamp 1677677812
transform 1 0 1248 0 -1 370
box -8 -3 16 105
use FILL  FILL_10310
timestamp 1677677812
transform 1 0 1256 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_417
timestamp 1677677812
transform -1 0 1304 0 -1 370
box -8 -3 46 105
use FILL  FILL_10311
timestamp 1677677812
transform 1 0 1304 0 -1 370
box -8 -3 16 105
use FILL  FILL_10312
timestamp 1677677812
transform 1 0 1312 0 -1 370
box -8 -3 16 105
use FILL  FILL_10314
timestamp 1677677812
transform 1 0 1320 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_664
timestamp 1677677812
transform 1 0 1328 0 -1 370
box -9 -3 26 105
use AOI22X1  AOI22X1_394
timestamp 1677677812
transform -1 0 1384 0 -1 370
box -8 -3 46 105
use FILL  FILL_10335
timestamp 1677677812
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use FILL  FILL_10336
timestamp 1677677812
transform 1 0 1392 0 -1 370
box -8 -3 16 105
use FILL  FILL_10337
timestamp 1677677812
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use FILL  FILL_10338
timestamp 1677677812
transform 1 0 1408 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_570
timestamp 1677677812
transform -1 0 1512 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_665
timestamp 1677677812
transform 1 0 1512 0 -1 370
box -9 -3 26 105
use FILL  FILL_10339
timestamp 1677677812
transform 1 0 1528 0 -1 370
box -8 -3 16 105
use FILL  FILL_10340
timestamp 1677677812
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use FILL  FILL_10341
timestamp 1677677812
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_10342
timestamp 1677677812
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use FILL  FILL_10343
timestamp 1677677812
transform 1 0 1560 0 -1 370
box -8 -3 16 105
use FILL  FILL_10344
timestamp 1677677812
transform 1 0 1568 0 -1 370
box -8 -3 16 105
use FILL  FILL_10345
timestamp 1677677812
transform 1 0 1576 0 -1 370
box -8 -3 16 105
use FILL  FILL_10346
timestamp 1677677812
transform 1 0 1584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10347
timestamp 1677677812
transform 1 0 1592 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_571
timestamp 1677677812
transform 1 0 1600 0 -1 370
box -8 -3 104 105
use FILL  FILL_10348
timestamp 1677677812
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_10349
timestamp 1677677812
transform 1 0 1704 0 -1 370
box -8 -3 16 105
use FILL  FILL_10350
timestamp 1677677812
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use FILL  FILL_10351
timestamp 1677677812
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_419
timestamp 1677677812
transform -1 0 1768 0 -1 370
box -8 -3 46 105
use FILL  FILL_10352
timestamp 1677677812
transform 1 0 1768 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_420
timestamp 1677677812
transform -1 0 1816 0 -1 370
box -8 -3 46 105
use FILL  FILL_10353
timestamp 1677677812
transform 1 0 1816 0 -1 370
box -8 -3 16 105
use FILL  FILL_10354
timestamp 1677677812
transform 1 0 1824 0 -1 370
box -8 -3 16 105
use FILL  FILL_10355
timestamp 1677677812
transform 1 0 1832 0 -1 370
box -8 -3 16 105
use FILL  FILL_10356
timestamp 1677677812
transform 1 0 1840 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_572
timestamp 1677677812
transform -1 0 1944 0 -1 370
box -8 -3 104 105
use FILL  FILL_10357
timestamp 1677677812
transform 1 0 1944 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_666
timestamp 1677677812
transform 1 0 1952 0 -1 370
box -9 -3 26 105
use FILL  FILL_10358
timestamp 1677677812
transform 1 0 1968 0 -1 370
box -8 -3 16 105
use FILL  FILL_10359
timestamp 1677677812
transform 1 0 1976 0 -1 370
box -8 -3 16 105
use FILL  FILL_10361
timestamp 1677677812
transform 1 0 1984 0 -1 370
box -8 -3 16 105
use FILL  FILL_10365
timestamp 1677677812
transform 1 0 1992 0 -1 370
box -8 -3 16 105
use FILL  FILL_10366
timestamp 1677677812
transform 1 0 2000 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_396
timestamp 1677677812
transform -1 0 2048 0 -1 370
box -8 -3 46 105
use FILL  FILL_10367
timestamp 1677677812
transform 1 0 2048 0 -1 370
box -8 -3 16 105
use FILL  FILL_10369
timestamp 1677677812
transform 1 0 2056 0 -1 370
box -8 -3 16 105
use FILL  FILL_10370
timestamp 1677677812
transform 1 0 2064 0 -1 370
box -8 -3 16 105
use FILL  FILL_10371
timestamp 1677677812
transform 1 0 2072 0 -1 370
box -8 -3 16 105
use FILL  FILL_10373
timestamp 1677677812
transform 1 0 2080 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_668
timestamp 1677677812
transform 1 0 2088 0 -1 370
box -9 -3 26 105
use FILL  FILL_10378
timestamp 1677677812
transform 1 0 2104 0 -1 370
box -8 -3 16 105
use FILL  FILL_10379
timestamp 1677677812
transform 1 0 2112 0 -1 370
box -8 -3 16 105
use FILL  FILL_10380
timestamp 1677677812
transform 1 0 2120 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_575
timestamp 1677677812
transform 1 0 2128 0 -1 370
box -8 -3 104 105
use FILL  FILL_10381
timestamp 1677677812
transform 1 0 2224 0 -1 370
box -8 -3 16 105
use FILL  FILL_10382
timestamp 1677677812
transform 1 0 2232 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_576
timestamp 1677677812
transform 1 0 2240 0 -1 370
box -8 -3 104 105
use FILL  FILL_10383
timestamp 1677677812
transform 1 0 2336 0 -1 370
box -8 -3 16 105
use FILL  FILL_10395
timestamp 1677677812
transform 1 0 2344 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_577
timestamp 1677677812
transform -1 0 2448 0 -1 370
box -8 -3 104 105
use FILL  FILL_10396
timestamp 1677677812
transform 1 0 2448 0 -1 370
box -8 -3 16 105
use FILL  FILL_10398
timestamp 1677677812
transform 1 0 2456 0 -1 370
box -8 -3 16 105
use FILL  FILL_10400
timestamp 1677677812
transform 1 0 2464 0 -1 370
box -8 -3 16 105
use FILL  FILL_10402
timestamp 1677677812
transform 1 0 2472 0 -1 370
box -8 -3 16 105
use FILL  FILL_10404
timestamp 1677677812
transform 1 0 2480 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_177
timestamp 1677677812
transform 1 0 2488 0 -1 370
box -8 -3 34 105
use FILL  FILL_10405
timestamp 1677677812
transform 1 0 2520 0 -1 370
box -8 -3 16 105
use FILL  FILL_10406
timestamp 1677677812
transform 1 0 2528 0 -1 370
box -8 -3 16 105
use FILL  FILL_10407
timestamp 1677677812
transform 1 0 2536 0 -1 370
box -8 -3 16 105
use FILL  FILL_10408
timestamp 1677677812
transform 1 0 2544 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_77
timestamp 1677677812
transform -1 0 2584 0 -1 370
box -8 -3 40 105
use FILL  FILL_10409
timestamp 1677677812
transform 1 0 2584 0 -1 370
box -8 -3 16 105
use FILL  FILL_10410
timestamp 1677677812
transform 1 0 2592 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_116
timestamp 1677677812
transform 1 0 2600 0 -1 370
box -8 -3 32 105
use FILL  FILL_10420
timestamp 1677677812
transform 1 0 2624 0 -1 370
box -8 -3 16 105
use FILL  FILL_10421
timestamp 1677677812
transform 1 0 2632 0 -1 370
box -8 -3 16 105
use FILL  FILL_10422
timestamp 1677677812
transform 1 0 2640 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_671
timestamp 1677677812
transform -1 0 2664 0 -1 370
box -9 -3 26 105
use FILL  FILL_10423
timestamp 1677677812
transform 1 0 2664 0 -1 370
box -8 -3 16 105
use FILL  FILL_10424
timestamp 1677677812
transform 1 0 2672 0 -1 370
box -8 -3 16 105
use FILL  FILL_10425
timestamp 1677677812
transform 1 0 2680 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_117
timestamp 1677677812
transform 1 0 2688 0 -1 370
box -8 -3 32 105
use FILL  FILL_10426
timestamp 1677677812
transform 1 0 2712 0 -1 370
box -8 -3 16 105
use FILL  FILL_10427
timestamp 1677677812
transform 1 0 2720 0 -1 370
box -8 -3 16 105
use FILL  FILL_10428
timestamp 1677677812
transform 1 0 2728 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_582
timestamp 1677677812
transform 1 0 2736 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_672
timestamp 1677677812
transform -1 0 2848 0 -1 370
box -9 -3 26 105
use FILL  FILL_10429
timestamp 1677677812
transform 1 0 2848 0 -1 370
box -8 -3 16 105
use AOI22X1  AOI22X1_397
timestamp 1677677812
transform 1 0 2856 0 -1 370
box -8 -3 46 105
use FILL  FILL_10430
timestamp 1677677812
transform 1 0 2896 0 -1 370
box -8 -3 16 105
use FILL  FILL_10431
timestamp 1677677812
transform 1 0 2904 0 -1 370
box -8 -3 16 105
use FILL  FILL_10432
timestamp 1677677812
transform 1 0 2912 0 -1 370
box -8 -3 16 105
use FILL  FILL_10433
timestamp 1677677812
transform 1 0 2920 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_583
timestamp 1677677812
transform 1 0 2928 0 -1 370
box -8 -3 104 105
use NAND2X1  NAND2X1_47
timestamp 1677677812
transform 1 0 3024 0 -1 370
box -8 -3 32 105
use BUFX2  BUFX2_115
timestamp 1677677812
transform 1 0 3048 0 -1 370
box -5 -3 28 105
use FILL  FILL_10434
timestamp 1677677812
transform 1 0 3072 0 -1 370
box -8 -3 16 105
use FILL  FILL_10439
timestamp 1677677812
transform 1 0 3080 0 -1 370
box -8 -3 16 105
use BUFX2  BUFX2_116
timestamp 1677677812
transform 1 0 3088 0 -1 370
box -5 -3 28 105
use FILL  FILL_10440
timestamp 1677677812
transform 1 0 3112 0 -1 370
box -8 -3 16 105
use FILL  FILL_10441
timestamp 1677677812
transform 1 0 3120 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_674
timestamp 1677677812
transform 1 0 3128 0 -1 370
box -9 -3 26 105
use FILL  FILL_10442
timestamp 1677677812
transform 1 0 3144 0 -1 370
box -8 -3 16 105
use FILL  FILL_10443
timestamp 1677677812
transform 1 0 3152 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_586
timestamp 1677677812
transform 1 0 3160 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_675
timestamp 1677677812
transform 1 0 3256 0 -1 370
box -9 -3 26 105
use NOR2X1  NOR2X1_118
timestamp 1677677812
transform 1 0 3272 0 -1 370
box -8 -3 32 105
use FILL  FILL_10444
timestamp 1677677812
transform 1 0 3296 0 -1 370
box -8 -3 16 105
use FILL  FILL_10445
timestamp 1677677812
transform 1 0 3304 0 -1 370
box -8 -3 16 105
use FILL  FILL_10446
timestamp 1677677812
transform 1 0 3312 0 -1 370
box -8 -3 16 105
use FILL  FILL_10448
timestamp 1677677812
transform 1 0 3320 0 -1 370
box -8 -3 16 105
use FILL  FILL_10450
timestamp 1677677812
transform 1 0 3328 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_50
timestamp 1677677812
transform 1 0 3336 0 -1 370
box -8 -3 32 105
use FILL  FILL_10457
timestamp 1677677812
transform 1 0 3360 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_51
timestamp 1677677812
transform 1 0 3368 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_676
timestamp 1677677812
transform 1 0 3392 0 -1 370
box -9 -3 26 105
use INVX2  INVX2_677
timestamp 1677677812
transform 1 0 3408 0 -1 370
box -9 -3 26 105
use FILL  FILL_10458
timestamp 1677677812
transform 1 0 3424 0 -1 370
box -8 -3 16 105
use FILL  FILL_10460
timestamp 1677677812
transform 1 0 3432 0 -1 370
box -8 -3 16 105
use FILL  FILL_10462
timestamp 1677677812
transform 1 0 3440 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_52
timestamp 1677677812
transform 1 0 3448 0 -1 370
box -8 -3 32 105
use FILL  FILL_10468
timestamp 1677677812
transform 1 0 3472 0 -1 370
box -8 -3 16 105
use FILL  FILL_10469
timestamp 1677677812
transform 1 0 3480 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_181
timestamp 1677677812
transform 1 0 3488 0 -1 370
box -8 -3 34 105
use FILL  FILL_10470
timestamp 1677677812
transform 1 0 3520 0 -1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_182
timestamp 1677677812
transform 1 0 3528 0 -1 370
box -8 -3 34 105
use FILL  FILL_10471
timestamp 1677677812
transform 1 0 3560 0 -1 370
box -8 -3 16 105
use FILL  FILL_10472
timestamp 1677677812
transform 1 0 3568 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_678
timestamp 1677677812
transform 1 0 3576 0 -1 370
box -9 -3 26 105
use FILL  FILL_10473
timestamp 1677677812
transform 1 0 3592 0 -1 370
box -8 -3 16 105
use FILL  FILL_10474
timestamp 1677677812
transform 1 0 3600 0 -1 370
box -8 -3 16 105
use FILL  FILL_10475
timestamp 1677677812
transform 1 0 3608 0 -1 370
box -8 -3 16 105
use FILL  FILL_10476
timestamp 1677677812
transform 1 0 3616 0 -1 370
box -8 -3 16 105
use FILL  FILL_10477
timestamp 1677677812
transform 1 0 3624 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_421
timestamp 1677677812
transform 1 0 3632 0 -1 370
box -8 -3 46 105
use FILL  FILL_10478
timestamp 1677677812
transform 1 0 3672 0 -1 370
box -8 -3 16 105
use FILL  FILL_10480
timestamp 1677677812
transform 1 0 3680 0 -1 370
box -8 -3 16 105
use FILL  FILL_10482
timestamp 1677677812
transform 1 0 3688 0 -1 370
box -8 -3 16 105
use FILL  FILL_10483
timestamp 1677677812
transform 1 0 3696 0 -1 370
box -8 -3 16 105
use FILL  FILL_10484
timestamp 1677677812
transform 1 0 3704 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_679
timestamp 1677677812
transform -1 0 3728 0 -1 370
box -9 -3 26 105
use FILL  FILL_10485
timestamp 1677677812
transform 1 0 3728 0 -1 370
box -8 -3 16 105
use FILL  FILL_10487
timestamp 1677677812
transform 1 0 3736 0 -1 370
box -8 -3 16 105
use FILL  FILL_10489
timestamp 1677677812
transform 1 0 3744 0 -1 370
box -8 -3 16 105
use FILL  FILL_10495
timestamp 1677677812
transform 1 0 3752 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_592
timestamp 1677677812
transform 1 0 3760 0 -1 370
box -8 -3 104 105
use FILL  FILL_10496
timestamp 1677677812
transform 1 0 3856 0 -1 370
box -8 -3 16 105
use FILL  FILL_10497
timestamp 1677677812
transform 1 0 3864 0 -1 370
box -8 -3 16 105
use FILL  FILL_10498
timestamp 1677677812
transform 1 0 3872 0 -1 370
box -8 -3 16 105
use FILL  FILL_10499
timestamp 1677677812
transform 1 0 3880 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_423
timestamp 1677677812
transform 1 0 3888 0 -1 370
box -8 -3 46 105
use FILL  FILL_10500
timestamp 1677677812
transform 1 0 3928 0 -1 370
box -8 -3 16 105
use FILL  FILL_10501
timestamp 1677677812
transform 1 0 3936 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_424
timestamp 1677677812
transform -1 0 3984 0 -1 370
box -8 -3 46 105
use FILL  FILL_10502
timestamp 1677677812
transform 1 0 3984 0 -1 370
box -8 -3 16 105
use FILL  FILL_10503
timestamp 1677677812
transform 1 0 3992 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_425
timestamp 1677677812
transform 1 0 4000 0 -1 370
box -8 -3 46 105
use FILL  FILL_10504
timestamp 1677677812
transform 1 0 4040 0 -1 370
box -8 -3 16 105
use FILL  FILL_10505
timestamp 1677677812
transform 1 0 4048 0 -1 370
box -8 -3 16 105
use FILL  FILL_10506
timestamp 1677677812
transform 1 0 4056 0 -1 370
box -8 -3 16 105
use FILL  FILL_10507
timestamp 1677677812
transform 1 0 4064 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_426
timestamp 1677677812
transform -1 0 4112 0 -1 370
box -8 -3 46 105
use FILL  FILL_10508
timestamp 1677677812
transform 1 0 4112 0 -1 370
box -8 -3 16 105
use FILL  FILL_10509
timestamp 1677677812
transform 1 0 4120 0 -1 370
box -8 -3 16 105
use FILL  FILL_10510
timestamp 1677677812
transform 1 0 4128 0 -1 370
box -8 -3 16 105
use FILL  FILL_10511
timestamp 1677677812
transform 1 0 4136 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_427
timestamp 1677677812
transform 1 0 4144 0 -1 370
box -8 -3 46 105
use FILL  FILL_10512
timestamp 1677677812
transform 1 0 4184 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_596
timestamp 1677677812
transform 1 0 4192 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_684
timestamp 1677677812
transform -1 0 4304 0 -1 370
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_597
timestamp 1677677812
transform 1 0 4304 0 -1 370
box -8 -3 104 105
use INVX2  INVX2_685
timestamp 1677677812
transform 1 0 4400 0 -1 370
box -9 -3 26 105
use FILL  FILL_10526
timestamp 1677677812
transform 1 0 4416 0 -1 370
box -8 -3 16 105
use FILL  FILL_10527
timestamp 1677677812
transform 1 0 4424 0 -1 370
box -8 -3 16 105
use FILL  FILL_10528
timestamp 1677677812
transform 1 0 4432 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_432
timestamp 1677677812
transform 1 0 4440 0 -1 370
box -8 -3 46 105
use FILL  FILL_10529
timestamp 1677677812
transform 1 0 4480 0 -1 370
box -8 -3 16 105
use FILL  FILL_10530
timestamp 1677677812
transform 1 0 4488 0 -1 370
box -8 -3 16 105
use FILL  FILL_10531
timestamp 1677677812
transform 1 0 4496 0 -1 370
box -8 -3 16 105
use FILL  FILL_10532
timestamp 1677677812
transform 1 0 4504 0 -1 370
box -8 -3 16 105
use FILL  FILL_10533
timestamp 1677677812
transform 1 0 4512 0 -1 370
box -8 -3 16 105
use FILL  FILL_10534
timestamp 1677677812
transform 1 0 4520 0 -1 370
box -8 -3 16 105
use FILL  FILL_10535
timestamp 1677677812
transform 1 0 4528 0 -1 370
box -8 -3 16 105
use FILL  FILL_10536
timestamp 1677677812
transform 1 0 4536 0 -1 370
box -8 -3 16 105
use FILL  FILL_10537
timestamp 1677677812
transform 1 0 4544 0 -1 370
box -8 -3 16 105
use FILL  FILL_10538
timestamp 1677677812
transform 1 0 4552 0 -1 370
box -8 -3 16 105
use FILL  FILL_10539
timestamp 1677677812
transform 1 0 4560 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_598
timestamp 1677677812
transform 1 0 4568 0 -1 370
box -8 -3 104 105
use FILL  FILL_10540
timestamp 1677677812
transform 1 0 4664 0 -1 370
box -8 -3 16 105
use FILL  FILL_10541
timestamp 1677677812
transform 1 0 4672 0 -1 370
box -8 -3 16 105
use FILL  FILL_10542
timestamp 1677677812
transform 1 0 4680 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_433
timestamp 1677677812
transform 1 0 4688 0 -1 370
box -8 -3 46 105
use INVX2  INVX2_686
timestamp 1677677812
transform -1 0 4744 0 -1 370
box -9 -3 26 105
use FILL  FILL_10543
timestamp 1677677812
transform 1 0 4744 0 -1 370
box -8 -3 16 105
use FILL  FILL_10544
timestamp 1677677812
transform 1 0 4752 0 -1 370
box -8 -3 16 105
use FILL  FILL_10545
timestamp 1677677812
transform 1 0 4760 0 -1 370
box -8 -3 16 105
use FILL  FILL_10546
timestamp 1677677812
transform 1 0 4768 0 -1 370
box -8 -3 16 105
use FILL  FILL_10547
timestamp 1677677812
transform 1 0 4776 0 -1 370
box -8 -3 16 105
use FILL  FILL_10548
timestamp 1677677812
transform 1 0 4784 0 -1 370
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_89
timestamp 1677677812
transform 1 0 4843 0 1 270
box -10 -3 10 3
use M3_M2  M3_M2_8523
timestamp 1677677812
transform 1 0 164 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8546
timestamp 1677677812
transform 1 0 132 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8547
timestamp 1677677812
transform 1 0 172 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9610
timestamp 1677677812
transform 1 0 132 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9611
timestamp 1677677812
transform 1 0 164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9612
timestamp 1677677812
transform 1 0 172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9751
timestamp 1677677812
transform 1 0 84 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8632
timestamp 1677677812
transform 1 0 84 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8633
timestamp 1677677812
transform 1 0 148 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8497
timestamp 1677677812
transform 1 0 220 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8524
timestamp 1677677812
transform 1 0 196 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8548
timestamp 1677677812
transform 1 0 188 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8549
timestamp 1677677812
transform 1 0 228 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8550
timestamp 1677677812
transform 1 0 300 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9613
timestamp 1677677812
transform 1 0 188 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9614
timestamp 1677677812
transform 1 0 204 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9615
timestamp 1677677812
transform 1 0 220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9616
timestamp 1677677812
transform 1 0 228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9617
timestamp 1677677812
transform 1 0 244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9618
timestamp 1677677812
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9619
timestamp 1677677812
transform 1 0 284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9752
timestamp 1677677812
transform 1 0 188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9753
timestamp 1677677812
transform 1 0 196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9754
timestamp 1677677812
transform 1 0 212 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9755
timestamp 1677677812
transform 1 0 220 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9756
timestamp 1677677812
transform 1 0 228 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9757
timestamp 1677677812
transform 1 0 252 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8634
timestamp 1677677812
transform 1 0 220 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8635
timestamp 1677677812
transform 1 0 252 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8687
timestamp 1677677812
transform 1 0 228 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8594
timestamp 1677677812
transform 1 0 292 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8498
timestamp 1677677812
transform 1 0 348 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8511
timestamp 1677677812
transform 1 0 340 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8491
timestamp 1677677812
transform 1 0 404 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8512
timestamp 1677677812
transform 1 0 380 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8513
timestamp 1677677812
transform 1 0 396 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8514
timestamp 1677677812
transform 1 0 428 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8551
timestamp 1677677812
transform 1 0 340 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8552
timestamp 1677677812
transform 1 0 364 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9620
timestamp 1677677812
transform 1 0 300 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9621
timestamp 1677677812
transform 1 0 308 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9622
timestamp 1677677812
transform 1 0 324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9623
timestamp 1677677812
transform 1 0 340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9624
timestamp 1677677812
transform 1 0 348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9625
timestamp 1677677812
transform 1 0 364 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9626
timestamp 1677677812
transform 1 0 380 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8595
timestamp 1677677812
transform 1 0 388 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8525
timestamp 1677677812
transform 1 0 460 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9627
timestamp 1677677812
transform 1 0 396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9628
timestamp 1677677812
transform 1 0 412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9629
timestamp 1677677812
transform 1 0 428 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9630
timestamp 1677677812
transform 1 0 452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9758
timestamp 1677677812
transform 1 0 276 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9759
timestamp 1677677812
transform 1 0 292 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9760
timestamp 1677677812
transform 1 0 300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9761
timestamp 1677677812
transform 1 0 332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9762
timestamp 1677677812
transform 1 0 340 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9763
timestamp 1677677812
transform 1 0 356 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9764
timestamp 1677677812
transform 1 0 380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9765
timestamp 1677677812
transform 1 0 388 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9766
timestamp 1677677812
transform 1 0 404 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8636
timestamp 1677677812
transform 1 0 276 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8637
timestamp 1677677812
transform 1 0 300 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8638
timestamp 1677677812
transform 1 0 340 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8619
timestamp 1677677812
transform 1 0 412 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9767
timestamp 1677677812
transform 1 0 420 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9768
timestamp 1677677812
transform 1 0 428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9769
timestamp 1677677812
transform 1 0 444 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8639
timestamp 1677677812
transform 1 0 380 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8620
timestamp 1677677812
transform 1 0 452 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8553
timestamp 1677677812
transform 1 0 468 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9770
timestamp 1677677812
transform 1 0 460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9771
timestamp 1677677812
transform 1 0 468 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8640
timestamp 1677677812
transform 1 0 428 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8688
timestamp 1677677812
transform 1 0 420 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9631
timestamp 1677677812
transform 1 0 476 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9632
timestamp 1677677812
transform 1 0 532 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8554
timestamp 1677677812
transform 1 0 548 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9633
timestamp 1677677812
transform 1 0 556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9772
timestamp 1677677812
transform 1 0 548 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8499
timestamp 1677677812
transform 1 0 580 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8555
timestamp 1677677812
transform 1 0 612 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9634
timestamp 1677677812
transform 1 0 636 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8556
timestamp 1677677812
transform 1 0 668 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8596
timestamp 1677677812
transform 1 0 652 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9635
timestamp 1677677812
transform 1 0 660 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9773
timestamp 1677677812
transform 1 0 644 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9774
timestamp 1677677812
transform 1 0 652 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9775
timestamp 1677677812
transform 1 0 668 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9776
timestamp 1677677812
transform 1 0 676 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8641
timestamp 1677677812
transform 1 0 652 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8500
timestamp 1677677812
transform 1 0 692 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9636
timestamp 1677677812
transform 1 0 692 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8515
timestamp 1677677812
transform 1 0 716 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8516
timestamp 1677677812
transform 1 0 764 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9637
timestamp 1677677812
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9638
timestamp 1677677812
transform 1 0 716 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9639
timestamp 1677677812
transform 1 0 740 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8597
timestamp 1677677812
transform 1 0 756 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9640
timestamp 1677677812
transform 1 0 764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9641
timestamp 1677677812
transform 1 0 780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9777
timestamp 1677677812
transform 1 0 716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9778
timestamp 1677677812
transform 1 0 732 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8621
timestamp 1677677812
transform 1 0 740 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9779
timestamp 1677677812
transform 1 0 748 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9780
timestamp 1677677812
transform 1 0 756 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9781
timestamp 1677677812
transform 1 0 772 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8642
timestamp 1677677812
transform 1 0 716 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8643
timestamp 1677677812
transform 1 0 732 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8622
timestamp 1677677812
transform 1 0 780 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8644
timestamp 1677677812
transform 1 0 788 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9892
timestamp 1677677812
transform 1 0 796 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_8689
timestamp 1677677812
transform 1 0 772 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8598
timestamp 1677677812
transform 1 0 812 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9782
timestamp 1677677812
transform 1 0 812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9783
timestamp 1677677812
transform 1 0 820 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9784
timestamp 1677677812
transform 1 0 828 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9893
timestamp 1677677812
transform 1 0 828 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_8690
timestamp 1677677812
transform 1 0 828 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8557
timestamp 1677677812
transform 1 0 852 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9642
timestamp 1677677812
transform 1 0 852 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8645
timestamp 1677677812
transform 1 0 844 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8517
timestamp 1677677812
transform 1 0 868 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8526
timestamp 1677677812
transform 1 0 884 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9643
timestamp 1677677812
transform 1 0 884 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9644
timestamp 1677677812
transform 1 0 892 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8492
timestamp 1677677812
transform 1 0 956 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9645
timestamp 1677677812
transform 1 0 948 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9646
timestamp 1677677812
transform 1 0 996 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8623
timestamp 1677677812
transform 1 0 900 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9785
timestamp 1677677812
transform 1 0 980 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8501
timestamp 1677677812
transform 1 0 1044 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9647
timestamp 1677677812
transform 1 0 1004 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8599
timestamp 1677677812
transform 1 0 1020 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9648
timestamp 1677677812
transform 1 0 1028 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9649
timestamp 1677677812
transform 1 0 1044 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8624
timestamp 1677677812
transform 1 0 1004 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9786
timestamp 1677677812
transform 1 0 1012 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9787
timestamp 1677677812
transform 1 0 1020 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9788
timestamp 1677677812
transform 1 0 1036 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8625
timestamp 1677677812
transform 1 0 1044 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8646
timestamp 1677677812
transform 1 0 1036 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9650
timestamp 1677677812
transform 1 0 1092 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9789
timestamp 1677677812
transform 1 0 1068 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8518
timestamp 1677677812
transform 1 0 1164 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8502
timestamp 1677677812
transform 1 0 1236 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8558
timestamp 1677677812
transform 1 0 1220 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9651
timestamp 1677677812
transform 1 0 1156 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9652
timestamp 1677677812
transform 1 0 1164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9653
timestamp 1677677812
transform 1 0 1180 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9654
timestamp 1677677812
transform 1 0 1196 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9655
timestamp 1677677812
transform 1 0 1212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9656
timestamp 1677677812
transform 1 0 1228 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8600
timestamp 1677677812
transform 1 0 1236 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9657
timestamp 1677677812
transform 1 0 1244 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9790
timestamp 1677677812
transform 1 0 1164 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9791
timestamp 1677677812
transform 1 0 1188 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9792
timestamp 1677677812
transform 1 0 1196 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9793
timestamp 1677677812
transform 1 0 1220 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8647
timestamp 1677677812
transform 1 0 1156 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8648
timestamp 1677677812
transform 1 0 1188 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8519
timestamp 1677677812
transform 1 0 1276 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8493
timestamp 1677677812
transform 1 0 1292 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8527
timestamp 1677677812
transform 1 0 1284 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9794
timestamp 1677677812
transform 1 0 1284 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8649
timestamp 1677677812
transform 1 0 1284 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8503
timestamp 1677677812
transform 1 0 1372 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9658
timestamp 1677677812
transform 1 0 1340 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9795
timestamp 1677677812
transform 1 0 1372 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8691
timestamp 1677677812
transform 1 0 1372 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9796
timestamp 1677677812
transform 1 0 1388 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8504
timestamp 1677677812
transform 1 0 1428 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8559
timestamp 1677677812
transform 1 0 1404 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8528
timestamp 1677677812
transform 1 0 1436 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9659
timestamp 1677677812
transform 1 0 1404 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9660
timestamp 1677677812
transform 1 0 1420 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8650
timestamp 1677677812
transform 1 0 1396 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8601
timestamp 1677677812
transform 1 0 1428 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9661
timestamp 1677677812
transform 1 0 1436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9797
timestamp 1677677812
transform 1 0 1412 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9798
timestamp 1677677812
transform 1 0 1428 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9799
timestamp 1677677812
transform 1 0 1436 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8560
timestamp 1677677812
transform 1 0 1468 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9662
timestamp 1677677812
transform 1 0 1460 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9663
timestamp 1677677812
transform 1 0 1468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9800
timestamp 1677677812
transform 1 0 1468 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8651
timestamp 1677677812
transform 1 0 1468 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8529
timestamp 1677677812
transform 1 0 1524 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8561
timestamp 1677677812
transform 1 0 1516 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9664
timestamp 1677677812
transform 1 0 1508 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9665
timestamp 1677677812
transform 1 0 1524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9801
timestamp 1677677812
transform 1 0 1516 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9802
timestamp 1677677812
transform 1 0 1524 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8692
timestamp 1677677812
transform 1 0 1492 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8494
timestamp 1677677812
transform 1 0 1588 0 1 265
box -3 -3 3 3
use M3_M2  M3_M2_8520
timestamp 1677677812
transform 1 0 1572 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8562
timestamp 1677677812
transform 1 0 1604 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9666
timestamp 1677677812
transform 1 0 1572 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9667
timestamp 1677677812
transform 1 0 1588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9668
timestamp 1677677812
transform 1 0 1604 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8602
timestamp 1677677812
transform 1 0 1612 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9669
timestamp 1677677812
transform 1 0 1620 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9803
timestamp 1677677812
transform 1 0 1564 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9804
timestamp 1677677812
transform 1 0 1580 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9805
timestamp 1677677812
transform 1 0 1604 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9806
timestamp 1677677812
transform 1 0 1612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9807
timestamp 1677677812
transform 1 0 1628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8652
timestamp 1677677812
transform 1 0 1564 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8653
timestamp 1677677812
transform 1 0 1628 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8693
timestamp 1677677812
transform 1 0 1604 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8563
timestamp 1677677812
transform 1 0 1676 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9670
timestamp 1677677812
transform 1 0 1668 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8626
timestamp 1677677812
transform 1 0 1668 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9808
timestamp 1677677812
transform 1 0 1676 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8603
timestamp 1677677812
transform 1 0 1692 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9809
timestamp 1677677812
transform 1 0 1692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9671
timestamp 1677677812
transform 1 0 1700 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9672
timestamp 1677677812
transform 1 0 1708 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8654
timestamp 1677677812
transform 1 0 1708 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8564
timestamp 1677677812
transform 1 0 1732 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9673
timestamp 1677677812
transform 1 0 1732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9674
timestamp 1677677812
transform 1 0 1748 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9810
timestamp 1677677812
transform 1 0 1740 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8627
timestamp 1677677812
transform 1 0 1748 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_9811
timestamp 1677677812
transform 1 0 1756 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8565
timestamp 1677677812
transform 1 0 1772 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9675
timestamp 1677677812
transform 1 0 1764 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8505
timestamp 1677677812
transform 1 0 1804 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9676
timestamp 1677677812
transform 1 0 1788 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8604
timestamp 1677677812
transform 1 0 1796 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9677
timestamp 1677677812
transform 1 0 1804 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8605
timestamp 1677677812
transform 1 0 1812 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9812
timestamp 1677677812
transform 1 0 1780 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9813
timestamp 1677677812
transform 1 0 1796 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9814
timestamp 1677677812
transform 1 0 1804 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9815
timestamp 1677677812
transform 1 0 1828 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8694
timestamp 1677677812
transform 1 0 1828 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9678
timestamp 1677677812
transform 1 0 1844 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8506
timestamp 1677677812
transform 1 0 1876 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9679
timestamp 1677677812
transform 1 0 1860 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9680
timestamp 1677677812
transform 1 0 1876 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8628
timestamp 1677677812
transform 1 0 1860 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8530
timestamp 1677677812
transform 1 0 1908 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8566
timestamp 1677677812
transform 1 0 1900 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9681
timestamp 1677677812
transform 1 0 1908 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8655
timestamp 1677677812
transform 1 0 1900 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8606
timestamp 1677677812
transform 1 0 1916 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9816
timestamp 1677677812
transform 1 0 1916 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8531
timestamp 1677677812
transform 1 0 1932 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8567
timestamp 1677677812
transform 1 0 1932 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9817
timestamp 1677677812
transform 1 0 1932 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8507
timestamp 1677677812
transform 1 0 1956 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9818
timestamp 1677677812
transform 1 0 1948 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8656
timestamp 1677677812
transform 1 0 1948 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9682
timestamp 1677677812
transform 1 0 1956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9683
timestamp 1677677812
transform 1 0 1964 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8629
timestamp 1677677812
transform 1 0 1964 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8532
timestamp 1677677812
transform 1 0 1980 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8568
timestamp 1677677812
transform 1 0 1988 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9684
timestamp 1677677812
transform 1 0 1988 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8607
timestamp 1677677812
transform 1 0 1996 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9685
timestamp 1677677812
transform 1 0 2004 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9686
timestamp 1677677812
transform 1 0 2012 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9819
timestamp 1677677812
transform 1 0 1996 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8657
timestamp 1677677812
transform 1 0 1988 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8695
timestamp 1677677812
transform 1 0 2004 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8495
timestamp 1677677812
transform 1 0 2060 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9687
timestamp 1677677812
transform 1 0 2100 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9820
timestamp 1677677812
transform 1 0 2124 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8658
timestamp 1677677812
transform 1 0 2124 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8496
timestamp 1677677812
transform 1 0 2148 0 1 265
box -3 -3 3 3
use M2_M1  M2_M1_9688
timestamp 1677677812
transform 1 0 2148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9689
timestamp 1677677812
transform 1 0 2212 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9821
timestamp 1677677812
transform 1 0 2244 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8569
timestamp 1677677812
transform 1 0 2324 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9690
timestamp 1677677812
transform 1 0 2324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9822
timestamp 1677677812
transform 1 0 2276 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8696
timestamp 1677677812
transform 1 0 2340 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9691
timestamp 1677677812
transform 1 0 2372 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8570
timestamp 1677677812
transform 1 0 2412 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8571
timestamp 1677677812
transform 1 0 2460 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8533
timestamp 1677677812
transform 1 0 2476 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9692
timestamp 1677677812
transform 1 0 2412 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9693
timestamp 1677677812
transform 1 0 2468 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9823
timestamp 1677677812
transform 1 0 2388 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8608
timestamp 1677677812
transform 1 0 2484 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9694
timestamp 1677677812
transform 1 0 2492 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9824
timestamp 1677677812
transform 1 0 2476 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8534
timestamp 1677677812
transform 1 0 2524 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9601
timestamp 1677677812
transform 1 0 2516 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_8609
timestamp 1677677812
transform 1 0 2516 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9695
timestamp 1677677812
transform 1 0 2524 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9825
timestamp 1677677812
transform 1 0 2516 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8697
timestamp 1677677812
transform 1 0 2508 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8535
timestamp 1677677812
transform 1 0 2564 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9602
timestamp 1677677812
transform 1 0 2564 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9696
timestamp 1677677812
transform 1 0 2556 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9826
timestamp 1677677812
transform 1 0 2532 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9827
timestamp 1677677812
transform 1 0 2548 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8659
timestamp 1677677812
transform 1 0 2524 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8698
timestamp 1677677812
transform 1 0 2532 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8610
timestamp 1677677812
transform 1 0 2564 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9828
timestamp 1677677812
transform 1 0 2564 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8660
timestamp 1677677812
transform 1 0 2564 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8536
timestamp 1677677812
transform 1 0 2588 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9829
timestamp 1677677812
transform 1 0 2580 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8537
timestamp 1677677812
transform 1 0 2620 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8572
timestamp 1677677812
transform 1 0 2604 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9603
timestamp 1677677812
transform 1 0 2620 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9697
timestamp 1677677812
transform 1 0 2604 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9830
timestamp 1677677812
transform 1 0 2620 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8661
timestamp 1677677812
transform 1 0 2620 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8573
timestamp 1677677812
transform 1 0 2636 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9698
timestamp 1677677812
transform 1 0 2636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9699
timestamp 1677677812
transform 1 0 2652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9700
timestamp 1677677812
transform 1 0 2668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9831
timestamp 1677677812
transform 1 0 2628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8662
timestamp 1677677812
transform 1 0 2644 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8574
timestamp 1677677812
transform 1 0 2724 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9832
timestamp 1677677812
transform 1 0 2716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9833
timestamp 1677677812
transform 1 0 2724 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9604
timestamp 1677677812
transform 1 0 2748 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_8575
timestamp 1677677812
transform 1 0 2756 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9701
timestamp 1677677812
transform 1 0 2764 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9702
timestamp 1677677812
transform 1 0 2788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9703
timestamp 1677677812
transform 1 0 2804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9834
timestamp 1677677812
transform 1 0 2772 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9835
timestamp 1677677812
transform 1 0 2780 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9836
timestamp 1677677812
transform 1 0 2796 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8663
timestamp 1677677812
transform 1 0 2780 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8699
timestamp 1677677812
transform 1 0 2772 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9704
timestamp 1677677812
transform 1 0 2820 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8611
timestamp 1677677812
transform 1 0 2828 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_8664
timestamp 1677677812
transform 1 0 2820 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9837
timestamp 1677677812
transform 1 0 2836 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8612
timestamp 1677677812
transform 1 0 2852 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9838
timestamp 1677677812
transform 1 0 2852 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9839
timestamp 1677677812
transform 1 0 2868 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8538
timestamp 1677677812
transform 1 0 2924 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8576
timestamp 1677677812
transform 1 0 2916 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9705
timestamp 1677677812
transform 1 0 2916 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9706
timestamp 1677677812
transform 1 0 2932 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9707
timestamp 1677677812
transform 1 0 2940 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9840
timestamp 1677677812
transform 1 0 2908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9841
timestamp 1677677812
transform 1 0 2924 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8700
timestamp 1677677812
transform 1 0 2940 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8521
timestamp 1677677812
transform 1 0 3036 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_9708
timestamp 1677677812
transform 1 0 3044 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9842
timestamp 1677677812
transform 1 0 3068 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8665
timestamp 1677677812
transform 1 0 3068 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8522
timestamp 1677677812
transform 1 0 3084 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_8539
timestamp 1677677812
transform 1 0 3084 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9709
timestamp 1677677812
transform 1 0 3084 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8577
timestamp 1677677812
transform 1 0 3148 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9710
timestamp 1677677812
transform 1 0 3148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9843
timestamp 1677677812
transform 1 0 3172 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8666
timestamp 1677677812
transform 1 0 3172 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8667
timestamp 1677677812
transform 1 0 3188 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8578
timestamp 1677677812
transform 1 0 3260 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9711
timestamp 1677677812
transform 1 0 3260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9844
timestamp 1677677812
transform 1 0 3236 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8630
timestamp 1677677812
transform 1 0 3260 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_8668
timestamp 1677677812
transform 1 0 3236 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9845
timestamp 1677677812
transform 1 0 3332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9712
timestamp 1677677812
transform 1 0 3348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9846
timestamp 1677677812
transform 1 0 3348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9605
timestamp 1677677812
transform 1 0 3364 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_8613
timestamp 1677677812
transform 1 0 3380 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9606
timestamp 1677677812
transform 1 0 3404 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9713
timestamp 1677677812
transform 1 0 3388 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9714
timestamp 1677677812
transform 1 0 3396 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9847
timestamp 1677677812
transform 1 0 3380 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8540
timestamp 1677677812
transform 1 0 3420 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8614
timestamp 1677677812
transform 1 0 3412 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9848
timestamp 1677677812
transform 1 0 3412 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8669
timestamp 1677677812
transform 1 0 3412 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9607
timestamp 1677677812
transform 1 0 3436 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9849
timestamp 1677677812
transform 1 0 3436 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9608
timestamp 1677677812
transform 1 0 3452 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_9850
timestamp 1677677812
transform 1 0 3444 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8670
timestamp 1677677812
transform 1 0 3444 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8701
timestamp 1677677812
transform 1 0 3444 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8541
timestamp 1677677812
transform 1 0 3468 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9609
timestamp 1677677812
transform 1 0 3468 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_8579
timestamp 1677677812
transform 1 0 3476 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9715
timestamp 1677677812
transform 1 0 3476 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8580
timestamp 1677677812
transform 1 0 3524 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8581
timestamp 1677677812
transform 1 0 3540 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9716
timestamp 1677677812
transform 1 0 3540 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9851
timestamp 1677677812
transform 1 0 3492 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9717
timestamp 1677677812
transform 1 0 3580 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9718
timestamp 1677677812
transform 1 0 3588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9852
timestamp 1677677812
transform 1 0 3580 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8702
timestamp 1677677812
transform 1 0 3580 0 1 185
box -3 -3 3 3
use M2_M1  M2_M1_9719
timestamp 1677677812
transform 1 0 3604 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8542
timestamp 1677677812
transform 1 0 3636 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_9720
timestamp 1677677812
transform 1 0 3636 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9853
timestamp 1677677812
transform 1 0 3612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9854
timestamp 1677677812
transform 1 0 3628 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8582
timestamp 1677677812
transform 1 0 3652 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8543
timestamp 1677677812
transform 1 0 3676 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8583
timestamp 1677677812
transform 1 0 3668 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9855
timestamp 1677677812
transform 1 0 3668 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8671
timestamp 1677677812
transform 1 0 3684 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8508
timestamp 1677677812
transform 1 0 3708 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_8584
timestamp 1677677812
transform 1 0 3732 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9721
timestamp 1677677812
transform 1 0 3708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9722
timestamp 1677677812
transform 1 0 3724 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9723
timestamp 1677677812
transform 1 0 3732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9856
timestamp 1677677812
transform 1 0 3716 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9857
timestamp 1677677812
transform 1 0 3732 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8672
timestamp 1677677812
transform 1 0 3708 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8673
timestamp 1677677812
transform 1 0 3724 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8703
timestamp 1677677812
transform 1 0 3732 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8509
timestamp 1677677812
transform 1 0 3748 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9858
timestamp 1677677812
transform 1 0 3764 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8674
timestamp 1677677812
transform 1 0 3756 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9859
timestamp 1677677812
transform 1 0 3780 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9724
timestamp 1677677812
transform 1 0 3804 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9725
timestamp 1677677812
transform 1 0 3820 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9726
timestamp 1677677812
transform 1 0 3836 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9860
timestamp 1677677812
transform 1 0 3812 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9861
timestamp 1677677812
transform 1 0 3828 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8704
timestamp 1677677812
transform 1 0 3812 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8585
timestamp 1677677812
transform 1 0 3860 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8615
timestamp 1677677812
transform 1 0 3860 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9862
timestamp 1677677812
transform 1 0 3860 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9727
timestamp 1677677812
transform 1 0 3900 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9863
timestamp 1677677812
transform 1 0 3908 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9864
timestamp 1677677812
transform 1 0 3924 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8675
timestamp 1677677812
transform 1 0 3908 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8705
timestamp 1677677812
transform 1 0 3924 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8586
timestamp 1677677812
transform 1 0 3940 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9728
timestamp 1677677812
transform 1 0 3940 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8587
timestamp 1677677812
transform 1 0 4060 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9729
timestamp 1677677812
transform 1 0 3996 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9730
timestamp 1677677812
transform 1 0 4052 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9731
timestamp 1677677812
transform 1 0 4060 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9865
timestamp 1677677812
transform 1 0 3972 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8676
timestamp 1677677812
transform 1 0 3996 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8677
timestamp 1677677812
transform 1 0 4012 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8678
timestamp 1677677812
transform 1 0 4052 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8544
timestamp 1677677812
transform 1 0 4084 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8616
timestamp 1677677812
transform 1 0 4076 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9732
timestamp 1677677812
transform 1 0 4084 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9866
timestamp 1677677812
transform 1 0 4068 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9867
timestamp 1677677812
transform 1 0 4076 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9868
timestamp 1677677812
transform 1 0 4092 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9869
timestamp 1677677812
transform 1 0 4108 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8679
timestamp 1677677812
transform 1 0 4092 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8706
timestamp 1677677812
transform 1 0 4108 0 1 185
box -3 -3 3 3
use M3_M2  M3_M2_8588
timestamp 1677677812
transform 1 0 4124 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9733
timestamp 1677677812
transform 1 0 4124 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8589
timestamp 1677677812
transform 1 0 4228 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8617
timestamp 1677677812
transform 1 0 4140 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9734
timestamp 1677677812
transform 1 0 4164 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8618
timestamp 1677677812
transform 1 0 4204 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_9735
timestamp 1677677812
transform 1 0 4220 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9736
timestamp 1677677812
transform 1 0 4228 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9870
timestamp 1677677812
transform 1 0 4140 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8680
timestamp 1677677812
transform 1 0 4164 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8545
timestamp 1677677812
transform 1 0 4268 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_8590
timestamp 1677677812
transform 1 0 4252 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9737
timestamp 1677677812
transform 1 0 4252 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9738
timestamp 1677677812
transform 1 0 4268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9871
timestamp 1677677812
transform 1 0 4236 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9872
timestamp 1677677812
transform 1 0 4244 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9873
timestamp 1677677812
transform 1 0 4260 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8591
timestamp 1677677812
transform 1 0 4284 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9739
timestamp 1677677812
transform 1 0 4284 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9874
timestamp 1677677812
transform 1 0 4284 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9875
timestamp 1677677812
transform 1 0 4300 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9876
timestamp 1677677812
transform 1 0 4308 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8681
timestamp 1677677812
transform 1 0 4284 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8682
timestamp 1677677812
transform 1 0 4308 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9740
timestamp 1677677812
transform 1 0 4324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9741
timestamp 1677677812
transform 1 0 4348 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9877
timestamp 1677677812
transform 1 0 4332 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9878
timestamp 1677677812
transform 1 0 4348 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9879
timestamp 1677677812
transform 1 0 4396 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9880
timestamp 1677677812
transform 1 0 4404 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8683
timestamp 1677677812
transform 1 0 4404 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9742
timestamp 1677677812
transform 1 0 4436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9743
timestamp 1677677812
transform 1 0 4452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9881
timestamp 1677677812
transform 1 0 4444 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9882
timestamp 1677677812
transform 1 0 4460 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8684
timestamp 1677677812
transform 1 0 4476 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9883
timestamp 1677677812
transform 1 0 4508 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9884
timestamp 1677677812
transform 1 0 4516 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8685
timestamp 1677677812
transform 1 0 4516 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_8510
timestamp 1677677812
transform 1 0 4548 0 1 255
box -3 -3 3 3
use M2_M1  M2_M1_9744
timestamp 1677677812
transform 1 0 4548 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9745
timestamp 1677677812
transform 1 0 4564 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9746
timestamp 1677677812
transform 1 0 4588 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9885
timestamp 1677677812
transform 1 0 4556 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9886
timestamp 1677677812
transform 1 0 4572 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8686
timestamp 1677677812
transform 1 0 4588 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_9887
timestamp 1677677812
transform 1 0 4612 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9888
timestamp 1677677812
transform 1 0 4628 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9747
timestamp 1677677812
transform 1 0 4668 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9748
timestamp 1677677812
transform 1 0 4684 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_8592
timestamp 1677677812
transform 1 0 4708 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_8593
timestamp 1677677812
transform 1 0 4732 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_9749
timestamp 1677677812
transform 1 0 4732 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9750
timestamp 1677677812
transform 1 0 4788 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_9889
timestamp 1677677812
transform 1 0 4676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9890
timestamp 1677677812
transform 1 0 4692 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_9891
timestamp 1677677812
transform 1 0 4708 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_8631
timestamp 1677677812
transform 1 0 4780 0 1 205
box -3 -3 3 3
use top_level_VIA0  top_level_VIA0_90
timestamp 1677677812
transform 1 0 48 0 1 170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_599
timestamp 1677677812
transform 1 0 72 0 1 170
box -8 -3 104 105
use INVX2  INVX2_687
timestamp 1677677812
transform -1 0 184 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_398
timestamp 1677677812
transform -1 0 224 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_399
timestamp 1677677812
transform -1 0 264 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_400
timestamp 1677677812
transform 1 0 264 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_401
timestamp 1677677812
transform 1 0 304 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_402
timestamp 1677677812
transform 1 0 344 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_434
timestamp 1677677812
transform 1 0 384 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_435
timestamp 1677677812
transform 1 0 424 0 1 170
box -8 -3 46 105
use FILL  FILL_10549
timestamp 1677677812
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_10550
timestamp 1677677812
transform 1 0 472 0 1 170
box -8 -3 16 105
use INVX2  INVX2_688
timestamp 1677677812
transform 1 0 480 0 1 170
box -9 -3 26 105
use FILL  FILL_10551
timestamp 1677677812
transform 1 0 496 0 1 170
box -8 -3 16 105
use FILL  FILL_10552
timestamp 1677677812
transform 1 0 504 0 1 170
box -8 -3 16 105
use FILL  FILL_10553
timestamp 1677677812
transform 1 0 512 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8707
timestamp 1677677812
transform 1 0 532 0 1 175
box -3 -3 3 3
use FILL  FILL_10554
timestamp 1677677812
transform 1 0 520 0 1 170
box -8 -3 16 105
use FILL  FILL_10572
timestamp 1677677812
transform 1 0 528 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_403
timestamp 1677677812
transform 1 0 536 0 1 170
box -8 -3 46 105
use FILL  FILL_10574
timestamp 1677677812
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_10575
timestamp 1677677812
transform 1 0 584 0 1 170
box -8 -3 16 105
use FILL  FILL_10576
timestamp 1677677812
transform 1 0 592 0 1 170
box -8 -3 16 105
use FILL  FILL_10577
timestamp 1677677812
transform 1 0 600 0 1 170
box -8 -3 16 105
use FILL  FILL_10578
timestamp 1677677812
transform 1 0 608 0 1 170
box -8 -3 16 105
use FILL  FILL_10579
timestamp 1677677812
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_10580
timestamp 1677677812
transform 1 0 624 0 1 170
box -8 -3 16 105
use FILL  FILL_10581
timestamp 1677677812
transform 1 0 632 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_404
timestamp 1677677812
transform -1 0 680 0 1 170
box -8 -3 46 105
use FILL  FILL_10582
timestamp 1677677812
transform 1 0 680 0 1 170
box -8 -3 16 105
use INVX2  INVX2_691
timestamp 1677677812
transform 1 0 688 0 1 170
box -9 -3 26 105
use FILL  FILL_10583
timestamp 1677677812
transform 1 0 704 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_436
timestamp 1677677812
transform 1 0 712 0 1 170
box -8 -3 46 105
use M3_M2  M3_M2_8708
timestamp 1677677812
transform 1 0 772 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_437
timestamp 1677677812
transform 1 0 752 0 1 170
box -8 -3 46 105
use FILL  FILL_10584
timestamp 1677677812
transform 1 0 792 0 1 170
box -8 -3 16 105
use FILL  FILL_10585
timestamp 1677677812
transform 1 0 800 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_119
timestamp 1677677812
transform 1 0 808 0 1 170
box -8 -3 32 105
use FILL  FILL_10586
timestamp 1677677812
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_10594
timestamp 1677677812
transform 1 0 840 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_120
timestamp 1677677812
transform 1 0 848 0 1 170
box -8 -3 32 105
use FILL  FILL_10595
timestamp 1677677812
transform 1 0 872 0 1 170
box -8 -3 16 105
use FILL  FILL_10596
timestamp 1677677812
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_10597
timestamp 1677677812
transform 1 0 888 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_605
timestamp 1677677812
transform -1 0 992 0 1 170
box -8 -3 104 105
use INVX2  INVX2_693
timestamp 1677677812
transform -1 0 1008 0 1 170
box -9 -3 26 105
use AOI22X1  AOI22X1_406
timestamp 1677677812
transform -1 0 1048 0 1 170
box -8 -3 46 105
use FILL  FILL_10598
timestamp 1677677812
transform 1 0 1048 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_606
timestamp 1677677812
transform 1 0 1056 0 1 170
box -8 -3 104 105
use FILL  FILL_10599
timestamp 1677677812
transform 1 0 1152 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_407
timestamp 1677677812
transform 1 0 1160 0 1 170
box -8 -3 46 105
use OAI22X1  OAI22X1_438
timestamp 1677677812
transform -1 0 1240 0 1 170
box -8 -3 46 105
use FILL  FILL_10600
timestamp 1677677812
transform 1 0 1240 0 1 170
box -8 -3 16 105
use FILL  FILL_10601
timestamp 1677677812
transform 1 0 1248 0 1 170
box -8 -3 16 105
use FILL  FILL_10602
timestamp 1677677812
transform 1 0 1256 0 1 170
box -8 -3 16 105
use FILL  FILL_10603
timestamp 1677677812
transform 1 0 1264 0 1 170
box -8 -3 16 105
use FILL  FILL_10604
timestamp 1677677812
transform 1 0 1272 0 1 170
box -8 -3 16 105
use FILL  FILL_10610
timestamp 1677677812
transform 1 0 1280 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8709
timestamp 1677677812
transform 1 0 1348 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_8710
timestamp 1677677812
transform 1 0 1380 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_610
timestamp 1677677812
transform -1 0 1384 0 1 170
box -8 -3 104 105
use FILL  FILL_10611
timestamp 1677677812
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_10612
timestamp 1677677812
transform 1 0 1392 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_410
timestamp 1677677812
transform -1 0 1440 0 1 170
box -8 -3 46 105
use INVX2  INVX2_696
timestamp 1677677812
transform 1 0 1440 0 1 170
box -9 -3 26 105
use FILL  FILL_10613
timestamp 1677677812
transform 1 0 1456 0 1 170
box -8 -3 16 105
use FILL  FILL_10614
timestamp 1677677812
transform 1 0 1464 0 1 170
box -8 -3 16 105
use FILL  FILL_10615
timestamp 1677677812
transform 1 0 1472 0 1 170
box -8 -3 16 105
use FILL  FILL_10616
timestamp 1677677812
transform 1 0 1480 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_411
timestamp 1677677812
transform -1 0 1528 0 1 170
box -8 -3 46 105
use FILL  FILL_10617
timestamp 1677677812
transform 1 0 1528 0 1 170
box -8 -3 16 105
use FILL  FILL_10618
timestamp 1677677812
transform 1 0 1536 0 1 170
box -8 -3 16 105
use FILL  FILL_10619
timestamp 1677677812
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_10620
timestamp 1677677812
transform 1 0 1552 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_439
timestamp 1677677812
transform -1 0 1600 0 1 170
box -8 -3 46 105
use AOI22X1  AOI22X1_412
timestamp 1677677812
transform 1 0 1600 0 1 170
box -8 -3 46 105
use FILL  FILL_10621
timestamp 1677677812
transform 1 0 1640 0 1 170
box -8 -3 16 105
use FILL  FILL_10628
timestamp 1677677812
transform 1 0 1648 0 1 170
box -8 -3 16 105
use FILL  FILL_10630
timestamp 1677677812
transform 1 0 1656 0 1 170
box -8 -3 16 105
use FILL  FILL_10632
timestamp 1677677812
transform 1 0 1664 0 1 170
box -8 -3 16 105
use INVX2  INVX2_699
timestamp 1677677812
transform 1 0 1672 0 1 170
box -9 -3 26 105
use FILL  FILL_10633
timestamp 1677677812
transform 1 0 1688 0 1 170
box -8 -3 16 105
use FILL  FILL_10634
timestamp 1677677812
transform 1 0 1696 0 1 170
box -8 -3 16 105
use FILL  FILL_10635
timestamp 1677677812
transform 1 0 1704 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_413
timestamp 1677677812
transform 1 0 1712 0 1 170
box -8 -3 46 105
use FILL  FILL_10636
timestamp 1677677812
transform 1 0 1752 0 1 170
box -8 -3 16 105
use FILL  FILL_10637
timestamp 1677677812
transform 1 0 1760 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_414
timestamp 1677677812
transform -1 0 1808 0 1 170
box -8 -3 46 105
use INVX2  INVX2_700
timestamp 1677677812
transform 1 0 1808 0 1 170
box -9 -3 26 105
use FILL  FILL_10638
timestamp 1677677812
transform 1 0 1824 0 1 170
box -8 -3 16 105
use FILL  FILL_10639
timestamp 1677677812
transform 1 0 1832 0 1 170
box -8 -3 16 105
use FILL  FILL_10640
timestamp 1677677812
transform 1 0 1840 0 1 170
box -8 -3 16 105
use FILL  FILL_10641
timestamp 1677677812
transform 1 0 1848 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_415
timestamp 1677677812
transform -1 0 1896 0 1 170
box -8 -3 46 105
use FILL  FILL_10642
timestamp 1677677812
transform 1 0 1896 0 1 170
box -8 -3 16 105
use FILL  FILL_10643
timestamp 1677677812
transform 1 0 1904 0 1 170
box -8 -3 16 105
use FILL  FILL_10644
timestamp 1677677812
transform 1 0 1912 0 1 170
box -8 -3 16 105
use FILL  FILL_10645
timestamp 1677677812
transform 1 0 1920 0 1 170
box -8 -3 16 105
use INVX2  INVX2_701
timestamp 1677677812
transform 1 0 1928 0 1 170
box -9 -3 26 105
use FILL  FILL_10646
timestamp 1677677812
transform 1 0 1944 0 1 170
box -8 -3 16 105
use FILL  FILL_10647
timestamp 1677677812
transform 1 0 1952 0 1 170
box -8 -3 16 105
use FILL  FILL_10648
timestamp 1677677812
transform 1 0 1960 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_416
timestamp 1677677812
transform -1 0 2008 0 1 170
box -8 -3 46 105
use FILL  FILL_10649
timestamp 1677677812
transform 1 0 2008 0 1 170
box -8 -3 16 105
use FILL  FILL_10650
timestamp 1677677812
transform 1 0 2016 0 1 170
box -8 -3 16 105
use FILL  FILL_10651
timestamp 1677677812
transform 1 0 2024 0 1 170
box -8 -3 16 105
use FILL  FILL_10652
timestamp 1677677812
transform 1 0 2032 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8711
timestamp 1677677812
transform 1 0 2068 0 1 175
box -3 -3 3 3
use M3_M2  M3_M2_8712
timestamp 1677677812
transform 1 0 2084 0 1 175
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_614
timestamp 1677677812
transform -1 0 2136 0 1 170
box -8 -3 104 105
use FILL  FILL_10653
timestamp 1677677812
transform 1 0 2136 0 1 170
box -8 -3 16 105
use FILL  FILL_10654
timestamp 1677677812
transform 1 0 2144 0 1 170
box -8 -3 16 105
use FILL  FILL_10655
timestamp 1677677812
transform 1 0 2152 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_615
timestamp 1677677812
transform -1 0 2256 0 1 170
box -8 -3 104 105
use FILL  FILL_10656
timestamp 1677677812
transform 1 0 2256 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_616
timestamp 1677677812
transform 1 0 2264 0 1 170
box -8 -3 104 105
use FILL  FILL_10657
timestamp 1677677812
transform 1 0 2360 0 1 170
box -8 -3 16 105
use FILL  FILL_10658
timestamp 1677677812
transform 1 0 2368 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_617
timestamp 1677677812
transform 1 0 2376 0 1 170
box -8 -3 104 105
use FILL  FILL_10659
timestamp 1677677812
transform 1 0 2472 0 1 170
box -8 -3 16 105
use FILL  FILL_10660
timestamp 1677677812
transform 1 0 2480 0 1 170
box -8 -3 16 105
use FILL  FILL_10678
timestamp 1677677812
transform 1 0 2488 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_53
timestamp 1677677812
transform 1 0 2496 0 1 170
box -8 -3 32 105
use FILL  FILL_10679
timestamp 1677677812
transform 1 0 2520 0 1 170
box -8 -3 16 105
use INVX2  INVX2_703
timestamp 1677677812
transform 1 0 2528 0 1 170
box -9 -3 26 105
use NAND2X1  NAND2X1_54
timestamp 1677677812
transform 1 0 2544 0 1 170
box -8 -3 32 105
use FILL  FILL_10680
timestamp 1677677812
transform 1 0 2568 0 1 170
box -8 -3 16 105
use FILL  FILL_10681
timestamp 1677677812
transform 1 0 2576 0 1 170
box -8 -3 16 105
use FILL  FILL_10682
timestamp 1677677812
transform 1 0 2584 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_183
timestamp 1677677812
transform 1 0 2592 0 1 170
box -8 -3 34 105
use FILL  FILL_10683
timestamp 1677677812
transform 1 0 2624 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_417
timestamp 1677677812
transform 1 0 2632 0 1 170
box -8 -3 46 105
use FILL  FILL_10684
timestamp 1677677812
transform 1 0 2672 0 1 170
box -8 -3 16 105
use FILL  FILL_10685
timestamp 1677677812
transform 1 0 2680 0 1 170
box -8 -3 16 105
use FILL  FILL_10686
timestamp 1677677812
transform 1 0 2688 0 1 170
box -8 -3 16 105
use FILL  FILL_10687
timestamp 1677677812
transform 1 0 2696 0 1 170
box -8 -3 16 105
use INVX2  INVX2_704
timestamp 1677677812
transform -1 0 2720 0 1 170
box -9 -3 26 105
use FILL  FILL_10688
timestamp 1677677812
transform 1 0 2720 0 1 170
box -8 -3 16 105
use FILL  FILL_10689
timestamp 1677677812
transform 1 0 2728 0 1 170
box -8 -3 16 105
use FILL  FILL_10690
timestamp 1677677812
transform 1 0 2736 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_184
timestamp 1677677812
transform -1 0 2776 0 1 170
box -8 -3 34 105
use OAI22X1  OAI22X1_440
timestamp 1677677812
transform 1 0 2776 0 1 170
box -8 -3 46 105
use FILL  FILL_10691
timestamp 1677677812
transform 1 0 2816 0 1 170
box -8 -3 16 105
use FILL  FILL_10702
timestamp 1677677812
transform 1 0 2824 0 1 170
box -8 -3 16 105
use FILL  FILL_10704
timestamp 1677677812
transform 1 0 2832 0 1 170
box -8 -3 16 105
use INVX2  INVX2_706
timestamp 1677677812
transform -1 0 2856 0 1 170
box -9 -3 26 105
use FILL  FILL_10705
timestamp 1677677812
transform 1 0 2856 0 1 170
box -8 -3 16 105
use FILL  FILL_10706
timestamp 1677677812
transform 1 0 2864 0 1 170
box -8 -3 16 105
use FILL  FILL_10707
timestamp 1677677812
transform 1 0 2872 0 1 170
box -8 -3 16 105
use FILL  FILL_10708
timestamp 1677677812
transform 1 0 2880 0 1 170
box -8 -3 16 105
use FILL  FILL_10709
timestamp 1677677812
transform 1 0 2888 0 1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_418
timestamp 1677677812
transform 1 0 2896 0 1 170
box -8 -3 46 105
use FILL  FILL_10710
timestamp 1677677812
transform 1 0 2936 0 1 170
box -8 -3 16 105
use FILL  FILL_10716
timestamp 1677677812
transform 1 0 2944 0 1 170
box -8 -3 16 105
use FILL  FILL_10717
timestamp 1677677812
transform 1 0 2952 0 1 170
box -8 -3 16 105
use FILL  FILL_10718
timestamp 1677677812
transform 1 0 2960 0 1 170
box -8 -3 16 105
use INVX2  INVX2_709
timestamp 1677677812
transform -1 0 2984 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_627
timestamp 1677677812
transform -1 0 3080 0 1 170
box -8 -3 104 105
use FILL  FILL_10719
timestamp 1677677812
transform 1 0 3080 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_628
timestamp 1677677812
transform -1 0 3184 0 1 170
box -8 -3 104 105
use FILL  FILL_10720
timestamp 1677677812
transform 1 0 3184 0 1 170
box -8 -3 16 105
use FILL  FILL_10721
timestamp 1677677812
transform 1 0 3192 0 1 170
box -8 -3 16 105
use FILL  FILL_10722
timestamp 1677677812
transform 1 0 3200 0 1 170
box -8 -3 16 105
use FILL  FILL_10732
timestamp 1677677812
transform 1 0 3208 0 1 170
box -8 -3 16 105
use FILL  FILL_10734
timestamp 1677677812
transform 1 0 3216 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_631
timestamp 1677677812
transform 1 0 3224 0 1 170
box -8 -3 104 105
use FILL  FILL_10736
timestamp 1677677812
transform 1 0 3320 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_56
timestamp 1677677812
transform 1 0 3328 0 1 170
box -8 -3 32 105
use FILL  FILL_10738
timestamp 1677677812
transform 1 0 3352 0 1 170
box -8 -3 16 105
use FILL  FILL_10741
timestamp 1677677812
transform 1 0 3360 0 1 170
box -8 -3 16 105
use FILL  FILL_10743
timestamp 1677677812
transform 1 0 3368 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_57
timestamp 1677677812
transform 1 0 3376 0 1 170
box -8 -3 32 105
use FILL  FILL_10744
timestamp 1677677812
transform 1 0 3400 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8713
timestamp 1677677812
transform 1 0 3436 0 1 175
box -3 -3 3 3
use OAI21X1  OAI21X1_185
timestamp 1677677812
transform 1 0 3408 0 1 170
box -8 -3 34 105
use FILL  FILL_10745
timestamp 1677677812
transform 1 0 3440 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_58
timestamp 1677677812
transform 1 0 3448 0 1 170
box -8 -3 32 105
use FILL  FILL_10746
timestamp 1677677812
transform 1 0 3472 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_633
timestamp 1677677812
transform 1 0 3480 0 1 170
box -8 -3 104 105
use FILL  FILL_10747
timestamp 1677677812
transform 1 0 3576 0 1 170
box -8 -3 16 105
use FILL  FILL_10748
timestamp 1677677812
transform 1 0 3584 0 1 170
box -8 -3 16 105
use FILL  FILL_10753
timestamp 1677677812
transform 1 0 3592 0 1 170
box -8 -3 16 105
use FILL  FILL_10755
timestamp 1677677812
transform 1 0 3600 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_442
timestamp 1677677812
transform 1 0 3608 0 1 170
box -8 -3 46 105
use FILL  FILL_10757
timestamp 1677677812
transform 1 0 3648 0 1 170
box -8 -3 16 105
use FILL  FILL_10758
timestamp 1677677812
transform 1 0 3656 0 1 170
box -8 -3 16 105
use FILL  FILL_10759
timestamp 1677677812
transform 1 0 3664 0 1 170
box -8 -3 16 105
use FILL  FILL_10760
timestamp 1677677812
transform 1 0 3672 0 1 170
box -8 -3 16 105
use FILL  FILL_10761
timestamp 1677677812
transform 1 0 3680 0 1 170
box -8 -3 16 105
use FILL  FILL_10762
timestamp 1677677812
transform 1 0 3688 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_443
timestamp 1677677812
transform -1 0 3736 0 1 170
box -8 -3 46 105
use FILL  FILL_10763
timestamp 1677677812
transform 1 0 3736 0 1 170
box -8 -3 16 105
use FILL  FILL_10769
timestamp 1677677812
transform 1 0 3744 0 1 170
box -8 -3 16 105
use FILL  FILL_10770
timestamp 1677677812
transform 1 0 3752 0 1 170
box -8 -3 16 105
use INVX2  INVX2_712
timestamp 1677677812
transform 1 0 3760 0 1 170
box -9 -3 26 105
use FILL  FILL_10771
timestamp 1677677812
transform 1 0 3776 0 1 170
box -8 -3 16 105
use FILL  FILL_10772
timestamp 1677677812
transform 1 0 3784 0 1 170
box -8 -3 16 105
use FILL  FILL_10773
timestamp 1677677812
transform 1 0 3792 0 1 170
box -8 -3 16 105
use FILL  FILL_10774
timestamp 1677677812
transform 1 0 3800 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_444
timestamp 1677677812
transform 1 0 3808 0 1 170
box -8 -3 46 105
use FILL  FILL_10775
timestamp 1677677812
transform 1 0 3848 0 1 170
box -8 -3 16 105
use FILL  FILL_10776
timestamp 1677677812
transform 1 0 3856 0 1 170
box -8 -3 16 105
use FILL  FILL_10777
timestamp 1677677812
transform 1 0 3864 0 1 170
box -8 -3 16 105
use FILL  FILL_10778
timestamp 1677677812
transform 1 0 3872 0 1 170
box -8 -3 16 105
use FILL  FILL_10779
timestamp 1677677812
transform 1 0 3880 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_445
timestamp 1677677812
transform -1 0 3928 0 1 170
box -8 -3 46 105
use FILL  FILL_10780
timestamp 1677677812
transform 1 0 3928 0 1 170
box -8 -3 16 105
use FILL  FILL_10781
timestamp 1677677812
transform 1 0 3936 0 1 170
box -8 -3 16 105
use FILL  FILL_10782
timestamp 1677677812
transform 1 0 3944 0 1 170
box -8 -3 16 105
use FILL  FILL_10783
timestamp 1677677812
transform 1 0 3952 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_636
timestamp 1677677812
transform 1 0 3960 0 1 170
box -8 -3 104 105
use INVX2  INVX2_713
timestamp 1677677812
transform -1 0 4072 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_446
timestamp 1677677812
transform -1 0 4112 0 1 170
box -8 -3 46 105
use FILL  FILL_10784
timestamp 1677677812
transform 1 0 4112 0 1 170
box -8 -3 16 105
use FILL  FILL_10785
timestamp 1677677812
transform 1 0 4120 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_637
timestamp 1677677812
transform 1 0 4128 0 1 170
box -8 -3 104 105
use M3_M2  M3_M2_8714
timestamp 1677677812
transform 1 0 4244 0 1 175
box -3 -3 3 3
use INVX2  INVX2_714
timestamp 1677677812
transform -1 0 4240 0 1 170
box -9 -3 26 105
use OAI22X1  OAI22X1_447
timestamp 1677677812
transform 1 0 4240 0 1 170
box -8 -3 46 105
use FILL  FILL_10786
timestamp 1677677812
transform 1 0 4280 0 1 170
box -8 -3 16 105
use INVX2  INVX2_715
timestamp 1677677812
transform -1 0 4304 0 1 170
box -9 -3 26 105
use FILL  FILL_10787
timestamp 1677677812
transform 1 0 4304 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8715
timestamp 1677677812
transform 1 0 4348 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_448
timestamp 1677677812
transform -1 0 4352 0 1 170
box -8 -3 46 105
use INVX2  INVX2_716
timestamp 1677677812
transform -1 0 4368 0 1 170
box -9 -3 26 105
use FILL  FILL_10788
timestamp 1677677812
transform 1 0 4368 0 1 170
box -8 -3 16 105
use FILL  FILL_10789
timestamp 1677677812
transform 1 0 4376 0 1 170
box -8 -3 16 105
use FILL  FILL_10790
timestamp 1677677812
transform 1 0 4384 0 1 170
box -8 -3 16 105
use FILL  FILL_10791
timestamp 1677677812
transform 1 0 4392 0 1 170
box -8 -3 16 105
use FILL  FILL_10792
timestamp 1677677812
transform 1 0 4400 0 1 170
box -8 -3 16 105
use FILL  FILL_10808
timestamp 1677677812
transform 1 0 4408 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8716
timestamp 1677677812
transform 1 0 4428 0 1 175
box -3 -3 3 3
use FILL  FILL_10810
timestamp 1677677812
transform 1 0 4416 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8717
timestamp 1677677812
transform 1 0 4460 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_449
timestamp 1677677812
transform -1 0 4464 0 1 170
box -8 -3 46 105
use INVX2  INVX2_721
timestamp 1677677812
transform -1 0 4480 0 1 170
box -9 -3 26 105
use FILL  FILL_10811
timestamp 1677677812
transform 1 0 4480 0 1 170
box -8 -3 16 105
use FILL  FILL_10812
timestamp 1677677812
transform 1 0 4488 0 1 170
box -8 -3 16 105
use FILL  FILL_10813
timestamp 1677677812
transform 1 0 4496 0 1 170
box -8 -3 16 105
use FILL  FILL_10814
timestamp 1677677812
transform 1 0 4504 0 1 170
box -8 -3 16 105
use FILL  FILL_10815
timestamp 1677677812
transform 1 0 4512 0 1 170
box -8 -3 16 105
use FILL  FILL_10817
timestamp 1677677812
transform 1 0 4520 0 1 170
box -8 -3 16 105
use FILL  FILL_10818
timestamp 1677677812
transform 1 0 4528 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8718
timestamp 1677677812
transform 1 0 4572 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_450
timestamp 1677677812
transform -1 0 4576 0 1 170
box -8 -3 46 105
use INVX2  INVX2_722
timestamp 1677677812
transform -1 0 4592 0 1 170
box -9 -3 26 105
use FILL  FILL_10819
timestamp 1677677812
transform 1 0 4592 0 1 170
box -8 -3 16 105
use FILL  FILL_10820
timestamp 1677677812
transform 1 0 4600 0 1 170
box -8 -3 16 105
use FILL  FILL_10821
timestamp 1677677812
transform 1 0 4608 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8719
timestamp 1677677812
transform 1 0 4628 0 1 175
box -3 -3 3 3
use INVX2  INVX2_723
timestamp 1677677812
transform -1 0 4632 0 1 170
box -9 -3 26 105
use FILL  FILL_10822
timestamp 1677677812
transform 1 0 4632 0 1 170
box -8 -3 16 105
use FILL  FILL_10823
timestamp 1677677812
transform 1 0 4640 0 1 170
box -8 -3 16 105
use FILL  FILL_10824
timestamp 1677677812
transform 1 0 4648 0 1 170
box -8 -3 16 105
use M3_M2  M3_M2_8720
timestamp 1677677812
transform 1 0 4692 0 1 175
box -3 -3 3 3
use OAI22X1  OAI22X1_451
timestamp 1677677812
transform -1 0 4696 0 1 170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_644
timestamp 1677677812
transform 1 0 4696 0 1 170
box -8 -3 104 105
use top_level_VIA0  top_level_VIA0_91
timestamp 1677677812
transform 1 0 4819 0 1 170
box -10 -3 10 3
use top_level_VIA0  top_level_VIA0_92
timestamp 1677677812
transform 1 0 24 0 1 70
box -10 -3 10 3
use FILL  FILL_10555
timestamp 1677677812
transform 1 0 72 0 -1 170
box -8 -3 16 105
use FILL  FILL_10556
timestamp 1677677812
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_10557
timestamp 1677677812
transform 1 0 88 0 -1 170
box -8 -3 16 105
use FILL  FILL_10558
timestamp 1677677812
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_10559
timestamp 1677677812
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_10560
timestamp 1677677812
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_10561
timestamp 1677677812
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_10562
timestamp 1677677812
transform 1 0 128 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9895
timestamp 1677677812
transform 1 0 148 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9896
timestamp 1677677812
transform 1 0 244 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9957
timestamp 1677677812
transform 1 0 196 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9958
timestamp 1677677812
transform 1 0 228 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9959
timestamp 1677677812
transform 1 0 236 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8791
timestamp 1677677812
transform 1 0 196 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8792
timestamp 1677677812
transform 1 0 236 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_600
timestamp 1677677812
transform 1 0 136 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_689
timestamp 1677677812
transform -1 0 248 0 -1 170
box -9 -3 26 105
use FILL  FILL_10563
timestamp 1677677812
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_10564
timestamp 1677677812
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_10565
timestamp 1677677812
transform 1 0 264 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9897
timestamp 1677677812
transform 1 0 284 0 1 135
box -2 -2 2 2
use FILL  FILL_10566
timestamp 1677677812
transform 1 0 272 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9960
timestamp 1677677812
transform 1 0 300 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8793
timestamp 1677677812
transform 1 0 300 0 1 115
box -3 -3 3 3
use INVX2  INVX2_690
timestamp 1677677812
transform 1 0 280 0 -1 170
box -9 -3 26 105
use FILL  FILL_10567
timestamp 1677677812
transform 1 0 296 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8734
timestamp 1677677812
transform 1 0 316 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9898
timestamp 1677677812
transform 1 0 316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9961
timestamp 1677677812
transform 1 0 340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9962
timestamp 1677677812
transform 1 0 396 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8794
timestamp 1677677812
transform 1 0 340 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_601
timestamp 1677677812
transform 1 0 304 0 -1 170
box -8 -3 104 105
use FILL  FILL_10568
timestamp 1677677812
transform 1 0 400 0 -1 170
box -8 -3 16 105
use FILL  FILL_10569
timestamp 1677677812
transform 1 0 408 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8735
timestamp 1677677812
transform 1 0 508 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9899
timestamp 1677677812
transform 1 0 508 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9963
timestamp 1677677812
transform 1 0 428 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9964
timestamp 1677677812
transform 1 0 476 0 1 125
box -2 -2 2 2
use FILL  FILL_10570
timestamp 1677677812
transform 1 0 416 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_602
timestamp 1677677812
transform -1 0 520 0 -1 170
box -8 -3 104 105
use FILL  FILL_10571
timestamp 1677677812
transform 1 0 520 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9900
timestamp 1677677812
transform 1 0 540 0 1 135
box -2 -2 2 2
use FILL  FILL_10573
timestamp 1677677812
transform 1 0 528 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9965
timestamp 1677677812
transform 1 0 556 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8795
timestamp 1677677812
transform 1 0 556 0 1 115
box -3 -3 3 3
use INVX2  INVX2_692
timestamp 1677677812
transform 1 0 536 0 -1 170
box -9 -3 26 105
use FILL  FILL_10587
timestamp 1677677812
transform 1 0 552 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8736
timestamp 1677677812
transform 1 0 572 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9901
timestamp 1677677812
transform 1 0 572 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9966
timestamp 1677677812
transform 1 0 596 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9967
timestamp 1677677812
transform 1 0 652 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8796
timestamp 1677677812
transform 1 0 596 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_603
timestamp 1677677812
transform 1 0 560 0 -1 170
box -8 -3 104 105
use FILL  FILL_10588
timestamp 1677677812
transform 1 0 656 0 -1 170
box -8 -3 16 105
use FILL  FILL_10589
timestamp 1677677812
transform 1 0 664 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8737
timestamp 1677677812
transform 1 0 684 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9902
timestamp 1677677812
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9968
timestamp 1677677812
transform 1 0 708 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9969
timestamp 1677677812
transform 1 0 764 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9970
timestamp 1677677812
transform 1 0 772 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8797
timestamp 1677677812
transform 1 0 748 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_604
timestamp 1677677812
transform 1 0 672 0 -1 170
box -8 -3 104 105
use FILL  FILL_10590
timestamp 1677677812
transform 1 0 768 0 -1 170
box -8 -3 16 105
use FILL  FILL_10591
timestamp 1677677812
transform 1 0 776 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8738
timestamp 1677677812
transform 1 0 804 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9903
timestamp 1677677812
transform 1 0 804 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9904
timestamp 1677677812
transform 1 0 820 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9905
timestamp 1677677812
transform 1 0 828 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9971
timestamp 1677677812
transform 1 0 796 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9972
timestamp 1677677812
transform 1 0 812 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8798
timestamp 1677677812
transform 1 0 820 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8839
timestamp 1677677812
transform 1 0 796 0 1 95
box -3 -3 3 3
use FILL  FILL_10592
timestamp 1677677812
transform 1 0 784 0 -1 170
box -8 -3 16 105
use AOI22X1  AOI22X1_405
timestamp 1677677812
transform 1 0 792 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_8739
timestamp 1677677812
transform 1 0 844 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8774
timestamp 1677677812
transform 1 0 844 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8740
timestamp 1677677812
transform 1 0 940 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8775
timestamp 1677677812
transform 1 0 900 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9906
timestamp 1677677812
transform 1 0 940 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9973
timestamp 1677677812
transform 1 0 844 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9974
timestamp 1677677812
transform 1 0 852 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9975
timestamp 1677677812
transform 1 0 860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9976
timestamp 1677677812
transform 1 0 892 0 1 125
box -2 -2 2 2
use FILL  FILL_10593
timestamp 1677677812
transform 1 0 832 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8799
timestamp 1677677812
transform 1 0 852 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8800
timestamp 1677677812
transform 1 0 892 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8829
timestamp 1677677812
transform 1 0 860 0 1 105
box -3 -3 3 3
use INVX2  INVX2_694
timestamp 1677677812
transform 1 0 840 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_607
timestamp 1677677812
transform -1 0 952 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8741
timestamp 1677677812
transform 1 0 964 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8742
timestamp 1677677812
transform 1 0 980 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9907
timestamp 1677677812
transform 1 0 964 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8743
timestamp 1677677812
transform 1 0 1140 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9908
timestamp 1677677812
transform 1 0 1060 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8744
timestamp 1677677812
transform 1 0 1188 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9909
timestamp 1677677812
transform 1 0 1164 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9910
timestamp 1677677812
transform 1 0 1172 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9911
timestamp 1677677812
transform 1 0 1188 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9977
timestamp 1677677812
transform 1 0 996 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9978
timestamp 1677677812
transform 1 0 1044 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9979
timestamp 1677677812
transform 1 0 1108 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9980
timestamp 1677677812
transform 1 0 1140 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9981
timestamp 1677677812
transform 1 0 1148 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_608
timestamp 1677677812
transform 1 0 952 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8784
timestamp 1677677812
transform 1 0 1156 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9982
timestamp 1677677812
transform 1 0 1164 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8785
timestamp 1677677812
transform 1 0 1172 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_9983
timestamp 1677677812
transform 1 0 1180 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8801
timestamp 1677677812
transform 1 0 1108 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8802
timestamp 1677677812
transform 1 0 1148 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_609
timestamp 1677677812
transform 1 0 1048 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8840
timestamp 1677677812
transform 1 0 1164 0 1 95
box -3 -3 3 3
use INVX2  INVX2_695
timestamp 1677677812
transform -1 0 1160 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_9984
timestamp 1677677812
transform 1 0 1204 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8803
timestamp 1677677812
transform 1 0 1204 0 1 115
box -3 -3 3 3
use AOI22X1  AOI22X1_408
timestamp 1677677812
transform 1 0 1160 0 -1 170
box -8 -3 46 105
use FILL  FILL_10605
timestamp 1677677812
transform 1 0 1200 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9912
timestamp 1677677812
transform 1 0 1220 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8786
timestamp 1677677812
transform 1 0 1220 0 1 125
box -3 -3 3 3
use FILL  FILL_10606
timestamp 1677677812
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use FILL  FILL_10607
timestamp 1677677812
transform 1 0 1216 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9913
timestamp 1677677812
transform 1 0 1260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9914
timestamp 1677677812
transform 1 0 1268 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9985
timestamp 1677677812
transform 1 0 1236 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9986
timestamp 1677677812
transform 1 0 1252 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9987
timestamp 1677677812
transform 1 0 1268 0 1 125
box -2 -2 2 2
use FILL  FILL_10608
timestamp 1677677812
transform 1 0 1224 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8804
timestamp 1677677812
transform 1 0 1268 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8830
timestamp 1677677812
transform 1 0 1260 0 1 105
box -3 -3 3 3
use M2_M1  M2_M1_9915
timestamp 1677677812
transform 1 0 1380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9988
timestamp 1677677812
transform 1 0 1292 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9989
timestamp 1677677812
transform 1 0 1300 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9990
timestamp 1677677812
transform 1 0 1332 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8805
timestamp 1677677812
transform 1 0 1292 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8806
timestamp 1677677812
transform 1 0 1332 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8831
timestamp 1677677812
transform 1 0 1276 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_8832
timestamp 1677677812
transform 1 0 1300 0 1 105
box -3 -3 3 3
use AOI22X1  AOI22X1_409
timestamp 1677677812
transform 1 0 1232 0 -1 170
box -8 -3 46 105
use FILL  FILL_10609
timestamp 1677677812
transform 1 0 1272 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_697
timestamp 1677677812
transform 1 0 1280 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_611
timestamp 1677677812
transform -1 0 1392 0 -1 170
box -8 -3 104 105
use FILL  FILL_10622
timestamp 1677677812
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9916
timestamp 1677677812
transform 1 0 1492 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9991
timestamp 1677677812
transform 1 0 1412 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9992
timestamp 1677677812
transform 1 0 1460 0 1 125
box -2 -2 2 2
use FILL  FILL_10623
timestamp 1677677812
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_612
timestamp 1677677812
transform -1 0 1504 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8745
timestamp 1677677812
transform 1 0 1604 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9917
timestamp 1677677812
transform 1 0 1604 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9918
timestamp 1677677812
transform 1 0 1620 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9993
timestamp 1677677812
transform 1 0 1524 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9994
timestamp 1677677812
transform 1 0 1580 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9995
timestamp 1677677812
transform 1 0 1620 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8841
timestamp 1677677812
transform 1 0 1516 0 1 95
box -3 -3 3 3
use FILL  FILL_10624
timestamp 1677677812
transform 1 0 1504 0 -1 170
box -8 -3 16 105
use FILL  FILL_10625
timestamp 1677677812
transform 1 0 1512 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8807
timestamp 1677677812
transform 1 0 1580 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8808
timestamp 1677677812
transform 1 0 1620 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_613
timestamp 1677677812
transform -1 0 1616 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_698
timestamp 1677677812
transform 1 0 1616 0 -1 170
box -9 -3 26 105
use FILL  FILL_10626
timestamp 1677677812
transform 1 0 1632 0 -1 170
box -8 -3 16 105
use FILL  FILL_10627
timestamp 1677677812
transform 1 0 1640 0 -1 170
box -8 -3 16 105
use FILL  FILL_10629
timestamp 1677677812
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_10631
timestamp 1677677812
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8746
timestamp 1677677812
transform 1 0 1676 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9919
timestamp 1677677812
transform 1 0 1676 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9996
timestamp 1677677812
transform 1 0 1700 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9997
timestamp 1677677812
transform 1 0 1756 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_618
timestamp 1677677812
transform 1 0 1664 0 -1 170
box -8 -3 104 105
use FILL  FILL_10661
timestamp 1677677812
transform 1 0 1760 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9998
timestamp 1677677812
transform 1 0 1780 0 1 125
box -2 -2 2 2
use FILL  FILL_10662
timestamp 1677677812
transform 1 0 1768 0 -1 170
box -8 -3 16 105
use FILL  FILL_10663
timestamp 1677677812
transform 1 0 1776 0 -1 170
box -8 -3 16 105
use FILL  FILL_10664
timestamp 1677677812
transform 1 0 1784 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8747
timestamp 1677677812
transform 1 0 1876 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9920
timestamp 1677677812
transform 1 0 1876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9999
timestamp 1677677812
transform 1 0 1844 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_619
timestamp 1677677812
transform -1 0 1888 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8721
timestamp 1677677812
transform 1 0 1908 0 1 165
box -3 -3 3 3
use M2_M1  M2_M1_10000
timestamp 1677677812
transform 1 0 1900 0 1 125
box -2 -2 2 2
use FILL  FILL_10665
timestamp 1677677812
transform 1 0 1888 0 -1 170
box -8 -3 16 105
use FILL  FILL_10666
timestamp 1677677812
transform 1 0 1896 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9921
timestamp 1677677812
transform 1 0 1988 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10001
timestamp 1677677812
transform 1 0 1956 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8787
timestamp 1677677812
transform 1 0 1988 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_8809
timestamp 1677677812
transform 1 0 2004 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_620
timestamp 1677677812
transform -1 0 2000 0 -1 170
box -8 -3 104 105
use FILL  FILL_10667
timestamp 1677677812
transform 1 0 2000 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8748
timestamp 1677677812
transform 1 0 2100 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9922
timestamp 1677677812
transform 1 0 2100 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10002
timestamp 1677677812
transform 1 0 2020 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10003
timestamp 1677677812
transform 1 0 2052 0 1 125
box -2 -2 2 2
use FILL  FILL_10668
timestamp 1677677812
transform 1 0 2008 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8788
timestamp 1677677812
transform 1 0 2060 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_8810
timestamp 1677677812
transform 1 0 2052 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8833
timestamp 1677677812
transform 1 0 2076 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_8834
timestamp 1677677812
transform 1 0 2108 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_8846
timestamp 1677677812
transform 1 0 2092 0 1 85
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_621
timestamp 1677677812
transform -1 0 2112 0 -1 170
box -8 -3 104 105
use FILL  FILL_10669
timestamp 1677677812
transform 1 0 2112 0 -1 170
box -8 -3 16 105
use FILL  FILL_10670
timestamp 1677677812
transform 1 0 2120 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8722
timestamp 1677677812
transform 1 0 2220 0 1 165
box -3 -3 3 3
use M3_M2  M3_M2_8749
timestamp 1677677812
transform 1 0 2140 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9923
timestamp 1677677812
transform 1 0 2140 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10004
timestamp 1677677812
transform 1 0 2164 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10005
timestamp 1677677812
transform 1 0 2220 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8811
timestamp 1677677812
transform 1 0 2140 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8812
timestamp 1677677812
transform 1 0 2164 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8842
timestamp 1677677812
transform 1 0 2156 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_8843
timestamp 1677677812
transform 1 0 2180 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_8847
timestamp 1677677812
transform 1 0 2204 0 1 85
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_622
timestamp 1677677812
transform 1 0 2128 0 -1 170
box -8 -3 104 105
use FILL  FILL_10671
timestamp 1677677812
transform 1 0 2224 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8750
timestamp 1677677812
transform 1 0 2244 0 1 145
box -3 -3 3 3
use FILL  FILL_10672
timestamp 1677677812
transform 1 0 2232 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8751
timestamp 1677677812
transform 1 0 2260 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8752
timestamp 1677677812
transform 1 0 2276 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9924
timestamp 1677677812
transform 1 0 2260 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10006
timestamp 1677677812
transform 1 0 2284 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10007
timestamp 1677677812
transform 1 0 2340 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8835
timestamp 1677677812
transform 1 0 2252 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_8836
timestamp 1677677812
transform 1 0 2284 0 1 105
box -3 -3 3 3
use FILL  FILL_10673
timestamp 1677677812
transform 1 0 2240 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8844
timestamp 1677677812
transform 1 0 2276 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_8845
timestamp 1677677812
transform 1 0 2300 0 1 95
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_623
timestamp 1677677812
transform 1 0 2248 0 -1 170
box -8 -3 104 105
use FILL  FILL_10674
timestamp 1677677812
transform 1 0 2344 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8753
timestamp 1677677812
transform 1 0 2364 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8754
timestamp 1677677812
transform 1 0 2388 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9925
timestamp 1677677812
transform 1 0 2364 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10008
timestamp 1677677812
transform 1 0 2388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10009
timestamp 1677677812
transform 1 0 2412 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_624
timestamp 1677677812
transform 1 0 2352 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_9926
timestamp 1677677812
transform 1 0 2460 0 1 135
box -2 -2 2 2
use FILL  FILL_10675
timestamp 1677677812
transform 1 0 2448 0 -1 170
box -8 -3 16 105
use FILL  FILL_10676
timestamp 1677677812
transform 1 0 2456 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10010
timestamp 1677677812
transform 1 0 2484 0 1 125
box -2 -2 2 2
use INVX2  INVX2_702
timestamp 1677677812
transform 1 0 2464 0 -1 170
box -9 -3 26 105
use FILL  FILL_10677
timestamp 1677677812
transform 1 0 2480 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8755
timestamp 1677677812
transform 1 0 2580 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9927
timestamp 1677677812
transform 1 0 2580 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10011
timestamp 1677677812
transform 1 0 2500 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10012
timestamp 1677677812
transform 1 0 2556 0 1 125
box -2 -2 2 2
use FILL  FILL_10692
timestamp 1677677812
transform 1 0 2488 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10050
timestamp 1677677812
transform 1 0 2596 0 1 115
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_625
timestamp 1677677812
transform -1 0 2592 0 -1 170
box -8 -3 104 105
use FILL  FILL_10693
timestamp 1677677812
transform 1 0 2592 0 -1 170
box -8 -3 16 105
use FILL  FILL_10694
timestamp 1677677812
transform 1 0 2600 0 -1 170
box -8 -3 16 105
use FILL  FILL_10695
timestamp 1677677812
transform 1 0 2608 0 -1 170
box -8 -3 16 105
use FILL  FILL_10696
timestamp 1677677812
transform 1 0 2616 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8723
timestamp 1677677812
transform 1 0 2644 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8776
timestamp 1677677812
transform 1 0 2636 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8756
timestamp 1677677812
transform 1 0 2660 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8757
timestamp 1677677812
transform 1 0 2708 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9928
timestamp 1677677812
transform 1 0 2644 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9929
timestamp 1677677812
transform 1 0 2660 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10013
timestamp 1677677812
transform 1 0 2636 0 1 125
box -2 -2 2 2
use NAND2X1  NAND2X1_55
timestamp 1677677812
transform -1 0 2648 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_8789
timestamp 1677677812
transform 1 0 2660 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_10014
timestamp 1677677812
transform 1 0 2708 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_626
timestamp 1677677812
transform 1 0 2648 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8724
timestamp 1677677812
transform 1 0 2780 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9894
timestamp 1677677812
transform 1 0 2764 0 1 145
box -2 -2 2 2
use M3_M2  M3_M2_8758
timestamp 1677677812
transform 1 0 2772 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9930
timestamp 1677677812
transform 1 0 2772 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10015
timestamp 1677677812
transform 1 0 2764 0 1 125
box -2 -2 2 2
use INVX2  INVX2_705
timestamp 1677677812
transform 1 0 2744 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_10016
timestamp 1677677812
transform 1 0 2780 0 1 125
box -2 -2 2 2
use NOR2X1  NOR2X1_121
timestamp 1677677812
transform 1 0 2760 0 -1 170
box -8 -3 32 105
use FILL  FILL_10697
timestamp 1677677812
transform 1 0 2784 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8777
timestamp 1677677812
transform 1 0 2804 0 1 135
box -3 -3 3 3
use M3_M2  M3_M2_8813
timestamp 1677677812
transform 1 0 2804 0 1 115
box -3 -3 3 3
use FILL  FILL_10698
timestamp 1677677812
transform 1 0 2792 0 -1 170
box -8 -3 16 105
use FILL  FILL_10699
timestamp 1677677812
transform 1 0 2800 0 -1 170
box -8 -3 16 105
use FILL  FILL_10700
timestamp 1677677812
transform 1 0 2808 0 -1 170
box -8 -3 16 105
use FILL  FILL_10701
timestamp 1677677812
transform 1 0 2816 0 -1 170
box -8 -3 16 105
use FILL  FILL_10703
timestamp 1677677812
transform 1 0 2824 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8759
timestamp 1677677812
transform 1 0 2844 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9931
timestamp 1677677812
transform 1 0 2844 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9932
timestamp 1677677812
transform 1 0 2860 0 1 135
box -2 -2 2 2
use FILL  FILL_10711
timestamp 1677677812
transform 1 0 2832 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8778
timestamp 1677677812
transform 1 0 2868 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9933
timestamp 1677677812
transform 1 0 2876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10017
timestamp 1677677812
transform 1 0 2868 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10018
timestamp 1677677812
transform 1 0 2884 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8814
timestamp 1677677812
transform 1 0 2868 0 1 115
box -3 -3 3 3
use OAI22X1  OAI22X1_441
timestamp 1677677812
transform 1 0 2840 0 -1 170
box -8 -3 46 105
use M3_M2  M3_M2_8760
timestamp 1677677812
transform 1 0 2900 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9934
timestamp 1677677812
transform 1 0 2892 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10019
timestamp 1677677812
transform 1 0 2900 0 1 125
box -2 -2 2 2
use INVX2  INVX2_707
timestamp 1677677812
transform -1 0 2896 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_8725
timestamp 1677677812
transform 1 0 2908 0 1 155
box -3 -3 3 3
use FILL  FILL_10712
timestamp 1677677812
transform 1 0 2896 0 -1 170
box -8 -3 16 105
use FILL  FILL_10713
timestamp 1677677812
transform 1 0 2904 0 -1 170
box -8 -3 16 105
use FILL  FILL_10714
timestamp 1677677812
transform 1 0 2912 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9935
timestamp 1677677812
transform 1 0 2932 0 1 135
box -2 -2 2 2
use INVX2  INVX2_708
timestamp 1677677812
transform -1 0 2936 0 -1 170
box -9 -3 26 105
use FILL  FILL_10715
timestamp 1677677812
transform 1 0 2936 0 -1 170
box -8 -3 16 105
use FILL  FILL_10723
timestamp 1677677812
transform 1 0 2944 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8779
timestamp 1677677812
transform 1 0 2988 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9936
timestamp 1677677812
transform 1 0 3036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10020
timestamp 1677677812
transform 1 0 2988 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8790
timestamp 1677677812
transform 1 0 3036 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_8726
timestamp 1677677812
transform 1 0 3052 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_10021
timestamp 1677677812
transform 1 0 3052 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_629
timestamp 1677677812
transform -1 0 3048 0 -1 170
box -8 -3 104 105
use FILL  FILL_10724
timestamp 1677677812
transform 1 0 3048 0 -1 170
box -8 -3 16 105
use FILL  FILL_10725
timestamp 1677677812
transform 1 0 3056 0 -1 170
box -8 -3 16 105
use FILL  FILL_10726
timestamp 1677677812
transform 1 0 3064 0 -1 170
box -8 -3 16 105
use FILL  FILL_10727
timestamp 1677677812
transform 1 0 3072 0 -1 170
box -8 -3 16 105
use FILL  FILL_10728
timestamp 1677677812
transform 1 0 3080 0 -1 170
box -8 -3 16 105
use FILL  FILL_10729
timestamp 1677677812
transform 1 0 3088 0 -1 170
box -8 -3 16 105
use FILL  FILL_10730
timestamp 1677677812
transform 1 0 3096 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9937
timestamp 1677677812
transform 1 0 3188 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10022
timestamp 1677677812
transform 1 0 3164 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8815
timestamp 1677677812
transform 1 0 3164 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_630
timestamp 1677677812
transform -1 0 3200 0 -1 170
box -8 -3 104 105
use FILL  FILL_10731
timestamp 1677677812
transform 1 0 3200 0 -1 170
box -8 -3 16 105
use FILL  FILL_10733
timestamp 1677677812
transform 1 0 3208 0 -1 170
box -8 -3 16 105
use FILL  FILL_10735
timestamp 1677677812
transform 1 0 3216 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9938
timestamp 1677677812
transform 1 0 3236 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10023
timestamp 1677677812
transform 1 0 3260 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8816
timestamp 1677677812
transform 1 0 3260 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_632
timestamp 1677677812
transform 1 0 3224 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_8727
timestamp 1677677812
transform 1 0 3332 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9939
timestamp 1677677812
transform 1 0 3332 0 1 135
box -2 -2 2 2
use FILL  FILL_10737
timestamp 1677677812
transform 1 0 3320 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_710
timestamp 1677677812
transform 1 0 3328 0 -1 170
box -9 -3 26 105
use FILL  FILL_10739
timestamp 1677677812
transform 1 0 3344 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8728
timestamp 1677677812
transform 1 0 3364 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8761
timestamp 1677677812
transform 1 0 3372 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9940
timestamp 1677677812
transform 1 0 3372 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10024
timestamp 1677677812
transform 1 0 3364 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8837
timestamp 1677677812
transform 1 0 3364 0 1 105
box -3 -3 3 3
use FILL  FILL_10740
timestamp 1677677812
transform 1 0 3352 0 -1 170
box -8 -3 16 105
use FILL  FILL_10742
timestamp 1677677812
transform 1 0 3360 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8762
timestamp 1677677812
transform 1 0 3396 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9941
timestamp 1677677812
transform 1 0 3396 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10025
timestamp 1677677812
transform 1 0 3388 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_9942
timestamp 1677677812
transform 1 0 3420 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10051
timestamp 1677677812
transform 1 0 3396 0 1 115
box -2 -2 2 2
use NAND2X1  NAND2X1_59
timestamp 1677677812
transform 1 0 3368 0 -1 170
box -8 -3 32 105
use M3_M2  M3_M2_8817
timestamp 1677677812
transform 1 0 3404 0 1 115
box -3 -3 3 3
use M2_M1  M2_M1_10052
timestamp 1677677812
transform 1 0 3412 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_8818
timestamp 1677677812
transform 1 0 3420 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8838
timestamp 1677677812
transform 1 0 3412 0 1 105
box -3 -3 3 3
use NAND2X1  NAND2X1_60
timestamp 1677677812
transform 1 0 3392 0 -1 170
box -8 -3 32 105
use M2_M1  M2_M1_9943
timestamp 1677677812
transform 1 0 3444 0 1 135
box -2 -2 2 2
use OAI21X1  OAI21X1_186
timestamp 1677677812
transform 1 0 3416 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_8763
timestamp 1677677812
transform 1 0 3468 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8764
timestamp 1677677812
transform 1 0 3492 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8765
timestamp 1677677812
transform 1 0 3516 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9944
timestamp 1677677812
transform 1 0 3468 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10026
timestamp 1677677812
transform 1 0 3516 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10053
timestamp 1677677812
transform 1 0 3452 0 1 115
box -2 -2 2 2
use FILL  FILL_10749
timestamp 1677677812
transform 1 0 3448 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8819
timestamp 1677677812
transform 1 0 3492 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_634
timestamp 1677677812
transform 1 0 3456 0 -1 170
box -8 -3 104 105
use FILL  FILL_10750
timestamp 1677677812
transform 1 0 3552 0 -1 170
box -8 -3 16 105
use FILL  FILL_10751
timestamp 1677677812
transform 1 0 3560 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10027
timestamp 1677677812
transform 1 0 3588 0 1 125
box -2 -2 2 2
use INVX2  INVX2_711
timestamp 1677677812
transform 1 0 3568 0 -1 170
box -9 -3 26 105
use FILL  FILL_10752
timestamp 1677677812
transform 1 0 3584 0 -1 170
box -8 -3 16 105
use FILL  FILL_10754
timestamp 1677677812
transform 1 0 3592 0 -1 170
box -8 -3 16 105
use FILL  FILL_10756
timestamp 1677677812
transform 1 0 3600 0 -1 170
box -8 -3 16 105
use FILL  FILL_10764
timestamp 1677677812
transform 1 0 3608 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8766
timestamp 1677677812
transform 1 0 3628 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9945
timestamp 1677677812
transform 1 0 3628 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8780
timestamp 1677677812
transform 1 0 3676 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10028
timestamp 1677677812
transform 1 0 3676 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8820
timestamp 1677677812
transform 1 0 3628 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8781
timestamp 1677677812
transform 1 0 3716 0 1 135
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_635
timestamp 1677677812
transform 1 0 3616 0 -1 170
box -8 -3 104 105
use FILL  FILL_10765
timestamp 1677677812
transform 1 0 3712 0 -1 170
box -8 -3 16 105
use FILL  FILL_10766
timestamp 1677677812
transform 1 0 3720 0 -1 170
box -8 -3 16 105
use FILL  FILL_10767
timestamp 1677677812
transform 1 0 3728 0 -1 170
box -8 -3 16 105
use FILL  FILL_10768
timestamp 1677677812
transform 1 0 3736 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_10029
timestamp 1677677812
transform 1 0 3756 0 1 125
box -2 -2 2 2
use INVX2  INVX2_717
timestamp 1677677812
transform 1 0 3744 0 -1 170
box -9 -3 26 105
use FILL  FILL_10793
timestamp 1677677812
transform 1 0 3760 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8767
timestamp 1677677812
transform 1 0 3780 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9946
timestamp 1677677812
transform 1 0 3780 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8729
timestamp 1677677812
transform 1 0 3876 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9947
timestamp 1677677812
transform 1 0 3876 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10030
timestamp 1677677812
transform 1 0 3828 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10031
timestamp 1677677812
transform 1 0 3860 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10032
timestamp 1677677812
transform 1 0 3868 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8821
timestamp 1677677812
transform 1 0 3780 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8822
timestamp 1677677812
transform 1 0 3820 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8823
timestamp 1677677812
transform 1 0 3868 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_638
timestamp 1677677812
transform 1 0 3768 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_718
timestamp 1677677812
transform -1 0 3880 0 -1 170
box -9 -3 26 105
use FILL  FILL_10794
timestamp 1677677812
transform 1 0 3880 0 -1 170
box -8 -3 16 105
use FILL  FILL_10795
timestamp 1677677812
transform 1 0 3888 0 -1 170
box -8 -3 16 105
use FILL  FILL_10796
timestamp 1677677812
transform 1 0 3896 0 -1 170
box -8 -3 16 105
use FILL  FILL_10797
timestamp 1677677812
transform 1 0 3904 0 -1 170
box -8 -3 16 105
use FILL  FILL_10798
timestamp 1677677812
transform 1 0 3912 0 -1 170
box -8 -3 16 105
use FILL  FILL_10799
timestamp 1677677812
transform 1 0 3920 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8730
timestamp 1677677812
transform 1 0 3940 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8768
timestamp 1677677812
transform 1 0 3972 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9948
timestamp 1677677812
transform 1 0 3940 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8782
timestamp 1677677812
transform 1 0 4020 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_10033
timestamp 1677677812
transform 1 0 3964 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10034
timestamp 1677677812
transform 1 0 4020 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10035
timestamp 1677677812
transform 1 0 4036 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8824
timestamp 1677677812
transform 1 0 4020 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_639
timestamp 1677677812
transform 1 0 3928 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_719
timestamp 1677677812
transform -1 0 4040 0 -1 170
box -9 -3 26 105
use M2_M1  M2_M1_10036
timestamp 1677677812
transform 1 0 4052 0 1 125
box -2 -2 2 2
use FILL  FILL_10800
timestamp 1677677812
transform 1 0 4040 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_9949
timestamp 1677677812
transform 1 0 4060 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_8825
timestamp 1677677812
transform 1 0 4060 0 1 115
box -3 -3 3 3
use FILL  FILL_10801
timestamp 1677677812
transform 1 0 4048 0 -1 170
box -8 -3 16 105
use FILL  FILL_10802
timestamp 1677677812
transform 1 0 4056 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8731
timestamp 1677677812
transform 1 0 4164 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_8769
timestamp 1677677812
transform 1 0 4140 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8783
timestamp 1677677812
transform 1 0 4116 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_9950
timestamp 1677677812
transform 1 0 4164 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10037
timestamp 1677677812
transform 1 0 4084 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10038
timestamp 1677677812
transform 1 0 4116 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8826
timestamp 1677677812
transform 1 0 4084 0 1 115
box -3 -3 3 3
use INVX2  INVX2_720
timestamp 1677677812
transform -1 0 4080 0 -1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_640
timestamp 1677677812
transform -1 0 4176 0 -1 170
box -8 -3 104 105
use FILL  FILL_10803
timestamp 1677677812
transform 1 0 4176 0 -1 170
box -8 -3 16 105
use FILL  FILL_10804
timestamp 1677677812
transform 1 0 4184 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8732
timestamp 1677677812
transform 1 0 4204 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9951
timestamp 1677677812
transform 1 0 4204 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10039
timestamp 1677677812
transform 1 0 4252 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_641
timestamp 1677677812
transform 1 0 4192 0 -1 170
box -8 -3 104 105
use M2_M1  M2_M1_10040
timestamp 1677677812
transform 1 0 4300 0 1 125
box -2 -2 2 2
use FILL  FILL_10805
timestamp 1677677812
transform 1 0 4288 0 -1 170
box -8 -3 16 105
use FILL  FILL_10806
timestamp 1677677812
transform 1 0 4296 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8733
timestamp 1677677812
transform 1 0 4316 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_9952
timestamp 1677677812
transform 1 0 4316 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10041
timestamp 1677677812
transform 1 0 4340 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10042
timestamp 1677677812
transform 1 0 4396 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_642
timestamp 1677677812
transform 1 0 4304 0 -1 170
box -8 -3 104 105
use FILL  FILL_10807
timestamp 1677677812
transform 1 0 4400 0 -1 170
box -8 -3 16 105
use FILL  FILL_10809
timestamp 1677677812
transform 1 0 4408 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8770
timestamp 1677677812
transform 1 0 4428 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9953
timestamp 1677677812
transform 1 0 4428 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10043
timestamp 1677677812
transform 1 0 4452 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10044
timestamp 1677677812
transform 1 0 4508 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_643
timestamp 1677677812
transform 1 0 4416 0 -1 170
box -8 -3 104 105
use FILL  FILL_10816
timestamp 1677677812
transform 1 0 4512 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8771
timestamp 1677677812
transform 1 0 4532 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9954
timestamp 1677677812
transform 1 0 4532 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10045
timestamp 1677677812
transform 1 0 4556 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10046
timestamp 1677677812
transform 1 0 4612 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_645
timestamp 1677677812
transform 1 0 4520 0 -1 170
box -8 -3 104 105
use FILL  FILL_10825
timestamp 1677677812
transform 1 0 4616 0 -1 170
box -8 -3 16 105
use FILL  FILL_10826
timestamp 1677677812
transform 1 0 4624 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_8772
timestamp 1677677812
transform 1 0 4644 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_8773
timestamp 1677677812
transform 1 0 4708 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_9955
timestamp 1677677812
transform 1 0 4644 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_9956
timestamp 1677677812
transform 1 0 4740 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_10047
timestamp 1677677812
transform 1 0 4676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10048
timestamp 1677677812
transform 1 0 4724 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_10049
timestamp 1677677812
transform 1 0 4732 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_8827
timestamp 1677677812
transform 1 0 4684 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_8828
timestamp 1677677812
transform 1 0 4732 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_646
timestamp 1677677812
transform 1 0 4632 0 -1 170
box -8 -3 104 105
use INVX2  INVX2_724
timestamp 1677677812
transform -1 0 4744 0 -1 170
box -9 -3 26 105
use FILL  FILL_10827
timestamp 1677677812
transform 1 0 4744 0 -1 170
box -8 -3 16 105
use FILL  FILL_10828
timestamp 1677677812
transform 1 0 4752 0 -1 170
box -8 -3 16 105
use FILL  FILL_10829
timestamp 1677677812
transform 1 0 4760 0 -1 170
box -8 -3 16 105
use FILL  FILL_10830
timestamp 1677677812
transform 1 0 4768 0 -1 170
box -8 -3 16 105
use FILL  FILL_10831
timestamp 1677677812
transform 1 0 4776 0 -1 170
box -8 -3 16 105
use FILL  FILL_10832
timestamp 1677677812
transform 1 0 4784 0 -1 170
box -8 -3 16 105
use top_level_VIA0  top_level_VIA0_93
timestamp 1677677812
transform 1 0 4843 0 1 70
box -10 -3 10 3
use top_level_VIA1  top_level_VIA1_4
timestamp 1677677812
transform 1 0 48 0 1 47
box -10 -10 10 10
use top_level_VIA1  top_level_VIA1_6
timestamp 1677677812
transform 1 0 24 0 1 23
box -10 -10 10 10
use M3_M2  M3_M2_8848
timestamp 1677677812
transform 1 0 2020 0 1 35
box -3 -3 3 3
use M3_M2  M3_M2_8849
timestamp 1677677812
transform 1 0 2308 0 1 35
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_5
timestamp 1677677812
transform 1 0 4819 0 1 47
box -10 -10 10 10
use M3_M2  M3_M2_8850
timestamp 1677677812
transform 1 0 2060 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8851
timestamp 1677677812
transform 1 0 2324 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8852
timestamp 1677677812
transform 1 0 2364 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_8853
timestamp 1677677812
transform 1 0 2668 0 1 15
box -3 -3 3 3
use top_level_VIA1  top_level_VIA1_7
timestamp 1677677812
transform 1 0 4843 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal2 2668 1 2668 1 4 clka
rlabel metal3 2 2015 2 2015 4 clkb
rlabel metal2 2372 1 2372 1 4 reset
rlabel metal2 2532 1 2532 1 4 we_ins
rlabel metal2 2108 1 2108 1 4 load[15]
rlabel metal2 2076 1 2076 1 4 load[14]
rlabel metal2 2036 1 2036 1 4 load[13]
rlabel metal2 2092 1 2092 1 4 load[12]
rlabel metal2 2060 1 2060 1 4 load[11]
rlabel metal2 2020 1 2020 1 4 load[10]
rlabel metal2 2124 1 2124 1 4 load[9]
rlabel metal2 2252 1 2252 1 4 load[8]
rlabel metal2 2212 1 2212 1 4 load[7]
rlabel metal2 2140 1 2140 1 4 load[6]
rlabel metal2 2004 1 2004 1 4 load[5]
rlabel metal2 2276 1 2276 1 4 load[4]
rlabel metal2 2172 1 2172 1 4 load[3]
rlabel metal2 2236 1 2236 1 4 load[2]
rlabel metal2 2156 1 2156 1 4 load[1]
rlabel metal2 1988 1 1988 1 4 load[0]
rlabel metal2 4060 1 4060 1 4 reg_0_out[7]
rlabel metal2 3860 1 3860 1 4 reg_0_out[6]
rlabel metal2 4100 1 4100 1 4 reg_0_out[5]
rlabel metal2 3844 1 3844 1 4 reg_0_out[4]
rlabel metal2 3708 1 3708 1 4 reg_0_out[3]
rlabel metal2 3684 1 3684 1 4 reg_0_out[2]
rlabel metal2 4084 1 4084 1 4 reg_0_out[1]
rlabel metal2 3940 1 3940 1 4 reg_0_out[0]
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
<< end >>

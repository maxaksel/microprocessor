magic
tech scmos
timestamp 1682952543
<< nwell >>
rect -8 48 46 105
<< ntransistor >>
rect 9 6 11 26
rect 14 6 16 26
rect 26 6 28 26
rect 31 6 33 26
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
rect 31 54 33 94
<< ndiffusion >>
rect 4 6 9 26
rect 11 6 14 26
rect 16 6 26 26
rect 28 6 31 26
rect 33 6 38 26
<< pdiffusion >>
rect 2 54 7 94
rect 9 54 15 94
rect 17 54 23 94
rect 25 54 31 94
rect 33 54 38 94
<< psubstratepdiff >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
<< nsubstratendiff >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 7 49 9 54
rect 15 53 17 54
rect 14 51 17 53
rect 6 47 10 49
rect 4 45 10 47
rect 4 29 6 45
rect 14 41 16 51
rect 10 37 16 41
rect 23 43 25 54
rect 31 53 33 54
rect 31 51 35 53
rect 33 47 38 51
rect 23 40 29 43
rect 4 27 11 29
rect 9 26 11 27
rect 14 26 16 37
rect 24 39 29 40
rect 24 29 26 39
rect 33 31 35 47
rect 31 29 35 31
rect 24 27 28 29
rect 26 26 28 27
rect 31 26 33 29
rect 9 4 11 6
rect 14 4 16 6
rect 26 4 28 6
rect 31 4 33 6
<< genericcontact >>
rect -1 99 1 101
rect 15 99 17 101
rect 31 99 33 101
rect 11 91 13 93
rect 3 89 5 91
rect 19 90 21 92
rect 35 90 37 92
rect 11 86 13 88
rect 3 84 5 86
rect 19 85 21 87
rect 27 85 29 87
rect 35 85 37 87
rect 11 81 13 83
rect 3 79 5 81
rect 19 80 21 82
rect 27 80 29 82
rect 35 80 37 82
rect 11 76 13 78
rect 3 74 5 76
rect 19 75 21 77
rect 27 75 29 77
rect 35 75 37 77
rect 11 71 13 73
rect 3 69 5 71
rect 19 70 21 72
rect 27 70 29 72
rect 35 70 37 72
rect 11 66 13 68
rect 3 64 5 66
rect 19 65 21 67
rect 27 65 29 67
rect 35 65 37 67
rect 11 61 13 63
rect 3 59 5 61
rect 19 60 21 62
rect 27 60 29 62
rect 35 60 37 62
rect 19 55 21 57
rect 27 55 29 57
rect 35 55 37 57
rect 35 48 37 50
rect 7 46 9 48
rect 26 40 28 42
rect 11 38 13 40
rect 5 22 7 24
rect 20 22 22 24
rect 35 22 37 24
rect 5 17 7 19
rect 20 17 22 19
rect 35 17 37 19
rect 5 12 7 14
rect 20 12 22 14
rect 35 12 37 14
rect 5 7 7 9
rect 20 7 22 9
rect 35 7 37 9
rect -1 -1 1 1
rect 15 -1 17 1
rect 31 -1 33 1
<< metal1 >>
rect -2 97 42 103
rect 2 57 6 94
rect 10 60 14 97
rect 18 91 38 94
rect 18 57 22 91
rect 2 54 22 57
rect 26 54 30 88
rect 34 54 38 91
rect 26 51 29 54
rect 6 47 10 49
rect 19 48 29 51
rect 19 47 22 48
rect 2 44 10 47
rect 2 43 6 44
rect 18 43 22 47
rect 34 43 38 51
rect 10 33 14 41
rect 19 26 22 43
rect 25 39 29 43
rect 26 37 29 39
rect 26 33 30 37
rect 4 3 8 26
rect 17 6 25 26
rect 34 3 38 26
rect -2 -3 42 3
<< m1p >>
rect 2 43 6 47
rect 18 43 22 47
rect 34 43 38 47
rect 10 33 14 37
rect 26 33 30 37
<< labels >>
rlabel metal1 4 0 4 0 8 gnd
rlabel metal1 4 100 4 100 6 vdd
rlabel metal1 36 45 36 45 6 C
rlabel metal1 28 35 28 35 6 D
rlabel metal1 20 45 20 45 6 Y
rlabel metal1 4 45 4 45 6 A
rlabel metal1 12 35 12 35 6 B
<< end >>
